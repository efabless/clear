magic
tech sky130A
magscale 1 2
timestamp 1681041584
<< viali >>
rect 3985 24361 4019 24395
rect 6561 24361 6595 24395
rect 11713 24361 11747 24395
rect 23857 24361 23891 24395
rect 25789 24361 25823 24395
rect 31309 24361 31343 24395
rect 34161 24361 34195 24395
rect 39313 24361 39347 24395
rect 44741 24361 44775 24395
rect 27169 24293 27203 24327
rect 29009 24293 29043 24327
rect 36369 24293 36403 24327
rect 37473 24293 37507 24327
rect 38669 24293 38703 24327
rect 3249 24225 3283 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 13553 24225 13587 24259
rect 16129 24225 16163 24259
rect 16865 24225 16899 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25053 24225 25087 24259
rect 25237 24225 25271 24259
rect 26341 24225 26375 24259
rect 27629 24225 27663 24259
rect 27721 24225 27755 24259
rect 29745 24225 29779 24259
rect 30021 24225 30055 24259
rect 37013 24225 37047 24259
rect 40049 24225 40083 24259
rect 40325 24225 40359 24259
rect 2237 24157 2271 24191
rect 3893 24157 3927 24191
rect 4169 24157 4203 24191
rect 4629 24157 4663 24191
rect 6469 24157 6503 24191
rect 6745 24157 6779 24191
rect 7389 24157 7423 24191
rect 9321 24157 9355 24191
rect 9965 24157 9999 24191
rect 11897 24157 11931 24191
rect 12541 24157 12575 24191
rect 14473 24157 14507 24191
rect 15117 24157 15151 24191
rect 18981 24157 19015 24191
rect 19625 24157 19659 24191
rect 20085 24157 20119 24191
rect 22017 24157 22051 24191
rect 24041 24157 24075 24191
rect 26157 24157 26191 24191
rect 26249 24157 26283 24191
rect 28549 24157 28583 24191
rect 29193 24157 29227 24191
rect 31493 24157 31527 24191
rect 32505 24157 32539 24191
rect 33333 24157 33367 24191
rect 34069 24157 34103 24191
rect 36553 24157 36587 24191
rect 37657 24157 37691 24191
rect 38485 24157 38519 24191
rect 39221 24157 39255 24191
rect 41429 24157 41463 24191
rect 42441 24157 42475 24191
rect 44373 24157 44407 24191
rect 45201 24157 45235 24191
rect 45937 24157 45971 24191
rect 46673 24157 46707 24191
rect 47225 24157 47259 24191
rect 47777 24157 47811 24191
rect 48605 24157 48639 24191
rect 10977 24089 11011 24123
rect 17141 24089 17175 24123
rect 27537 24089 27571 24123
rect 32781 24089 32815 24123
rect 34989 24089 35023 24123
rect 35725 24089 35759 24123
rect 37933 24089 37967 24123
rect 1593 24021 1627 24055
rect 1685 24021 1719 24055
rect 9137 24021 9171 24055
rect 14289 24021 14323 24055
rect 18613 24021 18647 24055
rect 19441 24021 19475 24055
rect 24593 24021 24627 24055
rect 24961 24021 24995 24055
rect 28365 24021 28399 24055
rect 30941 24021 30975 24055
rect 31861 24021 31895 24055
rect 32321 24021 32355 24055
rect 33425 24021 33459 24055
rect 35081 24021 35115 24055
rect 35817 24021 35851 24055
rect 36829 24021 36863 24055
rect 42073 24021 42107 24055
rect 44189 24021 44223 24055
rect 45385 24021 45419 24055
rect 46121 24021 46155 24055
rect 46857 24021 46891 24055
rect 47961 24021 47995 24055
rect 49249 24021 49283 24055
rect 1777 23817 1811 23851
rect 11897 23817 11931 23851
rect 12265 23817 12299 23851
rect 12357 23817 12391 23851
rect 24225 23817 24259 23851
rect 29377 23817 29411 23851
rect 33425 23817 33459 23851
rect 34069 23817 34103 23851
rect 34805 23817 34839 23851
rect 38485 23817 38519 23851
rect 39037 23817 39071 23851
rect 39865 23817 39899 23851
rect 40325 23817 40359 23851
rect 40693 23817 40727 23851
rect 46305 23817 46339 23851
rect 47593 23817 47627 23851
rect 1593 23749 1627 23783
rect 3985 23749 4019 23783
rect 9137 23749 9171 23783
rect 10977 23749 11011 23783
rect 14289 23749 14323 23783
rect 16129 23749 16163 23783
rect 18981 23749 19015 23783
rect 21189 23749 21223 23783
rect 22293 23749 22327 23783
rect 25145 23749 25179 23783
rect 30113 23749 30147 23783
rect 32965 23749 32999 23783
rect 35633 23749 35667 23783
rect 38669 23749 38703 23783
rect 46213 23749 46247 23783
rect 2145 23681 2179 23715
rect 2789 23681 2823 23715
rect 4813 23681 4847 23715
rect 7113 23681 7147 23715
rect 7205 23681 7239 23715
rect 7941 23681 7975 23715
rect 9873 23681 9907 23715
rect 13277 23681 13311 23715
rect 15117 23681 15151 23715
rect 16865 23681 16899 23715
rect 18705 23681 18739 23715
rect 21005 23681 21039 23715
rect 29561 23681 29595 23715
rect 30297 23681 30331 23715
rect 30849 23681 30883 23715
rect 31033 23681 31067 23715
rect 31501 23685 31535 23719
rect 33977 23681 34011 23715
rect 34713 23681 34747 23715
rect 35449 23681 35483 23715
rect 36277 23681 36311 23715
rect 36921 23681 36955 23715
rect 37289 23681 37323 23715
rect 37933 23681 37967 23715
rect 38209 23681 38243 23715
rect 40877 23681 40911 23715
rect 41521 23681 41555 23715
rect 41797 23681 41831 23715
rect 42625 23681 42659 23715
rect 43729 23681 43763 23715
rect 44833 23681 44867 23715
rect 45569 23681 45603 23715
rect 46765 23681 46799 23715
rect 47317 23681 47351 23715
rect 47961 23681 47995 23715
rect 48697 23681 48731 23715
rect 5457 23613 5491 23647
rect 6469 23613 6503 23647
rect 7389 23613 7423 23647
rect 12541 23613 12575 23647
rect 17877 23613 17911 23647
rect 22017 23613 22051 23647
rect 24869 23613 24903 23647
rect 27169 23613 27203 23647
rect 27445 23613 27479 23647
rect 32321 23613 32355 23647
rect 6745 23545 6779 23579
rect 21649 23545 21683 23579
rect 30665 23545 30699 23579
rect 36737 23545 36771 23579
rect 41337 23545 41371 23579
rect 44373 23545 44407 23579
rect 45017 23545 45051 23579
rect 2237 23477 2271 23511
rect 6561 23477 6595 23511
rect 11529 23477 11563 23511
rect 20453 23477 20487 23511
rect 23765 23477 23799 23511
rect 26617 23477 26651 23511
rect 28917 23477 28951 23511
rect 31309 23477 31343 23511
rect 31861 23477 31895 23511
rect 36093 23477 36127 23511
rect 37749 23477 37783 23511
rect 43269 23477 43303 23511
rect 45753 23477 45787 23511
rect 46949 23477 46983 23511
rect 48145 23477 48179 23511
rect 49341 23477 49375 23511
rect 14473 23273 14507 23307
rect 20348 23273 20382 23307
rect 25789 23273 25823 23307
rect 27524 23273 27558 23307
rect 29009 23273 29043 23307
rect 30002 23273 30036 23307
rect 36645 23273 36679 23307
rect 36829 23273 36863 23307
rect 37289 23273 37323 23307
rect 44005 23273 44039 23307
rect 44649 23273 44683 23307
rect 49341 23273 49375 23307
rect 18889 23205 18923 23239
rect 26801 23205 26835 23239
rect 32597 23205 32631 23239
rect 33333 23205 33367 23239
rect 34069 23205 34103 23239
rect 34897 23205 34931 23239
rect 37013 23205 37047 23239
rect 4721 23137 4755 23171
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 11529 23137 11563 23171
rect 13277 23137 13311 23171
rect 16497 23137 16531 23171
rect 20085 23137 20119 23171
rect 21833 23137 21867 23171
rect 22569 23137 22603 23171
rect 25145 23137 25179 23171
rect 26341 23137 26375 23171
rect 27261 23137 27295 23171
rect 47501 23137 47535 23171
rect 1777 23069 1811 23103
rect 3433 23069 3467 23103
rect 3617 23069 3651 23103
rect 5365 23069 5399 23103
rect 7205 23069 7239 23103
rect 9321 23069 9355 23103
rect 13921 23069 13955 23103
rect 14381 23069 14415 23103
rect 15485 23069 15519 23103
rect 17141 23069 17175 23103
rect 19625 23069 19659 23103
rect 22293 23069 22327 23103
rect 24961 23069 24995 23103
rect 29745 23069 29779 23103
rect 31861 23069 31895 23103
rect 35081 23069 35115 23103
rect 35725 23069 35759 23103
rect 41153 23069 41187 23103
rect 43361 23069 43395 23103
rect 47685 23069 47719 23103
rect 47961 23069 47995 23103
rect 48697 23069 48731 23103
rect 2789 23001 2823 23035
rect 3801 23001 3835 23035
rect 4077 23001 4111 23035
rect 9597 23001 9631 23035
rect 11805 23001 11839 23035
rect 17417 23001 17451 23035
rect 26249 23001 26283 23035
rect 32413 23001 32447 23035
rect 33149 23001 33183 23035
rect 33885 23001 33919 23035
rect 34437 23001 34471 23035
rect 4169 22933 4203 22967
rect 4537 22933 4571 22967
rect 4629 22933 4663 22967
rect 9045 22933 9079 22967
rect 11069 22933 11103 22967
rect 13645 22933 13679 22967
rect 14933 22933 14967 22967
rect 19441 22933 19475 22967
rect 24041 22933 24075 22967
rect 24593 22933 24627 22967
rect 25053 22933 25087 22967
rect 26157 22933 26191 22967
rect 29377 22933 29411 22967
rect 31493 22933 31527 22967
rect 31953 22933 31987 22967
rect 35541 22933 35575 22967
rect 36185 22933 36219 22967
rect 42441 22933 42475 22967
rect 48145 22933 48179 22967
rect 3801 22729 3835 22763
rect 6469 22729 6503 22763
rect 14565 22729 14599 22763
rect 18613 22729 18647 22763
rect 21465 22729 21499 22763
rect 25697 22729 25731 22763
rect 25789 22729 25823 22763
rect 27169 22729 27203 22763
rect 30573 22729 30607 22763
rect 32965 22729 32999 22763
rect 33241 22729 33275 22763
rect 35081 22729 35115 22763
rect 39957 22729 39991 22763
rect 47777 22729 47811 22763
rect 10701 22661 10735 22695
rect 12725 22661 12759 22695
rect 16129 22661 16163 22695
rect 17141 22661 17175 22695
rect 22201 22661 22235 22695
rect 22477 22661 22511 22695
rect 31677 22661 31711 22695
rect 31861 22661 31895 22695
rect 47685 22661 47719 22695
rect 1777 22593 1811 22627
rect 4813 22593 4847 22627
rect 7113 22593 7147 22627
rect 7205 22593 7239 22627
rect 8125 22593 8159 22627
rect 9965 22593 9999 22627
rect 11805 22593 11839 22627
rect 15025 22593 15059 22627
rect 19257 22593 19291 22627
rect 19717 22593 19751 22627
rect 23121 22593 23155 22627
rect 27537 22593 27571 22627
rect 28365 22593 28399 22627
rect 30941 22593 30975 22627
rect 32413 22593 32447 22627
rect 33885 22593 33919 22627
rect 34989 22593 35023 22627
rect 37565 22593 37599 22627
rect 37841 22593 37875 22627
rect 43913 22593 43947 22627
rect 48053 22593 48087 22627
rect 48329 22593 48363 22627
rect 49065 22593 49099 22627
rect 2789 22525 2823 22559
rect 3893 22525 3927 22559
rect 4077 22525 4111 22559
rect 5089 22525 5123 22559
rect 7297 22525 7331 22559
rect 8677 22525 8711 22559
rect 12449 22525 12483 22559
rect 16865 22525 16899 22559
rect 19993 22525 20027 22559
rect 23397 22525 23431 22559
rect 25881 22525 25915 22559
rect 26525 22525 26559 22559
rect 26709 22525 26743 22559
rect 27629 22525 27663 22559
rect 27721 22525 27755 22559
rect 28641 22525 28675 22559
rect 31033 22525 31067 22559
rect 31125 22525 31159 22559
rect 33057 22525 33091 22559
rect 33609 22525 33643 22559
rect 38117 22525 38151 22559
rect 44557 22525 44591 22559
rect 6745 22457 6779 22491
rect 11989 22457 12023 22491
rect 34713 22457 34747 22491
rect 49249 22457 49283 22491
rect 3433 22389 3467 22423
rect 14197 22389 14231 22423
rect 19073 22389 19107 22423
rect 21925 22389 21959 22423
rect 24869 22389 24903 22423
rect 25329 22389 25363 22423
rect 26433 22389 26467 22423
rect 30113 22389 30147 22423
rect 32505 22389 32539 22423
rect 35357 22389 35391 22423
rect 39589 22389 39623 22423
rect 48513 22389 48547 22423
rect 23305 22185 23339 22219
rect 24593 22185 24627 22219
rect 26052 22185 26086 22219
rect 29561 22185 29595 22219
rect 29745 22185 29779 22219
rect 8769 22117 8803 22151
rect 27537 22117 27571 22151
rect 33885 22117 33919 22151
rect 2053 22049 2087 22083
rect 4629 22049 4663 22083
rect 5825 22049 5859 22083
rect 7941 22049 7975 22083
rect 8953 22049 8987 22083
rect 9873 22049 9907 22083
rect 11253 22049 11287 22083
rect 13369 22049 13403 22083
rect 15669 22049 15703 22083
rect 17141 22049 17175 22083
rect 20085 22049 20119 22083
rect 23949 22049 23983 22083
rect 25237 22049 25271 22083
rect 29193 22049 29227 22083
rect 30573 22049 30607 22083
rect 30757 22049 30791 22083
rect 34253 22049 34287 22083
rect 1777 21981 1811 22015
rect 3985 21981 4019 22015
rect 6285 21981 6319 22015
rect 6929 21981 6963 22015
rect 8585 21981 8619 22015
rect 10517 21981 10551 22015
rect 12541 21981 12575 22015
rect 15209 21981 15243 22015
rect 19533 21981 19567 22015
rect 20361 21981 20395 22015
rect 23673 21981 23707 22015
rect 23765 21981 23799 22015
rect 25789 21981 25823 22015
rect 28825 21981 28859 22015
rect 31861 21981 31895 22015
rect 32229 21981 32263 22015
rect 32597 21981 32631 22015
rect 32873 21981 32907 22015
rect 34069 21981 34103 22015
rect 48605 21981 48639 22015
rect 49065 21981 49099 22015
rect 3433 21913 3467 21947
rect 14381 21913 14415 21947
rect 14933 21913 14967 21947
rect 17417 21913 17451 21947
rect 21281 21913 21315 21947
rect 22661 21913 22695 21947
rect 24961 21913 24995 21947
rect 25053 21913 25087 21947
rect 29285 21913 29319 21947
rect 31401 21913 31435 21947
rect 3617 21845 3651 21879
rect 6101 21845 6135 21879
rect 9321 21845 9355 21879
rect 9689 21845 9723 21879
rect 9781 21845 9815 21879
rect 14473 21845 14507 21879
rect 18889 21845 18923 21879
rect 19625 21845 19659 21879
rect 22109 21845 22143 21879
rect 22385 21845 22419 21879
rect 27997 21845 28031 21879
rect 28641 21845 28675 21879
rect 30113 21845 30147 21879
rect 30481 21845 30515 21879
rect 31493 21845 31527 21879
rect 32137 21845 32171 21879
rect 33701 21845 33735 21879
rect 48421 21845 48455 21879
rect 49249 21845 49283 21879
rect 6469 21641 6503 21675
rect 9413 21641 9447 21675
rect 10977 21641 11011 21675
rect 11161 21641 11195 21675
rect 16037 21641 16071 21675
rect 20821 21641 20855 21675
rect 21005 21641 21039 21675
rect 23029 21641 23063 21675
rect 25973 21641 26007 21675
rect 27261 21641 27295 21675
rect 27721 21641 27755 21675
rect 31125 21641 31159 21675
rect 33241 21641 33275 21675
rect 4353 21573 4387 21607
rect 7941 21573 7975 21607
rect 15945 21573 15979 21607
rect 23673 21573 23707 21607
rect 26065 21573 26099 21607
rect 1777 21505 1811 21539
rect 3433 21505 3467 21539
rect 5641 21505 5675 21539
rect 7021 21505 7055 21539
rect 10241 21505 10275 21539
rect 12173 21505 12207 21539
rect 12265 21505 12299 21539
rect 13093 21505 13127 21539
rect 16865 21505 16899 21539
rect 21281 21505 21315 21539
rect 22385 21505 22419 21539
rect 23397 21505 23431 21539
rect 27629 21505 27663 21539
rect 31033 21505 31067 21539
rect 31677 21505 31711 21539
rect 32413 21505 32447 21539
rect 32873 21505 32907 21539
rect 47961 21505 47995 21539
rect 2053 21437 2087 21471
rect 5733 21437 5767 21471
rect 5917 21437 5951 21471
rect 7665 21437 7699 21471
rect 10333 21437 10367 21471
rect 10517 21437 10551 21471
rect 12357 21437 12391 21471
rect 13369 21437 13403 21471
rect 16221 21437 16255 21471
rect 17325 21437 17359 21471
rect 18705 21437 18739 21471
rect 18981 21437 19015 21471
rect 22477 21437 22511 21471
rect 22661 21437 22695 21471
rect 25145 21437 25179 21471
rect 26249 21437 26283 21471
rect 26709 21437 26743 21471
rect 27813 21437 27847 21471
rect 28457 21437 28491 21471
rect 28733 21437 28767 21471
rect 31217 21437 31251 21471
rect 33609 21437 33643 21471
rect 49157 21437 49191 21471
rect 7205 21369 7239 21403
rect 15577 21369 15611 21403
rect 22017 21369 22051 21403
rect 25605 21369 25639 21403
rect 33057 21369 33091 21403
rect 5273 21301 5307 21335
rect 6561 21301 6595 21335
rect 9689 21301 9723 21335
rect 9873 21301 9907 21335
rect 11345 21301 11379 21335
rect 11805 21301 11839 21335
rect 14841 21301 14875 21335
rect 15301 21301 15335 21335
rect 20453 21301 20487 21335
rect 30205 21301 30239 21335
rect 30665 21301 30699 21335
rect 31861 21301 31895 21335
rect 32505 21301 32539 21335
rect 33425 21301 33459 21335
rect 47685 21301 47719 21335
rect 3433 21097 3467 21131
rect 10977 21097 11011 21131
rect 27813 21097 27847 21131
rect 32505 21097 32539 21131
rect 49433 21097 49467 21131
rect 5089 21029 5123 21063
rect 7849 21029 7883 21063
rect 22109 21029 22143 21063
rect 4261 20961 4295 20995
rect 5733 20961 5767 20995
rect 8309 20961 8343 20995
rect 8493 20961 8527 20995
rect 9597 20961 9631 20995
rect 12541 20961 12575 20995
rect 14289 20961 14323 20995
rect 15117 20961 15151 20995
rect 16221 20961 16255 20995
rect 16405 20961 16439 20995
rect 17601 20961 17635 20995
rect 18797 20961 18831 20995
rect 19717 20961 19751 20995
rect 21557 20961 21591 20995
rect 22753 20961 22787 20995
rect 23765 20961 23799 20995
rect 23857 20961 23891 20995
rect 25237 20961 25271 20995
rect 25697 20961 25731 20995
rect 26065 20961 26099 20995
rect 26341 20961 26375 20995
rect 28549 20961 28583 20995
rect 30021 20961 30055 20995
rect 1777 20893 1811 20927
rect 3985 20893 4019 20927
rect 5457 20893 5491 20927
rect 7757 20893 7791 20927
rect 8217 20893 8251 20927
rect 9137 20893 9171 20927
rect 11989 20893 12023 20927
rect 17417 20893 17451 20927
rect 18521 20893 18555 20927
rect 19441 20893 19475 20927
rect 21833 20893 21867 20927
rect 28273 20893 28307 20927
rect 29745 20893 29779 20927
rect 31125 20893 31159 20927
rect 32689 20893 32723 20927
rect 32965 20893 32999 20927
rect 2789 20825 2823 20859
rect 3617 20825 3651 20859
rect 11345 20825 11379 20859
rect 13737 20825 13771 20859
rect 15025 20825 15059 20859
rect 25053 20825 25087 20859
rect 31861 20825 31895 20859
rect 7205 20757 7239 20791
rect 7573 20757 7607 20791
rect 11437 20757 11471 20791
rect 13921 20757 13955 20791
rect 14565 20757 14599 20791
rect 14933 20757 14967 20791
rect 15761 20757 15795 20791
rect 16129 20757 16163 20791
rect 16957 20757 16991 20791
rect 17325 20757 17359 20791
rect 18153 20757 18187 20791
rect 18613 20757 18647 20791
rect 21189 20757 21223 20791
rect 22477 20757 22511 20791
rect 22569 20757 22603 20791
rect 23305 20757 23339 20791
rect 23673 20757 23707 20791
rect 24685 20757 24719 20791
rect 25145 20757 25179 20791
rect 31217 20757 31251 20791
rect 31953 20757 31987 20791
rect 5641 20553 5675 20587
rect 13001 20553 13035 20587
rect 16129 20553 16163 20587
rect 17509 20553 17543 20587
rect 18245 20553 18279 20587
rect 18521 20553 18555 20587
rect 18889 20553 18923 20587
rect 23397 20553 23431 20587
rect 24041 20553 24075 20587
rect 26525 20553 26559 20587
rect 27629 20553 27663 20587
rect 30941 20553 30975 20587
rect 8769 20485 8803 20519
rect 11805 20485 11839 20519
rect 22753 20485 22787 20519
rect 31585 20485 31619 20519
rect 32137 20485 32171 20519
rect 1777 20417 1811 20451
rect 3433 20417 3467 20451
rect 6561 20417 6595 20451
rect 12909 20417 12943 20451
rect 13737 20417 13771 20451
rect 16037 20417 16071 20451
rect 17417 20417 17451 20451
rect 18981 20417 19015 20451
rect 19717 20417 19751 20451
rect 22017 20417 22051 20451
rect 24317 20417 24351 20451
rect 26801 20417 26835 20451
rect 27537 20417 27571 20451
rect 31033 20417 31067 20451
rect 2789 20349 2823 20383
rect 3893 20349 3927 20383
rect 5733 20349 5767 20383
rect 5825 20349 5859 20383
rect 7021 20349 7055 20383
rect 9413 20349 9447 20383
rect 9689 20349 9723 20383
rect 12449 20349 12483 20383
rect 13185 20349 13219 20383
rect 14013 20349 14047 20383
rect 16865 20349 16899 20383
rect 17693 20349 17727 20383
rect 19073 20349 19107 20383
rect 19993 20349 20027 20383
rect 24593 20349 24627 20383
rect 26065 20349 26099 20383
rect 27721 20349 27755 20383
rect 28365 20349 28399 20383
rect 28641 20349 28675 20383
rect 31125 20349 31159 20383
rect 31769 20349 31803 20383
rect 17049 20281 17083 20315
rect 27169 20281 27203 20315
rect 5273 20213 5307 20247
rect 8401 20213 8435 20247
rect 8861 20213 8895 20247
rect 11161 20213 11195 20247
rect 11897 20213 11931 20247
rect 12541 20213 12575 20247
rect 15485 20213 15519 20247
rect 16681 20213 16715 20247
rect 21465 20213 21499 20247
rect 26433 20213 26467 20247
rect 30113 20213 30147 20247
rect 30573 20213 30607 20247
rect 3341 20009 3375 20043
rect 3801 20009 3835 20043
rect 3985 20009 4019 20043
rect 4169 20009 4203 20043
rect 6285 20009 6319 20043
rect 8493 20009 8527 20043
rect 10885 20009 10919 20043
rect 11345 20009 11379 20043
rect 11437 20009 11471 20043
rect 13001 20009 13035 20043
rect 14289 20009 14323 20043
rect 18705 20009 18739 20043
rect 30757 20009 30791 20043
rect 16773 19941 16807 19975
rect 17233 19941 17267 19975
rect 24685 19941 24719 19975
rect 29745 19941 29779 19975
rect 2789 19873 2823 19907
rect 4537 19873 4571 19907
rect 6745 19873 6779 19907
rect 9137 19873 9171 19907
rect 12357 19873 12391 19907
rect 13645 19873 13679 19907
rect 14841 19873 14875 19907
rect 16957 19873 16991 19907
rect 17693 19873 17727 19907
rect 17877 19873 17911 19907
rect 20545 19873 20579 19907
rect 23857 19873 23891 19907
rect 25145 19873 25179 19907
rect 25237 19873 25271 19907
rect 28641 19873 28675 19907
rect 31309 19873 31343 19907
rect 1777 19805 1811 19839
rect 12173 19805 12207 19839
rect 12265 19805 12299 19839
rect 14565 19805 14599 19839
rect 17601 19805 17635 19839
rect 18889 19805 18923 19839
rect 20269 19805 20303 19839
rect 22569 19805 22603 19839
rect 23765 19805 23799 19839
rect 25881 19805 25915 19839
rect 27905 19805 27939 19839
rect 28365 19805 28399 19839
rect 29929 19805 29963 19839
rect 30205 19805 30239 19839
rect 31217 19805 31251 19839
rect 3617 19737 3651 19771
rect 4813 19737 4847 19771
rect 7021 19737 7055 19771
rect 9413 19737 9447 19771
rect 13461 19737 13495 19771
rect 19625 19737 19659 19771
rect 22753 19737 22787 19771
rect 26157 19737 26191 19771
rect 11805 19669 11839 19703
rect 13369 19669 13403 19703
rect 16313 19669 16347 19703
rect 18429 19669 18463 19703
rect 19717 19669 19751 19703
rect 22017 19669 22051 19703
rect 23305 19669 23339 19703
rect 23673 19669 23707 19703
rect 25053 19669 25087 19703
rect 27629 19669 27663 19703
rect 30389 19669 30423 19703
rect 31125 19669 31159 19703
rect 5273 19465 5307 19499
rect 5733 19465 5767 19499
rect 10425 19465 10459 19499
rect 10885 19465 10919 19499
rect 14841 19465 14875 19499
rect 17233 19465 17267 19499
rect 17877 19465 17911 19499
rect 19073 19465 19107 19499
rect 21465 19465 21499 19499
rect 22385 19465 22419 19499
rect 23673 19465 23707 19499
rect 26433 19465 26467 19499
rect 27721 19465 27755 19499
rect 30481 19465 30515 19499
rect 4353 19397 4387 19431
rect 5641 19397 5675 19431
rect 9321 19397 9355 19431
rect 18337 19397 18371 19431
rect 22477 19397 22511 19431
rect 24133 19397 24167 19431
rect 27261 19397 27295 19431
rect 28549 19397 28583 19431
rect 1777 19329 1811 19363
rect 2789 19329 2823 19363
rect 3617 19329 3651 19363
rect 6653 19329 6687 19363
rect 7481 19329 7515 19363
rect 8585 19329 8619 19363
rect 10333 19329 10367 19363
rect 10793 19329 10827 19363
rect 11713 19329 11747 19363
rect 14749 19329 14783 19363
rect 15669 19329 15703 19363
rect 17417 19329 17451 19363
rect 18245 19329 18279 19363
rect 19257 19329 19291 19363
rect 24041 19329 24075 19363
rect 24961 19329 24995 19363
rect 30665 19329 30699 19363
rect 31125 19329 31159 19363
rect 5917 19261 5951 19295
rect 10977 19261 11011 19295
rect 11989 19261 12023 19295
rect 13461 19261 13495 19295
rect 13921 19261 13955 19295
rect 14933 19261 14967 19295
rect 16957 19261 16991 19295
rect 18429 19261 18463 19295
rect 19717 19261 19751 19295
rect 22661 19261 22695 19295
rect 24317 19261 24351 19295
rect 25789 19261 25823 19295
rect 26985 19261 27019 19295
rect 28273 19261 28307 19295
rect 30941 19261 30975 19295
rect 10149 19193 10183 19227
rect 15853 19193 15887 19227
rect 23305 19193 23339 19227
rect 27445 19193 27479 19227
rect 14105 19125 14139 19159
rect 14381 19125 14415 19159
rect 16221 19125 16255 19159
rect 16405 19125 16439 19159
rect 16773 19125 16807 19159
rect 17693 19125 17727 19159
rect 19980 19125 20014 19159
rect 22017 19125 22051 19159
rect 23121 19125 23155 19159
rect 27905 19125 27939 19159
rect 30021 19125 30055 19159
rect 3893 18921 3927 18955
rect 9413 18921 9447 18955
rect 11621 18921 11655 18955
rect 22937 18921 22971 18955
rect 27169 18921 27203 18955
rect 14197 18853 14231 18887
rect 18153 18853 18187 18887
rect 25145 18853 25179 18887
rect 3985 18785 4019 18819
rect 6837 18785 6871 18819
rect 8585 18785 8619 18819
rect 9045 18785 9079 18819
rect 9873 18785 9907 18819
rect 9965 18785 9999 18819
rect 12173 18785 12207 18819
rect 15209 18785 15243 18819
rect 17509 18785 17543 18819
rect 18705 18785 18739 18819
rect 20361 18785 20395 18819
rect 21189 18785 21223 18819
rect 21465 18785 21499 18819
rect 24593 18785 24627 18819
rect 25421 18785 25455 18819
rect 27629 18785 27663 18819
rect 30205 18785 30239 18819
rect 30297 18785 30331 18819
rect 30849 18785 30883 18819
rect 1777 18717 1811 18751
rect 4629 18717 4663 18751
rect 10609 18717 10643 18751
rect 14565 18717 14599 18751
rect 18613 18717 18647 18751
rect 19625 18717 19659 18751
rect 23581 18717 23615 18751
rect 24041 18717 24075 18751
rect 27905 18717 27939 18751
rect 2789 18649 2823 18683
rect 3617 18649 3651 18683
rect 4905 18649 4939 18683
rect 7113 18649 7147 18683
rect 10977 18649 11011 18683
rect 12817 18649 12851 18683
rect 13553 18649 13587 18683
rect 15485 18649 15519 18683
rect 25697 18649 25731 18683
rect 3341 18581 3375 18615
rect 6377 18581 6411 18615
rect 9781 18581 9815 18615
rect 11069 18581 11103 18615
rect 11989 18581 12023 18615
rect 12081 18581 12115 18615
rect 14657 18581 14691 18615
rect 16957 18581 16991 18615
rect 18521 18581 18555 18615
rect 19349 18581 19383 18615
rect 20821 18581 20855 18615
rect 23397 18581 23431 18615
rect 24133 18581 24167 18615
rect 29745 18581 29779 18615
rect 30113 18581 30147 18615
rect 9781 18377 9815 18411
rect 10425 18377 10459 18411
rect 12357 18377 12391 18411
rect 15393 18377 15427 18411
rect 17325 18377 17359 18411
rect 19901 18377 19935 18411
rect 20729 18377 20763 18411
rect 24869 18377 24903 18411
rect 26801 18377 26835 18411
rect 27169 18377 27203 18411
rect 30757 18377 30791 18411
rect 31493 18377 31527 18411
rect 9965 18309 9999 18343
rect 14473 18309 14507 18343
rect 16221 18309 16255 18343
rect 18153 18309 18187 18343
rect 21097 18309 21131 18343
rect 25329 18309 25363 18343
rect 26065 18309 26099 18343
rect 28365 18309 28399 18343
rect 1777 18241 1811 18275
rect 3617 18241 3651 18275
rect 5641 18241 5675 18275
rect 5733 18241 5767 18275
rect 6745 18241 6779 18275
rect 8493 18241 8527 18275
rect 10793 18241 10827 18275
rect 12449 18241 12483 18275
rect 13645 18241 13679 18275
rect 17233 18241 17267 18275
rect 18337 18241 18371 18275
rect 19993 18241 20027 18275
rect 22017 18241 22051 18275
rect 26525 18241 26559 18275
rect 28089 18241 28123 18275
rect 30665 18241 30699 18275
rect 31309 18241 31343 18275
rect 2053 18173 2087 18207
rect 3893 18173 3927 18207
rect 5917 18173 5951 18207
rect 7297 18173 7331 18207
rect 9229 18173 9263 18207
rect 10885 18173 10919 18207
rect 11069 18173 11103 18207
rect 12633 18173 12667 18207
rect 13185 18173 13219 18207
rect 15485 18173 15519 18207
rect 15669 18173 15703 18207
rect 17509 18173 17543 18207
rect 18889 18173 18923 18207
rect 20085 18173 20119 18207
rect 21189 18173 21223 18207
rect 21281 18173 21315 18207
rect 22569 18173 22603 18207
rect 22845 18173 22879 18207
rect 23121 18173 23155 18207
rect 23397 18173 23431 18207
rect 30849 18173 30883 18207
rect 11989 18105 12023 18139
rect 15025 18105 15059 18139
rect 19533 18105 19567 18139
rect 30297 18105 30331 18139
rect 5273 18037 5307 18071
rect 10057 18037 10091 18071
rect 11713 18037 11747 18071
rect 13369 18037 13403 18071
rect 16037 18037 16071 18071
rect 16405 18037 16439 18071
rect 16865 18037 16899 18071
rect 29837 18037 29871 18071
rect 3617 17833 3651 17867
rect 10609 17833 10643 17867
rect 13737 17833 13771 17867
rect 21925 17833 21959 17867
rect 30941 17833 30975 17867
rect 4445 17765 4479 17799
rect 6653 17765 6687 17799
rect 7849 17765 7883 17799
rect 20729 17765 20763 17799
rect 26617 17765 26651 17799
rect 29745 17765 29779 17799
rect 7389 17697 7423 17731
rect 8401 17697 8435 17731
rect 9873 17697 9907 17731
rect 11161 17697 11195 17731
rect 12265 17697 12299 17731
rect 16313 17697 16347 17731
rect 16589 17697 16623 17731
rect 19441 17697 19475 17731
rect 19717 17697 19751 17731
rect 21281 17697 21315 17731
rect 24869 17697 24903 17731
rect 27077 17697 27111 17731
rect 28825 17697 28859 17731
rect 29193 17697 29227 17731
rect 30297 17697 30331 17731
rect 31493 17697 31527 17731
rect 1777 17629 1811 17663
rect 3801 17629 3835 17663
rect 4905 17629 4939 17663
rect 8217 17629 8251 17663
rect 9137 17629 9171 17663
rect 11069 17629 11103 17663
rect 11713 17629 11747 17663
rect 11989 17629 12023 17663
rect 21097 17629 21131 17663
rect 22293 17629 22327 17663
rect 31309 17629 31343 17663
rect 31401 17629 31435 17663
rect 2513 17561 2547 17595
rect 3433 17561 3467 17595
rect 4261 17561 4295 17595
rect 5181 17561 5215 17595
rect 7205 17561 7239 17595
rect 8309 17561 8343 17595
rect 10977 17561 11011 17595
rect 14381 17561 14415 17595
rect 18337 17561 18371 17595
rect 21189 17561 21223 17595
rect 22569 17561 22603 17595
rect 25145 17561 25179 17595
rect 27353 17561 27387 17595
rect 30113 17561 30147 17595
rect 14473 17493 14507 17527
rect 14933 17493 14967 17527
rect 15117 17493 15151 17527
rect 15393 17493 15427 17527
rect 16037 17493 16071 17527
rect 18061 17493 18095 17527
rect 18705 17493 18739 17527
rect 21741 17493 21775 17527
rect 24041 17493 24075 17527
rect 24409 17493 24443 17527
rect 30205 17493 30239 17527
rect 4905 17289 4939 17323
rect 5089 17289 5123 17323
rect 5641 17289 5675 17323
rect 6837 17289 6871 17323
rect 8033 17289 8067 17323
rect 11897 17289 11931 17323
rect 12541 17289 12575 17323
rect 13737 17289 13771 17323
rect 16129 17289 16163 17323
rect 22017 17289 22051 17323
rect 22385 17289 22419 17323
rect 29837 17289 29871 17323
rect 30573 17289 30607 17323
rect 30849 17289 30883 17323
rect 30941 17289 30975 17323
rect 4353 17221 4387 17255
rect 7205 17221 7239 17255
rect 9965 17221 9999 17255
rect 10793 17221 10827 17255
rect 14197 17221 14231 17255
rect 14749 17221 14783 17255
rect 18429 17221 18463 17255
rect 24961 17221 24995 17255
rect 26801 17221 26835 17255
rect 1777 17153 1811 17187
rect 3617 17153 3651 17187
rect 8401 17153 8435 17187
rect 9873 17153 9907 17187
rect 11805 17153 11839 17187
rect 12909 17153 12943 17187
rect 13001 17153 13035 17187
rect 14105 17153 14139 17187
rect 14933 17153 14967 17187
rect 15669 17153 15703 17187
rect 16313 17153 16347 17187
rect 17233 17153 17267 17187
rect 21097 17153 21131 17187
rect 23673 17153 23707 17187
rect 24409 17153 24443 17187
rect 24685 17153 24719 17187
rect 27813 17153 27847 17187
rect 2053 17085 2087 17119
rect 5733 17085 5767 17119
rect 5917 17085 5951 17119
rect 6469 17085 6503 17119
rect 7297 17085 7331 17119
rect 7481 17085 7515 17119
rect 8493 17085 8527 17119
rect 8677 17085 8711 17119
rect 10057 17085 10091 17119
rect 13093 17085 13127 17119
rect 14381 17085 14415 17119
rect 17325 17085 17359 17119
rect 17417 17085 17451 17119
rect 18153 17085 18187 17119
rect 21189 17085 21223 17119
rect 21373 17085 21407 17119
rect 22477 17085 22511 17119
rect 22569 17085 22603 17119
rect 23765 17085 23799 17119
rect 23857 17085 23891 17119
rect 26433 17085 26467 17119
rect 27169 17085 27203 17119
rect 28089 17085 28123 17119
rect 5273 17017 5307 17051
rect 9505 17017 9539 17051
rect 15485 17017 15519 17051
rect 20361 17017 20395 17051
rect 9137 16949 9171 16983
rect 10885 16949 10919 16983
rect 11345 16949 11379 16983
rect 15209 16949 15243 16983
rect 16865 16949 16899 16983
rect 19901 16949 19935 16983
rect 20177 16949 20211 16983
rect 20729 16949 20763 16983
rect 23305 16949 23339 16983
rect 29561 16949 29595 16983
rect 3433 16677 3467 16711
rect 3617 16677 3651 16711
rect 6101 16677 6135 16711
rect 9413 16677 9447 16711
rect 9781 16677 9815 16711
rect 12449 16677 12483 16711
rect 13001 16677 13035 16711
rect 4537 16609 4571 16643
rect 7113 16609 7147 16643
rect 7297 16609 7331 16643
rect 8493 16609 8527 16643
rect 10701 16609 10735 16643
rect 11713 16609 11747 16643
rect 11897 16609 11931 16643
rect 12725 16609 12759 16643
rect 13461 16609 13495 16643
rect 13645 16609 13679 16643
rect 15485 16609 15519 16643
rect 15669 16609 15703 16643
rect 16773 16609 16807 16643
rect 19717 16609 19751 16643
rect 22477 16609 22511 16643
rect 22569 16609 22603 16643
rect 23765 16609 23799 16643
rect 25329 16609 25363 16643
rect 25973 16609 26007 16643
rect 27077 16609 27111 16643
rect 27169 16609 27203 16643
rect 28457 16609 28491 16643
rect 1777 16541 1811 16575
rect 3985 16541 4019 16575
rect 10425 16541 10459 16575
rect 10517 16541 10551 16575
rect 14565 16541 14599 16575
rect 15393 16541 15427 16575
rect 16221 16541 16255 16575
rect 17601 16541 17635 16575
rect 18245 16541 18279 16575
rect 19441 16541 19475 16575
rect 22385 16541 22419 16575
rect 23581 16541 23615 16575
rect 28181 16541 28215 16575
rect 28273 16541 28307 16575
rect 2513 16473 2547 16507
rect 5917 16473 5951 16507
rect 7021 16473 7055 16507
rect 8217 16473 8251 16507
rect 9229 16473 9263 16507
rect 13369 16473 13403 16507
rect 21465 16473 21499 16507
rect 26985 16473 27019 16507
rect 6653 16405 6687 16439
rect 7849 16405 7883 16439
rect 8309 16405 8343 16439
rect 10057 16405 10091 16439
rect 11253 16405 11287 16439
rect 11621 16405 11655 16439
rect 12265 16405 12299 16439
rect 14381 16405 14415 16439
rect 15025 16405 15059 16439
rect 16037 16405 16071 16439
rect 16405 16405 16439 16439
rect 17417 16405 17451 16439
rect 18061 16405 18095 16439
rect 18705 16405 18739 16439
rect 22017 16405 22051 16439
rect 23213 16405 23247 16439
rect 23673 16405 23707 16439
rect 24685 16405 24719 16439
rect 25053 16405 25087 16439
rect 25145 16405 25179 16439
rect 25697 16405 25731 16439
rect 26617 16405 26651 16439
rect 27813 16405 27847 16439
rect 7297 16201 7331 16235
rect 10241 16201 10275 16235
rect 10609 16201 10643 16235
rect 11621 16201 11655 16235
rect 13737 16201 13771 16235
rect 16957 16201 16991 16235
rect 17141 16201 17175 16235
rect 17417 16201 17451 16235
rect 17877 16201 17911 16235
rect 19717 16201 19751 16235
rect 20545 16201 20579 16235
rect 26617 16201 26651 16235
rect 26985 16201 27019 16235
rect 27721 16201 27755 16235
rect 4353 16133 4387 16167
rect 5733 16133 5767 16167
rect 14657 16133 14691 16167
rect 24409 16133 24443 16167
rect 24593 16133 24627 16167
rect 1777 16065 1811 16099
rect 3525 16065 3559 16099
rect 5641 16065 5675 16099
rect 7665 16065 7699 16099
rect 8493 16065 8527 16099
rect 11161 16065 11195 16099
rect 11989 16065 12023 16099
rect 14749 16065 14783 16099
rect 16313 16065 16347 16099
rect 17785 16065 17819 16099
rect 18613 16065 18647 16099
rect 18889 16065 18923 16099
rect 20453 16065 20487 16099
rect 21465 16065 21499 16099
rect 23673 16065 23707 16099
rect 23765 16065 23799 16099
rect 24869 16065 24903 16099
rect 2053 15997 2087 16031
rect 5917 15997 5951 16031
rect 6653 15997 6687 16031
rect 7757 15997 7791 16031
rect 7941 15997 7975 16031
rect 8769 15997 8803 16031
rect 12265 15997 12299 16031
rect 14841 15997 14875 16031
rect 15485 15997 15519 16031
rect 17969 15997 18003 16031
rect 20729 15997 20763 16031
rect 22017 15997 22051 16031
rect 22293 15997 22327 16031
rect 23949 15997 23983 16031
rect 25145 15997 25179 16031
rect 10977 15929 11011 15963
rect 20085 15929 20119 15963
rect 5273 15861 5307 15895
rect 14289 15861 14323 15895
rect 16129 15861 16163 15895
rect 16681 15861 16715 15895
rect 21281 15861 21315 15895
rect 23305 15861 23339 15895
rect 7849 15657 7883 15691
rect 9321 15657 9355 15691
rect 13553 15657 13587 15691
rect 15853 15657 15887 15691
rect 19901 15657 19935 15691
rect 22477 15657 22511 15691
rect 24501 15657 24535 15691
rect 7481 15589 7515 15623
rect 22845 15589 22879 15623
rect 2053 15521 2087 15555
rect 4445 15521 4479 15555
rect 4629 15521 4663 15555
rect 5641 15521 5675 15555
rect 5825 15521 5859 15555
rect 6837 15521 6871 15555
rect 6929 15521 6963 15555
rect 8493 15521 8527 15555
rect 10241 15521 10275 15555
rect 11437 15521 11471 15555
rect 12725 15521 12759 15555
rect 14933 15521 14967 15555
rect 15117 15521 15151 15555
rect 16497 15521 16531 15555
rect 20269 15521 20303 15555
rect 25789 15521 25823 15555
rect 1777 15453 1811 15487
rect 11345 15453 11379 15487
rect 13737 15453 13771 15487
rect 14841 15453 14875 15487
rect 17049 15453 17083 15487
rect 19625 15453 19659 15487
rect 23121 15453 23155 15487
rect 3341 15385 3375 15419
rect 5549 15385 5583 15419
rect 6745 15385 6779 15419
rect 8217 15385 8251 15419
rect 9229 15385 9263 15419
rect 12449 15385 12483 15419
rect 13277 15385 13311 15419
rect 16221 15385 16255 15419
rect 17325 15385 17359 15419
rect 20545 15385 20579 15419
rect 23949 15385 23983 15419
rect 25697 15385 25731 15419
rect 3617 15317 3651 15351
rect 3985 15317 4019 15351
rect 4353 15317 4387 15351
rect 5181 15317 5215 15351
rect 6377 15317 6411 15351
rect 8309 15317 8343 15351
rect 9781 15317 9815 15351
rect 9873 15317 9907 15351
rect 10885 15317 10919 15351
rect 11253 15317 11287 15351
rect 12081 15317 12115 15351
rect 12541 15317 12575 15351
rect 14105 15317 14139 15351
rect 14473 15317 14507 15351
rect 15485 15317 15519 15351
rect 16313 15317 16347 15351
rect 18797 15317 18831 15351
rect 19441 15317 19475 15351
rect 22017 15317 22051 15351
rect 22385 15317 22419 15351
rect 25237 15317 25271 15351
rect 25605 15317 25639 15351
rect 26249 15317 26283 15351
rect 26525 15317 26559 15351
rect 3525 15113 3559 15147
rect 6745 15113 6779 15147
rect 7665 15113 7699 15147
rect 9597 15113 9631 15147
rect 18429 15113 18463 15147
rect 23765 15113 23799 15147
rect 27077 15113 27111 15147
rect 7757 15045 7791 15079
rect 9689 15045 9723 15079
rect 10793 15045 10827 15079
rect 16773 15045 16807 15079
rect 20913 15045 20947 15079
rect 22293 15045 22327 15079
rect 25145 15045 25179 15079
rect 1777 14977 1811 15011
rect 3709 14977 3743 15011
rect 4169 14977 4203 15011
rect 6653 14977 6687 15011
rect 8585 14977 8619 15011
rect 10885 14977 10919 15011
rect 11713 14977 11747 15011
rect 11989 14977 12023 15011
rect 13369 14977 13403 15011
rect 13461 14977 13495 15011
rect 14013 14977 14047 15011
rect 17141 14977 17175 15011
rect 19165 14977 19199 15011
rect 20085 14977 20119 15011
rect 22017 14977 22051 15011
rect 24869 14977 24903 15011
rect 2053 14909 2087 14943
rect 4445 14909 4479 14943
rect 7849 14909 7883 14943
rect 9873 14909 9907 14943
rect 10977 14909 11011 14943
rect 13553 14909 13587 14943
rect 14565 14909 14599 14943
rect 14841 14909 14875 14943
rect 20177 14909 20211 14943
rect 20361 14909 20395 14943
rect 10425 14841 10459 14875
rect 13001 14841 13035 14875
rect 19717 14841 19751 14875
rect 5917 14773 5951 14807
rect 7297 14773 7331 14807
rect 8677 14773 8711 14807
rect 9229 14773 9263 14807
rect 14197 14773 14231 14807
rect 16313 14773 16347 14807
rect 19349 14773 19383 14807
rect 20729 14773 20763 14807
rect 24041 14773 24075 14807
rect 24225 14773 24259 14807
rect 26617 14773 26651 14807
rect 3985 14569 4019 14603
rect 9413 14569 9447 14603
rect 11621 14569 11655 14603
rect 13737 14569 13771 14603
rect 14381 14569 14415 14603
rect 18613 14569 18647 14603
rect 19441 14569 19475 14603
rect 21741 14501 21775 14535
rect 24041 14501 24075 14535
rect 26893 14501 26927 14535
rect 2053 14433 2087 14467
rect 4813 14433 4847 14467
rect 7205 14433 7239 14467
rect 8309 14433 8343 14467
rect 8493 14433 8527 14467
rect 10057 14433 10091 14467
rect 11161 14433 11195 14467
rect 12265 14433 12299 14467
rect 14657 14433 14691 14467
rect 14933 14433 14967 14467
rect 16865 14433 16899 14467
rect 21097 14433 21131 14467
rect 22293 14433 22327 14467
rect 25145 14433 25179 14467
rect 26249 14433 26283 14467
rect 26341 14433 26375 14467
rect 1777 14365 1811 14399
rect 5457 14365 5491 14399
rect 9873 14365 9907 14399
rect 11989 14365 12023 14399
rect 18889 14365 18923 14399
rect 19625 14365 19659 14399
rect 20913 14365 20947 14399
rect 21557 14365 21591 14399
rect 4629 14297 4663 14331
rect 5733 14297 5767 14331
rect 10977 14297 11011 14331
rect 14105 14297 14139 14331
rect 17141 14297 17175 14331
rect 22569 14297 22603 14331
rect 25053 14297 25087 14331
rect 26157 14297 26191 14331
rect 26985 14297 27019 14331
rect 3341 14229 3375 14263
rect 3525 14229 3559 14263
rect 4261 14229 4295 14263
rect 4721 14229 4755 14263
rect 7849 14229 7883 14263
rect 8217 14229 8251 14263
rect 9045 14229 9079 14263
rect 9781 14229 9815 14263
rect 10609 14229 10643 14263
rect 11069 14229 11103 14263
rect 16405 14229 16439 14263
rect 20545 14229 20579 14263
rect 21005 14229 21039 14263
rect 24593 14229 24627 14263
rect 24961 14229 24995 14263
rect 25789 14229 25823 14263
rect 3433 14025 3467 14059
rect 4077 14025 4111 14059
rect 5641 14025 5675 14059
rect 6561 14025 6595 14059
rect 6929 14025 6963 14059
rect 7297 14025 7331 14059
rect 8125 14025 8159 14059
rect 11989 14025 12023 14059
rect 12357 14025 12391 14059
rect 13185 14025 13219 14059
rect 14749 14025 14783 14059
rect 14841 14025 14875 14059
rect 15577 14025 15611 14059
rect 18889 14025 18923 14059
rect 19441 14025 19475 14059
rect 20085 14025 20119 14059
rect 23397 14025 23431 14059
rect 24961 14025 24995 14059
rect 4537 13957 4571 13991
rect 5733 13957 5767 13991
rect 6469 13957 6503 13991
rect 8493 13957 8527 13991
rect 8585 13957 8619 13991
rect 11621 13957 11655 13991
rect 12449 13957 12483 13991
rect 13645 13957 13679 13991
rect 21833 13957 21867 13991
rect 22661 13957 22695 13991
rect 25053 13957 25087 13991
rect 25605 13957 25639 13991
rect 1777 13889 1811 13923
rect 3617 13889 3651 13923
rect 4445 13889 4479 13923
rect 7389 13889 7423 13923
rect 13553 13889 13587 13923
rect 15945 13889 15979 13923
rect 16037 13889 16071 13923
rect 19625 13889 19659 13923
rect 20453 13889 20487 13923
rect 20545 13889 20579 13923
rect 22569 13889 22603 13923
rect 23765 13889 23799 13923
rect 23857 13889 23891 13923
rect 25789 13889 25823 13923
rect 2053 13821 2087 13855
rect 4721 13821 4755 13855
rect 5917 13821 5951 13855
rect 7481 13821 7515 13855
rect 8677 13821 8711 13855
rect 9321 13821 9355 13855
rect 11069 13821 11103 13855
rect 12633 13821 12667 13855
rect 13829 13821 13863 13855
rect 14933 13821 14967 13855
rect 16221 13821 16255 13855
rect 17141 13821 17175 13855
rect 20729 13821 20763 13855
rect 22845 13821 22879 13855
rect 24041 13821 24075 13855
rect 25237 13821 25271 13855
rect 26157 13821 26191 13855
rect 14381 13753 14415 13787
rect 22201 13753 22235 13787
rect 25973 13753 26007 13787
rect 5273 13685 5307 13719
rect 9584 13685 9618 13719
rect 16681 13685 16715 13719
rect 17404 13685 17438 13719
rect 24593 13685 24627 13719
rect 3433 13481 3467 13515
rect 16037 13481 16071 13515
rect 18889 13481 18923 13515
rect 22109 13481 22143 13515
rect 22569 13481 22603 13515
rect 23949 13481 23983 13515
rect 24133 13481 24167 13515
rect 6377 13413 6411 13447
rect 11529 13413 11563 13447
rect 11713 13413 11747 13447
rect 13737 13413 13771 13447
rect 2053 13345 2087 13379
rect 4169 13345 4203 13379
rect 6745 13345 6779 13379
rect 8493 13345 8527 13379
rect 9137 13345 9171 13379
rect 9413 13345 9447 13379
rect 10885 13345 10919 13379
rect 10977 13345 11011 13379
rect 11989 13345 12023 13379
rect 14565 13345 14599 13379
rect 16497 13345 16531 13379
rect 17141 13345 17175 13379
rect 20361 13345 20395 13379
rect 23489 13345 23523 13379
rect 1777 13277 1811 13311
rect 6193 13277 6227 13311
rect 14289 13277 14323 13311
rect 4445 13209 4479 13243
rect 7021 13209 7055 13243
rect 10793 13209 10827 13243
rect 12265 13209 12299 13243
rect 17417 13209 17451 13243
rect 20637 13209 20671 13243
rect 23213 13209 23247 13243
rect 23305 13209 23339 13243
rect 24593 13209 24627 13243
rect 25421 13209 25455 13243
rect 3525 13141 3559 13175
rect 3893 13141 3927 13175
rect 5917 13141 5951 13175
rect 10425 13141 10459 13175
rect 19349 13141 19383 13175
rect 19441 13141 19475 13175
rect 22845 13141 22879 13175
rect 3617 12937 3651 12971
rect 4813 12937 4847 12971
rect 5733 12937 5767 12971
rect 6469 12937 6503 12971
rect 7297 12937 7331 12971
rect 12541 12937 12575 12971
rect 13737 12937 13771 12971
rect 16129 12937 16163 12971
rect 17785 12937 17819 12971
rect 18153 12937 18187 12971
rect 21097 12937 21131 12971
rect 24777 12937 24811 12971
rect 3525 12869 3559 12903
rect 4261 12869 4295 12903
rect 11345 12869 11379 12903
rect 11897 12869 11931 12903
rect 15669 12869 15703 12903
rect 18981 12869 19015 12903
rect 23305 12869 23339 12903
rect 1593 12801 1627 12835
rect 1869 12801 1903 12835
rect 2789 12801 2823 12835
rect 5641 12801 5675 12835
rect 7205 12801 7239 12835
rect 10701 12801 10735 12835
rect 12909 12801 12943 12835
rect 14105 12801 14139 12835
rect 14933 12801 14967 12835
rect 16313 12801 16347 12835
rect 18245 12801 18279 12835
rect 21189 12801 21223 12835
rect 23029 12801 23063 12835
rect 4445 12733 4479 12767
rect 5917 12733 5951 12767
rect 7389 12733 7423 12767
rect 8033 12733 8067 12767
rect 8309 12733 8343 12767
rect 10057 12733 10091 12767
rect 13001 12733 13035 12767
rect 13185 12733 13219 12767
rect 14197 12733 14231 12767
rect 14381 12733 14415 12767
rect 16865 12733 16899 12767
rect 18429 12733 18463 12767
rect 19809 12733 19843 12767
rect 21373 12733 21407 12767
rect 3157 12665 3191 12699
rect 10517 12665 10551 12699
rect 11161 12665 11195 12699
rect 25053 12665 25087 12699
rect 2973 12597 3007 12631
rect 4905 12597 4939 12631
rect 5273 12597 5307 12631
rect 6837 12597 6871 12631
rect 11621 12597 11655 12631
rect 20729 12597 20763 12631
rect 22201 12597 22235 12631
rect 3985 12393 4019 12427
rect 4629 12393 4663 12427
rect 7849 12393 7883 12427
rect 11805 12393 11839 12427
rect 13001 12393 13035 12427
rect 18061 12393 18095 12427
rect 18889 12393 18923 12427
rect 21833 12393 21867 12427
rect 3157 12325 3191 12359
rect 1869 12257 1903 12291
rect 4721 12257 4755 12291
rect 5365 12257 5399 12291
rect 7389 12257 7423 12291
rect 8401 12257 8435 12291
rect 9873 12257 9907 12291
rect 11253 12257 11287 12291
rect 12265 12257 12299 12291
rect 12357 12257 12391 12291
rect 13645 12257 13679 12291
rect 16589 12257 16623 12291
rect 19625 12257 19659 12291
rect 20085 12257 20119 12291
rect 22569 12257 22603 12291
rect 1593 12189 1627 12223
rect 2973 12189 3007 12223
rect 4169 12189 4203 12223
rect 8309 12189 8343 12223
rect 10977 12189 11011 12223
rect 11069 12189 11103 12223
rect 13461 12189 13495 12223
rect 15485 12189 15519 12223
rect 16313 12189 16347 12223
rect 22293 12189 22327 12223
rect 5641 12121 5675 12155
rect 9137 12121 9171 12155
rect 13369 12121 13403 12155
rect 14749 12121 14783 12155
rect 18521 12121 18555 12155
rect 20361 12121 20395 12155
rect 3525 12053 3559 12087
rect 8217 12053 8251 12087
rect 10609 12053 10643 12087
rect 12173 12053 12207 12087
rect 14105 12053 14139 12087
rect 14381 12053 14415 12087
rect 15945 12053 15979 12087
rect 18337 12053 18371 12087
rect 18981 12053 19015 12087
rect 19349 12053 19383 12087
rect 24041 12053 24075 12087
rect 24409 12053 24443 12087
rect 1501 11849 1535 11883
rect 1869 11849 1903 11883
rect 3433 11849 3467 11883
rect 4445 11849 4479 11883
rect 5273 11849 5307 11883
rect 5641 11849 5675 11883
rect 6745 11849 6779 11883
rect 12449 11849 12483 11883
rect 15577 11849 15611 11883
rect 17325 11849 17359 11883
rect 18153 11849 18187 11883
rect 1685 11781 1719 11815
rect 5733 11781 5767 11815
rect 11621 11781 11655 11815
rect 15209 11781 15243 11815
rect 18521 11781 18555 11815
rect 19165 11781 19199 11815
rect 22661 11781 22695 11815
rect 2421 11713 2455 11747
rect 4537 11713 4571 11747
rect 6377 11713 6411 11747
rect 7389 11713 7423 11747
rect 9597 11713 9631 11747
rect 12357 11713 12391 11747
rect 13185 11713 13219 11747
rect 15945 11713 15979 11747
rect 16037 11713 16071 11747
rect 2145 11645 2179 11679
rect 4721 11645 4755 11679
rect 5825 11645 5859 11679
rect 7665 11645 7699 11679
rect 10333 11645 10367 11679
rect 10977 11645 11011 11679
rect 12541 11645 12575 11679
rect 13461 11645 13495 11679
rect 16221 11645 16255 11679
rect 17417 11645 17451 11679
rect 17601 11645 17635 11679
rect 18613 11645 18647 11679
rect 18705 11645 18739 11679
rect 19717 11645 19751 11679
rect 19993 11645 20027 11679
rect 22385 11645 22419 11679
rect 24409 11577 24443 11611
rect 4077 11509 4111 11543
rect 9137 11509 9171 11543
rect 11989 11509 12023 11543
rect 14933 11509 14967 11543
rect 16957 11509 16991 11543
rect 19441 11509 19475 11543
rect 21465 11509 21499 11543
rect 21925 11509 21959 11543
rect 24133 11509 24167 11543
rect 3433 11305 3467 11339
rect 3617 11305 3651 11339
rect 6561 11305 6595 11339
rect 7849 11305 7883 11339
rect 13277 11305 13311 11339
rect 13553 11305 13587 11339
rect 16497 11305 16531 11339
rect 18889 11305 18923 11339
rect 22661 11305 22695 11339
rect 32045 11305 32079 11339
rect 1593 11237 1627 11271
rect 10333 11237 10367 11271
rect 14105 11237 14139 11271
rect 2237 11169 2271 11203
rect 4813 11169 4847 11203
rect 7021 11169 7055 11203
rect 8309 11169 8343 11203
rect 8493 11169 8527 11203
rect 9597 11169 9631 11203
rect 9689 11169 9723 11203
rect 10793 11169 10827 11203
rect 10977 11169 11011 11203
rect 11805 11169 11839 11203
rect 22937 11169 22971 11203
rect 29745 11169 29779 11203
rect 1777 11101 1811 11135
rect 2513 11101 2547 11135
rect 4077 11101 4111 11135
rect 8217 11101 8251 11135
rect 9505 11101 9539 11135
rect 11529 11101 11563 11135
rect 14749 11101 14783 11135
rect 17141 11101 17175 11135
rect 19533 11101 19567 11135
rect 20913 11101 20947 11135
rect 5089 11033 5123 11067
rect 7481 11033 7515 11067
rect 10701 11033 10735 11067
rect 15025 11033 15059 11067
rect 17417 11033 17451 11067
rect 20269 11033 20303 11067
rect 21189 11033 21223 11067
rect 30021 11033 30055 11067
rect 31769 11033 31803 11067
rect 4169 10965 4203 10999
rect 9137 10965 9171 10999
rect 13829 10965 13863 10999
rect 16773 10965 16807 10999
rect 1501 10761 1535 10795
rect 4629 10761 4663 10795
rect 5825 10761 5859 10795
rect 9965 10761 9999 10795
rect 10793 10761 10827 10795
rect 14841 10761 14875 10795
rect 19257 10761 19291 10795
rect 4813 10693 4847 10727
rect 9505 10693 9539 10727
rect 9873 10693 9907 10727
rect 17785 10693 17819 10727
rect 5365 10625 5399 10659
rect 7021 10625 7055 10659
rect 10701 10625 10735 10659
rect 14749 10625 14783 10659
rect 15945 10625 15979 10659
rect 17509 10625 17543 10659
rect 1869 10557 1903 10591
rect 2145 10557 2179 10591
rect 2421 10557 2455 10591
rect 3433 10557 3467 10591
rect 3709 10557 3743 10591
rect 7481 10557 7515 10591
rect 7757 10557 7791 10591
rect 10977 10557 11011 10591
rect 12081 10557 12115 10591
rect 12357 10557 12391 10591
rect 15025 10557 15059 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 16865 10557 16899 10591
rect 19717 10557 19751 10591
rect 19993 10557 20027 10591
rect 5181 10489 5215 10523
rect 10333 10489 10367 10523
rect 15577 10489 15611 10523
rect 21465 10489 21499 10523
rect 1685 10421 1719 10455
rect 6469 10421 6503 10455
rect 6837 10421 6871 10455
rect 11621 10421 11655 10455
rect 13829 10421 13863 10455
rect 14381 10421 14415 10455
rect 21833 10421 21867 10455
rect 22017 10421 22051 10455
rect 2697 10217 2731 10251
rect 3249 10217 3283 10251
rect 9137 10217 9171 10251
rect 10057 10217 10091 10251
rect 16589 10217 16623 10251
rect 16773 10217 16807 10251
rect 18889 10217 18923 10251
rect 21465 10217 21499 10251
rect 2973 10149 3007 10183
rect 3985 10149 4019 10183
rect 6377 10149 6411 10183
rect 6561 10149 6595 10183
rect 8585 10149 8619 10183
rect 14105 10149 14139 10183
rect 1593 10081 1627 10115
rect 4537 10081 4571 10115
rect 5825 10081 5859 10115
rect 6837 10081 6871 10115
rect 10701 10081 10735 10115
rect 13553 10081 13587 10115
rect 14841 10081 14875 10115
rect 19441 10081 19475 10115
rect 3157 10013 3191 10047
rect 3433 10013 3467 10047
rect 4261 10013 4295 10047
rect 10517 10013 10551 10047
rect 11253 10013 11287 10047
rect 14565 10013 14599 10047
rect 17141 10013 17175 10047
rect 7113 9945 7147 9979
rect 9413 9945 9447 9979
rect 11529 9945 11563 9979
rect 17417 9945 17451 9979
rect 19717 9945 19751 9979
rect 21649 9945 21683 9979
rect 1823 9877 1857 9911
rect 5365 9877 5399 9911
rect 10425 9877 10459 9911
rect 13001 9877 13035 9911
rect 16313 9877 16347 9911
rect 21189 9877 21223 9911
rect 6561 9673 6595 9707
rect 13829 9673 13863 9707
rect 13921 9673 13955 9707
rect 16221 9673 16255 9707
rect 1501 9605 1535 9639
rect 1685 9605 1719 9639
rect 3249 9605 3283 9639
rect 5641 9605 5675 9639
rect 5825 9605 5859 9639
rect 10793 9605 10827 9639
rect 11989 9605 12023 9639
rect 17141 9605 17175 9639
rect 19533 9605 19567 9639
rect 28641 9605 28675 9639
rect 1961 9537 1995 9571
rect 2237 9537 2271 9571
rect 3801 9537 3835 9571
rect 4261 9537 4295 9571
rect 7113 9537 7147 9571
rect 10701 9537 10735 9571
rect 19441 9537 19475 9571
rect 27537 9537 27571 9571
rect 4537 9469 4571 9503
rect 6837 9469 6871 9503
rect 8125 9469 8159 9503
rect 8401 9469 8435 9503
rect 10977 9469 11011 9503
rect 11713 9469 11747 9503
rect 14473 9469 14507 9503
rect 14749 9469 14783 9503
rect 16865 9469 16899 9503
rect 19717 9469 19751 9503
rect 27997 9469 28031 9503
rect 3617 9401 3651 9435
rect 13461 9401 13495 9435
rect 14105 9401 14139 9435
rect 19073 9401 19107 9435
rect 5549 9333 5583 9367
rect 9873 9333 9907 9367
rect 10333 9333 10367 9367
rect 18613 9333 18647 9367
rect 20085 9333 20119 9367
rect 27813 9333 27847 9367
rect 28457 9333 28491 9367
rect 3525 9129 3559 9163
rect 4629 9129 4663 9163
rect 5181 9129 5215 9163
rect 5457 9129 5491 9163
rect 7205 9129 7239 9163
rect 7849 9129 7883 9163
rect 10149 9129 10183 9163
rect 14289 9129 14323 9163
rect 17785 9129 17819 9163
rect 2881 9061 2915 9095
rect 15393 9061 15427 9095
rect 1593 8993 1627 9027
rect 1869 8993 1903 9027
rect 4721 8993 4755 9027
rect 6193 8993 6227 9027
rect 8493 8993 8527 9027
rect 9413 8993 9447 9027
rect 10793 8993 10827 9027
rect 11345 8993 11379 9027
rect 12633 8993 12667 9027
rect 14749 8993 14783 9027
rect 14933 8993 14967 9027
rect 16037 8993 16071 9027
rect 3065 8925 3099 8959
rect 3341 8925 3375 8959
rect 3893 8925 3927 8959
rect 3985 8925 4019 8959
rect 5917 8925 5951 8959
rect 7389 8925 7423 8959
rect 8217 8925 8251 8959
rect 11621 8925 11655 8959
rect 5549 8857 5583 8891
rect 10517 8857 10551 8891
rect 13553 8857 13587 8891
rect 14657 8857 14691 8891
rect 16313 8857 16347 8891
rect 8309 8789 8343 8823
rect 9045 8789 9079 8823
rect 10609 8789 10643 8823
rect 18153 8789 18187 8823
rect 18705 8789 18739 8823
rect 18981 8789 19015 8823
rect 3341 8585 3375 8619
rect 3617 8585 3651 8619
rect 3985 8585 4019 8619
rect 4629 8585 4663 8619
rect 5181 8585 5215 8619
rect 5825 8585 5859 8619
rect 6377 8585 6411 8619
rect 6653 8585 6687 8619
rect 8033 8585 8067 8619
rect 10149 8585 10183 8619
rect 10517 8585 10551 8619
rect 11161 8585 11195 8619
rect 11529 8585 11563 8619
rect 12173 8585 12207 8619
rect 12541 8585 12575 8619
rect 14289 8585 14323 8619
rect 15577 8585 15611 8619
rect 15945 8585 15979 8619
rect 7205 8517 7239 8551
rect 16037 8517 16071 8551
rect 1593 8449 1627 8483
rect 1869 8449 1903 8483
rect 3065 8449 3099 8483
rect 4169 8449 4203 8483
rect 4813 8449 4847 8483
rect 6009 8449 6043 8483
rect 7757 8449 7791 8483
rect 8677 8449 8711 8483
rect 12633 8449 12667 8483
rect 13645 8449 13679 8483
rect 14657 8449 14691 8483
rect 7389 8381 7423 8415
rect 8401 8381 8435 8415
rect 9689 8381 9723 8415
rect 10609 8381 10643 8415
rect 10793 8381 10827 8415
rect 12725 8381 12759 8415
rect 14749 8381 14783 8415
rect 14933 8381 14967 8415
rect 16221 8381 16255 8415
rect 6837 8313 6871 8347
rect 9873 8313 9907 8347
rect 2881 8245 2915 8279
rect 7849 8245 7883 8279
rect 1593 8041 1627 8075
rect 3341 8041 3375 8075
rect 3525 8041 3559 8075
rect 3893 8041 3927 8075
rect 4629 8041 4663 8075
rect 7573 8041 7607 8075
rect 9597 8041 9631 8075
rect 12449 8041 12483 8075
rect 13001 8041 13035 8075
rect 4261 7973 4295 8007
rect 7757 7973 7791 8007
rect 15209 7973 15243 8007
rect 3985 7905 4019 7939
rect 10057 7905 10091 7939
rect 10241 7905 10275 7939
rect 11529 7905 11563 7939
rect 13645 7905 13679 7939
rect 14105 7905 14139 7939
rect 1777 7837 1811 7871
rect 2421 7837 2455 7871
rect 3065 7837 3099 7871
rect 4445 7837 4479 7871
rect 11253 7837 11287 7871
rect 14841 7837 14875 7871
rect 15025 7837 15059 7871
rect 2237 7701 2271 7735
rect 2881 7701 2915 7735
rect 9965 7701 9999 7735
rect 13369 7701 13403 7735
rect 13461 7701 13495 7735
rect 15853 7701 15887 7735
rect 1593 7497 1627 7531
rect 2237 7497 2271 7531
rect 4353 7497 4387 7531
rect 9137 7497 9171 7531
rect 11897 7497 11931 7531
rect 13461 7497 13495 7531
rect 23949 7497 23983 7531
rect 1777 7361 1811 7395
rect 2421 7361 2455 7395
rect 3065 7361 3099 7395
rect 3709 7361 3743 7395
rect 9321 7361 9355 7395
rect 10793 7361 10827 7395
rect 12725 7361 12759 7395
rect 14289 7361 14323 7395
rect 22201 7361 22235 7395
rect 24225 7361 24259 7395
rect 4169 7293 4203 7327
rect 22477 7293 22511 7327
rect 3985 7225 4019 7259
rect 10609 7225 10643 7259
rect 2881 7157 2915 7191
rect 3525 7157 3559 7191
rect 12541 7157 12575 7191
rect 14105 7157 14139 7191
rect 3433 6953 3467 6987
rect 23213 6953 23247 6987
rect 3801 6817 3835 6851
rect 3985 6817 4019 6851
rect 10609 6817 10643 6851
rect 23765 6817 23799 6851
rect 1777 6749 1811 6783
rect 2421 6749 2455 6783
rect 3065 6749 3099 6783
rect 3525 6749 3559 6783
rect 4169 6749 4203 6783
rect 22937 6749 22971 6783
rect 1593 6613 1627 6647
rect 2237 6613 2271 6647
rect 2881 6613 2915 6647
rect 23397 6613 23431 6647
rect 2881 6409 2915 6443
rect 22845 6409 22879 6443
rect 3065 6273 3099 6307
rect 3341 6273 3375 6307
rect 22452 6273 22486 6307
rect 1593 6205 1627 6239
rect 1869 6205 1903 6239
rect 22523 6069 22557 6103
rect 2697 5865 2731 5899
rect 18889 5865 18923 5899
rect 21005 5865 21039 5899
rect 21741 5797 21775 5831
rect 1869 5729 1903 5763
rect 15577 5729 15611 5763
rect 17141 5729 17175 5763
rect 24869 5729 24903 5763
rect 26985 5729 27019 5763
rect 28825 5729 28859 5763
rect 1593 5661 1627 5695
rect 2881 5661 2915 5695
rect 15761 5661 15795 5695
rect 19349 5661 19383 5695
rect 20913 5661 20947 5695
rect 24685 5661 24719 5695
rect 17417 5593 17451 5627
rect 26525 5593 26559 5627
rect 27169 5593 27203 5627
rect 16221 5525 16255 5559
rect 21373 5525 21407 5559
rect 22891 5321 22925 5355
rect 1593 5185 1627 5219
rect 2697 5185 2731 5219
rect 15669 5185 15703 5219
rect 17509 5185 17543 5219
rect 22176 5185 22210 5219
rect 22788 5185 22822 5219
rect 1869 5117 1903 5151
rect 15853 5117 15887 5151
rect 17693 5117 17727 5151
rect 28641 5117 28675 5151
rect 28825 5117 28859 5151
rect 30021 5117 30055 5151
rect 2881 4981 2915 5015
rect 16313 4981 16347 5015
rect 18153 4981 18187 5015
rect 22247 4981 22281 5015
rect 2881 4777 2915 4811
rect 19533 4777 19567 4811
rect 20269 4777 20303 4811
rect 24731 4777 24765 4811
rect 1593 4641 1627 4675
rect 1869 4641 1903 4675
rect 25789 4641 25823 4675
rect 3065 4573 3099 4607
rect 3341 4573 3375 4607
rect 19441 4573 19475 4607
rect 24628 4573 24662 4607
rect 25973 4505 26007 4539
rect 27629 4505 27663 4539
rect 19901 4437 19935 4471
rect 1409 4233 1443 4267
rect 1869 4097 1903 4131
rect 2513 4097 2547 4131
rect 2973 4097 3007 4131
rect 4261 4097 4295 4131
rect 4537 4097 4571 4131
rect 15209 4097 15243 4131
rect 4077 3961 4111 3995
rect 3617 3893 3651 3927
rect 15025 3893 15059 3927
rect 3985 3689 4019 3723
rect 12081 3689 12115 3723
rect 2973 3621 3007 3655
rect 4629 3553 4663 3587
rect 1593 3485 1627 3519
rect 1869 3485 1903 3519
rect 3157 3485 3191 3519
rect 3433 3485 3467 3519
rect 4169 3485 4203 3519
rect 4445 3485 4479 3519
rect 11529 3485 11563 3519
rect 11621 3349 11655 3383
rect 14013 3145 14047 3179
rect 10793 3077 10827 3111
rect 12633 3077 12667 3111
rect 13921 3077 13955 3111
rect 15577 3077 15611 3111
rect 2881 3009 2915 3043
rect 3525 3009 3559 3043
rect 4169 3009 4203 3043
rect 6561 3009 6595 3043
rect 8769 3009 8803 3043
rect 17049 3009 17083 3043
rect 18337 3009 18371 3043
rect 20545 3009 20579 3043
rect 1593 2941 1627 2975
rect 1869 2941 1903 2975
rect 7205 2941 7239 2975
rect 9045 2941 9079 2975
rect 10517 2941 10551 2975
rect 3985 2873 4019 2907
rect 15761 2873 15795 2907
rect 12725 2805 12759 2839
rect 16865 2805 16899 2839
rect 18153 2805 18187 2839
rect 20361 2805 20395 2839
rect 2881 2601 2915 2635
rect 25513 2601 25547 2635
rect 28181 2601 28215 2635
rect 30849 2601 30883 2635
rect 33517 2601 33551 2635
rect 3525 2533 3559 2567
rect 1593 2465 1627 2499
rect 3801 2465 3835 2499
rect 4629 2465 4663 2499
rect 7297 2465 7331 2499
rect 9965 2465 9999 2499
rect 12633 2465 12667 2499
rect 15301 2465 15335 2499
rect 17969 2465 18003 2499
rect 20545 2465 20579 2499
rect 23121 2465 23155 2499
rect 36369 2465 36403 2499
rect 3065 2397 3099 2431
rect 4353 2397 4387 2431
rect 7021 2397 7055 2431
rect 9597 2397 9631 2431
rect 12357 2397 12391 2431
rect 15025 2397 15059 2431
rect 17509 2397 17543 2431
rect 20085 2397 20119 2431
rect 22661 2397 22695 2431
rect 25697 2397 25731 2431
rect 25973 2397 26007 2431
rect 28365 2397 28399 2431
rect 28641 2397 28675 2431
rect 31033 2397 31067 2431
rect 31309 2397 31343 2431
rect 33701 2397 33735 2431
rect 33977 2397 34011 2431
rect 36093 2397 36127 2431
rect 37289 2397 37323 2431
rect 3341 2329 3375 2363
rect 1823 2261 1857 2295
<< metal1 >>
rect 22830 25848 22836 25900
rect 22888 25888 22894 25900
rect 26786 25888 26792 25900
rect 22888 25860 26792 25888
rect 22888 25848 22894 25860
rect 26786 25848 26792 25860
rect 26844 25848 26850 25900
rect 25590 25780 25596 25832
rect 25648 25820 25654 25832
rect 29178 25820 29184 25832
rect 25648 25792 29184 25820
rect 25648 25780 25654 25792
rect 29178 25780 29184 25792
rect 29236 25780 29242 25832
rect 12158 25712 12164 25764
rect 12216 25752 12222 25764
rect 33686 25752 33692 25764
rect 12216 25724 33692 25752
rect 12216 25712 12222 25724
rect 33686 25712 33692 25724
rect 33744 25712 33750 25764
rect 10134 25644 10140 25696
rect 10192 25684 10198 25696
rect 26878 25684 26884 25696
rect 10192 25656 26884 25684
rect 10192 25644 10198 25656
rect 26878 25644 26884 25656
rect 26936 25644 26942 25696
rect 12802 25576 12808 25628
rect 12860 25616 12866 25628
rect 34790 25616 34796 25628
rect 12860 25588 34796 25616
rect 12860 25576 12866 25588
rect 34790 25576 34796 25588
rect 34848 25576 34854 25628
rect 10042 25508 10048 25560
rect 10100 25548 10106 25560
rect 33594 25548 33600 25560
rect 10100 25520 33600 25548
rect 10100 25508 10106 25520
rect 33594 25508 33600 25520
rect 33652 25508 33658 25560
rect 10778 25440 10784 25492
rect 10836 25480 10842 25492
rect 35618 25480 35624 25492
rect 10836 25452 35624 25480
rect 10836 25440 10842 25452
rect 35618 25440 35624 25452
rect 35676 25440 35682 25492
rect 15838 25372 15844 25424
rect 15896 25412 15902 25424
rect 32858 25412 32864 25424
rect 15896 25384 32864 25412
rect 15896 25372 15902 25384
rect 32858 25372 32864 25384
rect 32916 25372 32922 25424
rect 12250 25304 12256 25356
rect 12308 25344 12314 25356
rect 32214 25344 32220 25356
rect 12308 25316 32220 25344
rect 12308 25304 12314 25316
rect 32214 25304 32220 25316
rect 32272 25304 32278 25356
rect 13446 25236 13452 25288
rect 13504 25276 13510 25288
rect 32582 25276 32588 25288
rect 13504 25248 32588 25276
rect 13504 25236 13510 25248
rect 32582 25236 32588 25248
rect 32640 25236 32646 25288
rect 10226 25168 10232 25220
rect 10284 25208 10290 25220
rect 30282 25208 30288 25220
rect 10284 25180 30288 25208
rect 10284 25168 10290 25180
rect 30282 25168 30288 25180
rect 30340 25168 30346 25220
rect 15654 25100 15660 25152
rect 15712 25140 15718 25152
rect 27614 25140 27620 25152
rect 15712 25112 27620 25140
rect 15712 25100 15718 25112
rect 27614 25100 27620 25112
rect 27672 25100 27678 25152
rect 28258 25100 28264 25152
rect 28316 25140 28322 25152
rect 28718 25140 28724 25152
rect 28316 25112 28724 25140
rect 28316 25100 28322 25112
rect 28718 25100 28724 25112
rect 28776 25100 28782 25152
rect 3694 25032 3700 25084
rect 3752 25072 3758 25084
rect 7558 25072 7564 25084
rect 3752 25044 7564 25072
rect 3752 25032 3758 25044
rect 7558 25032 7564 25044
rect 7616 25032 7622 25084
rect 15470 25032 15476 25084
rect 15528 25072 15534 25084
rect 28442 25072 28448 25084
rect 15528 25044 28448 25072
rect 15528 25032 15534 25044
rect 28442 25032 28448 25044
rect 28500 25032 28506 25084
rect 15010 24964 15016 25016
rect 15068 25004 15074 25016
rect 25590 25004 25596 25016
rect 15068 24976 25596 25004
rect 15068 24964 15074 24976
rect 25590 24964 25596 24976
rect 25648 24964 25654 25016
rect 26142 24964 26148 25016
rect 26200 25004 26206 25016
rect 28994 25004 29000 25016
rect 26200 24976 29000 25004
rect 26200 24964 26206 24976
rect 28994 24964 29000 24976
rect 29052 24964 29058 25016
rect 14826 24896 14832 24948
rect 14884 24936 14890 24948
rect 39298 24936 39304 24948
rect 14884 24908 39304 24936
rect 14884 24896 14890 24908
rect 39298 24896 39304 24908
rect 39356 24896 39362 24948
rect 15194 24828 15200 24880
rect 15252 24868 15258 24880
rect 33502 24868 33508 24880
rect 15252 24840 33508 24868
rect 15252 24828 15258 24840
rect 33502 24828 33508 24840
rect 33560 24828 33566 24880
rect 25038 24760 25044 24812
rect 25096 24800 25102 24812
rect 30466 24800 30472 24812
rect 25096 24772 30472 24800
rect 25096 24760 25102 24772
rect 30466 24760 30472 24772
rect 30524 24760 30530 24812
rect 14274 24692 14280 24744
rect 14332 24732 14338 24744
rect 26234 24732 26240 24744
rect 14332 24704 26240 24732
rect 14332 24692 14338 24704
rect 26234 24692 26240 24704
rect 26292 24692 26298 24744
rect 27338 24692 27344 24744
rect 27396 24732 27402 24744
rect 29546 24732 29552 24744
rect 27396 24704 29552 24732
rect 27396 24692 27402 24704
rect 29546 24692 29552 24704
rect 29604 24692 29610 24744
rect 3050 24624 3056 24676
rect 3108 24664 3114 24676
rect 7282 24664 7288 24676
rect 3108 24636 7288 24664
rect 3108 24624 3114 24636
rect 7282 24624 7288 24636
rect 7340 24624 7346 24676
rect 14734 24624 14740 24676
rect 14792 24664 14798 24676
rect 30006 24664 30012 24676
rect 14792 24636 30012 24664
rect 14792 24624 14798 24636
rect 30006 24624 30012 24636
rect 30064 24624 30070 24676
rect 32490 24624 32496 24676
rect 32548 24664 32554 24676
rect 36262 24664 36268 24676
rect 32548 24636 36268 24664
rect 32548 24624 32554 24636
rect 36262 24624 36268 24636
rect 36320 24624 36326 24676
rect 3418 24556 3424 24608
rect 3476 24596 3482 24608
rect 12250 24596 12256 24608
rect 3476 24568 12256 24596
rect 3476 24556 3482 24568
rect 12250 24556 12256 24568
rect 12308 24556 12314 24608
rect 15930 24556 15936 24608
rect 15988 24596 15994 24608
rect 25682 24596 25688 24608
rect 15988 24568 25688 24596
rect 15988 24556 15994 24568
rect 25682 24556 25688 24568
rect 25740 24556 25746 24608
rect 27614 24556 27620 24608
rect 27672 24596 27678 24608
rect 34146 24596 34152 24608
rect 27672 24568 34152 24596
rect 27672 24556 27678 24568
rect 34146 24556 34152 24568
rect 34204 24556 34210 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 3973 24395 4031 24401
rect 3973 24361 3985 24395
rect 4019 24392 4031 24395
rect 6549 24395 6607 24401
rect 4019 24364 6500 24392
rect 4019 24361 4031 24364
rect 3973 24355 4031 24361
rect 1486 24284 1492 24336
rect 1544 24324 1550 24336
rect 6472 24324 6500 24364
rect 6549 24361 6561 24395
rect 6595 24392 6607 24395
rect 9674 24392 9680 24404
rect 6595 24364 9680 24392
rect 6595 24361 6607 24364
rect 6549 24355 6607 24361
rect 9674 24352 9680 24364
rect 9732 24352 9738 24404
rect 11701 24395 11759 24401
rect 11701 24361 11713 24395
rect 11747 24392 11759 24395
rect 23845 24395 23903 24401
rect 11747 24364 20208 24392
rect 11747 24361 11759 24364
rect 11701 24355 11759 24361
rect 14458 24324 14464 24336
rect 1544 24296 4660 24324
rect 6472 24296 13308 24324
rect 1544 24284 1550 24296
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3510 24256 3516 24268
rect 3283 24228 3516 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2406 24188 2412 24200
rect 2271 24160 2412 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2406 24148 2412 24160
rect 2464 24148 2470 24200
rect 3881 24191 3939 24197
rect 3881 24157 3893 24191
rect 3927 24188 3939 24191
rect 4157 24191 4215 24197
rect 4157 24188 4169 24191
rect 3927 24160 4169 24188
rect 3927 24157 3939 24160
rect 3881 24151 3939 24157
rect 4157 24157 4169 24160
rect 4203 24188 4215 24191
rect 4246 24188 4252 24200
rect 4203 24160 4252 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4246 24148 4252 24160
rect 4304 24148 4310 24200
rect 4632 24197 4660 24296
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 6822 24256 6828 24268
rect 5859 24228 6828 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 6822 24216 6828 24228
rect 6880 24216 6886 24268
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9214 24256 9220 24268
rect 8251 24228 9220 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 9214 24216 9220 24228
rect 9272 24216 9278 24268
rect 13170 24256 13176 24268
rect 9692 24228 13176 24256
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 6457 24191 6515 24197
rect 6457 24157 6469 24191
rect 6503 24188 6515 24191
rect 6638 24188 6644 24200
rect 6503 24160 6644 24188
rect 6503 24157 6515 24160
rect 6457 24151 6515 24157
rect 6638 24148 6644 24160
rect 6696 24188 6702 24200
rect 6733 24191 6791 24197
rect 6733 24188 6745 24191
rect 6696 24160 6745 24188
rect 6696 24148 6702 24160
rect 6733 24157 6745 24160
rect 6779 24157 6791 24191
rect 6733 24151 6791 24157
rect 7377 24191 7435 24197
rect 7377 24157 7389 24191
rect 7423 24188 7435 24191
rect 8570 24188 8576 24200
rect 7423 24160 8576 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 8570 24148 8576 24160
rect 8628 24148 8634 24200
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24188 9367 24191
rect 9692 24188 9720 24228
rect 13170 24216 13176 24228
rect 13228 24216 13234 24268
rect 9355 24160 9720 24188
rect 9953 24191 10011 24197
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 9953 24157 9965 24191
rect 9999 24188 10011 24191
rect 10134 24188 10140 24200
rect 9999 24160 10140 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 12434 24188 12440 24200
rect 11931 24160 12440 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 12434 24148 12440 24160
rect 12492 24148 12498 24200
rect 12529 24191 12587 24197
rect 12529 24157 12541 24191
rect 12575 24188 12587 24191
rect 12618 24188 12624 24200
rect 12575 24160 12624 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 12618 24148 12624 24160
rect 12676 24188 12682 24200
rect 12802 24188 12808 24200
rect 12676 24160 12808 24188
rect 12676 24148 12682 24160
rect 12802 24148 12808 24160
rect 12860 24148 12866 24200
rect 13280 24188 13308 24296
rect 13556 24296 14464 24324
rect 13556 24265 13584 24296
rect 14458 24284 14464 24296
rect 14516 24284 14522 24336
rect 13541 24259 13599 24265
rect 13541 24225 13553 24259
rect 13587 24225 13599 24259
rect 13541 24219 13599 24225
rect 16117 24259 16175 24265
rect 16117 24225 16129 24259
rect 16163 24256 16175 24259
rect 16206 24256 16212 24268
rect 16163 24228 16212 24256
rect 16163 24225 16175 24228
rect 16117 24219 16175 24225
rect 16206 24216 16212 24228
rect 16264 24216 16270 24268
rect 16853 24259 16911 24265
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 18690 24256 18696 24268
rect 16899 24228 18696 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 18690 24216 18696 24228
rect 18748 24216 18754 24268
rect 14182 24188 14188 24200
rect 13280 24160 14188 24188
rect 14182 24148 14188 24160
rect 14240 24148 14246 24200
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24188 15163 24191
rect 18969 24191 19027 24197
rect 18969 24188 18981 24191
rect 15151 24160 15516 24188
rect 18262 24160 18981 24188
rect 15151 24157 15163 24160
rect 15105 24151 15163 24157
rect 2774 24080 2780 24132
rect 2832 24120 2838 24132
rect 4430 24120 4436 24132
rect 2832 24092 4436 24120
rect 2832 24080 2838 24092
rect 4430 24080 4436 24092
rect 4488 24080 4494 24132
rect 10965 24123 11023 24129
rect 10965 24089 10977 24123
rect 11011 24120 11023 24123
rect 13814 24120 13820 24132
rect 11011 24092 13820 24120
rect 11011 24089 11023 24092
rect 10965 24083 11023 24089
rect 13814 24080 13820 24092
rect 13872 24080 13878 24132
rect 15378 24120 15384 24132
rect 13924 24092 15384 24120
rect 1581 24055 1639 24061
rect 1581 24021 1593 24055
rect 1627 24052 1639 24055
rect 1673 24055 1731 24061
rect 1673 24052 1685 24055
rect 1627 24024 1685 24052
rect 1627 24021 1639 24024
rect 1581 24015 1639 24021
rect 1673 24021 1685 24024
rect 1719 24052 1731 24055
rect 3510 24052 3516 24064
rect 1719 24024 3516 24052
rect 1719 24021 1731 24024
rect 1673 24015 1731 24021
rect 3510 24012 3516 24024
rect 3568 24012 3574 24064
rect 3694 24012 3700 24064
rect 3752 24052 3758 24064
rect 8754 24052 8760 24064
rect 3752 24024 8760 24052
rect 3752 24012 3758 24024
rect 8754 24012 8760 24024
rect 8812 24012 8818 24064
rect 9125 24055 9183 24061
rect 9125 24021 9137 24055
rect 9171 24052 9183 24055
rect 12066 24052 12072 24064
rect 9171 24024 12072 24052
rect 9171 24021 9183 24024
rect 9125 24015 9183 24021
rect 12066 24012 12072 24024
rect 12124 24012 12130 24064
rect 12434 24012 12440 24064
rect 12492 24052 12498 24064
rect 13924 24052 13952 24092
rect 15378 24080 15384 24092
rect 15436 24080 15442 24132
rect 12492 24024 13952 24052
rect 12492 24012 12498 24024
rect 14274 24012 14280 24064
rect 14332 24012 14338 24064
rect 15488 24052 15516 24160
rect 18969 24157 18981 24160
rect 19015 24188 19027 24191
rect 19058 24188 19064 24200
rect 19015 24160 19064 24188
rect 19015 24157 19027 24160
rect 18969 24151 19027 24157
rect 19058 24148 19064 24160
rect 19116 24148 19122 24200
rect 19150 24148 19156 24200
rect 19208 24188 19214 24200
rect 19613 24191 19671 24197
rect 19613 24188 19625 24191
rect 19208 24160 19625 24188
rect 19208 24148 19214 24160
rect 19613 24157 19625 24160
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 19794 24148 19800 24200
rect 19852 24188 19858 24200
rect 20073 24191 20131 24197
rect 20073 24188 20085 24191
rect 19852 24160 20085 24188
rect 19852 24148 19858 24160
rect 20073 24157 20085 24160
rect 20119 24157 20131 24191
rect 20180 24188 20208 24364
rect 23845 24361 23857 24395
rect 23891 24392 23903 24395
rect 23891 24364 25636 24392
rect 23891 24361 23903 24364
rect 23845 24355 23903 24361
rect 25608 24324 25636 24364
rect 25682 24352 25688 24404
rect 25740 24392 25746 24404
rect 25777 24395 25835 24401
rect 25777 24392 25789 24395
rect 25740 24364 25789 24392
rect 25740 24352 25746 24364
rect 25777 24361 25789 24364
rect 25823 24361 25835 24395
rect 25777 24355 25835 24361
rect 25866 24352 25872 24404
rect 25924 24392 25930 24404
rect 29086 24392 29092 24404
rect 25924 24364 29092 24392
rect 25924 24352 25930 24364
rect 29086 24352 29092 24364
rect 29144 24352 29150 24404
rect 31297 24395 31355 24401
rect 31297 24392 31309 24395
rect 29196 24364 31309 24392
rect 25608 24296 26464 24324
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 21542 24216 21548 24268
rect 21600 24256 21606 24268
rect 22465 24259 22523 24265
rect 22465 24256 22477 24259
rect 21600 24228 22477 24256
rect 21600 24216 21606 24228
rect 22465 24225 22477 24228
rect 22511 24225 22523 24259
rect 22465 24219 22523 24225
rect 25038 24216 25044 24268
rect 25096 24216 25102 24268
rect 25225 24259 25283 24265
rect 25225 24225 25237 24259
rect 25271 24225 25283 24259
rect 25225 24219 25283 24225
rect 22005 24191 22063 24197
rect 22005 24188 22017 24191
rect 20180 24160 22017 24188
rect 20073 24151 20131 24157
rect 22005 24157 22017 24160
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 24026 24148 24032 24200
rect 24084 24188 24090 24200
rect 24946 24188 24952 24200
rect 24084 24160 24952 24188
rect 24084 24148 24090 24160
rect 24946 24148 24952 24160
rect 25004 24148 25010 24200
rect 25240 24188 25268 24219
rect 25314 24216 25320 24268
rect 25372 24256 25378 24268
rect 26329 24259 26387 24265
rect 26329 24256 26341 24259
rect 25372 24228 26341 24256
rect 25372 24216 25378 24228
rect 26329 24225 26341 24228
rect 26375 24225 26387 24259
rect 26436 24256 26464 24296
rect 26510 24284 26516 24336
rect 26568 24324 26574 24336
rect 27157 24327 27215 24333
rect 27157 24324 27169 24327
rect 26568 24296 27169 24324
rect 26568 24284 26574 24296
rect 27157 24293 27169 24296
rect 27203 24293 27215 24327
rect 27157 24287 27215 24293
rect 27890 24284 27896 24336
rect 27948 24324 27954 24336
rect 28997 24327 29055 24333
rect 28997 24324 29009 24327
rect 27948 24296 29009 24324
rect 27948 24284 27954 24296
rect 28997 24293 29009 24296
rect 29043 24293 29055 24327
rect 28997 24287 29055 24293
rect 27617 24259 27675 24265
rect 27617 24256 27629 24259
rect 26436 24228 27629 24256
rect 26329 24219 26387 24225
rect 27617 24225 27629 24228
rect 27663 24225 27675 24259
rect 27617 24219 27675 24225
rect 27709 24259 27767 24265
rect 27709 24225 27721 24259
rect 27755 24225 27767 24259
rect 27709 24219 27767 24225
rect 25866 24188 25872 24200
rect 25240 24160 25872 24188
rect 25866 24148 25872 24160
rect 25924 24148 25930 24200
rect 25958 24148 25964 24200
rect 26016 24188 26022 24200
rect 26145 24191 26203 24197
rect 26145 24188 26157 24191
rect 26016 24160 26157 24188
rect 26016 24148 26022 24160
rect 26145 24157 26157 24160
rect 26191 24157 26203 24191
rect 26145 24151 26203 24157
rect 26234 24148 26240 24200
rect 26292 24148 26298 24200
rect 26418 24148 26424 24200
rect 26476 24188 26482 24200
rect 27724 24188 27752 24219
rect 27798 24216 27804 24268
rect 27856 24256 27862 24268
rect 29196 24256 29224 24364
rect 31297 24361 31309 24364
rect 31343 24361 31355 24395
rect 31297 24355 31355 24361
rect 34146 24352 34152 24404
rect 34204 24352 34210 24404
rect 35728 24364 39252 24392
rect 29748 24296 30328 24324
rect 27856 24228 29224 24256
rect 27856 24216 27862 24228
rect 29270 24216 29276 24268
rect 29328 24256 29334 24268
rect 29748 24265 29776 24296
rect 29733 24259 29791 24265
rect 29733 24256 29745 24259
rect 29328 24228 29745 24256
rect 29328 24216 29334 24228
rect 29733 24225 29745 24228
rect 29779 24225 29791 24259
rect 29733 24219 29791 24225
rect 30006 24216 30012 24268
rect 30064 24216 30070 24268
rect 30300 24256 30328 24296
rect 30374 24284 30380 24336
rect 30432 24324 30438 24336
rect 35728 24324 35756 24364
rect 30432 24296 35756 24324
rect 30432 24284 30438 24296
rect 35802 24284 35808 24336
rect 35860 24324 35866 24336
rect 36357 24327 36415 24333
rect 36357 24324 36369 24327
rect 35860 24296 36369 24324
rect 35860 24284 35866 24296
rect 36357 24293 36369 24296
rect 36403 24293 36415 24327
rect 36357 24287 36415 24293
rect 36906 24284 36912 24336
rect 36964 24324 36970 24336
rect 37461 24327 37519 24333
rect 37461 24324 37473 24327
rect 36964 24296 37473 24324
rect 36964 24284 36970 24296
rect 37461 24293 37473 24296
rect 37507 24293 37519 24327
rect 37461 24287 37519 24293
rect 38654 24284 38660 24336
rect 38712 24284 38718 24336
rect 39224 24324 39252 24364
rect 39298 24352 39304 24404
rect 39356 24352 39362 24404
rect 44726 24352 44732 24404
rect 44784 24352 44790 24404
rect 40678 24324 40684 24336
rect 39224 24296 40684 24324
rect 40678 24284 40684 24296
rect 40736 24284 40742 24336
rect 37001 24259 37059 24265
rect 37001 24256 37013 24259
rect 30300 24228 37013 24256
rect 37001 24225 37013 24228
rect 37047 24225 37059 24259
rect 37001 24219 37059 24225
rect 39574 24216 39580 24268
rect 39632 24256 39638 24268
rect 40037 24259 40095 24265
rect 40037 24256 40049 24259
rect 39632 24228 40049 24256
rect 39632 24216 39638 24228
rect 40037 24225 40049 24228
rect 40083 24225 40095 24259
rect 40037 24219 40095 24225
rect 40126 24216 40132 24268
rect 40184 24256 40190 24268
rect 40313 24259 40371 24265
rect 40313 24256 40325 24259
rect 40184 24228 40325 24256
rect 40184 24216 40190 24228
rect 40313 24225 40325 24228
rect 40359 24225 40371 24259
rect 40313 24219 40371 24225
rect 28537 24191 28595 24197
rect 28537 24188 28549 24191
rect 26476 24160 27752 24188
rect 28184 24184 28304 24188
rect 28460 24184 28549 24188
rect 28184 24160 28549 24184
rect 26476 24148 26482 24160
rect 17129 24123 17187 24129
rect 17129 24089 17141 24123
rect 17175 24120 17187 24123
rect 17218 24120 17224 24132
rect 17175 24092 17224 24120
rect 17175 24089 17187 24092
rect 17129 24083 17187 24089
rect 17218 24080 17224 24092
rect 17276 24080 17282 24132
rect 18782 24080 18788 24132
rect 18840 24120 18846 24132
rect 25314 24120 25320 24132
rect 18840 24092 25320 24120
rect 18840 24080 18846 24092
rect 25314 24080 25320 24092
rect 25372 24080 25378 24132
rect 25498 24080 25504 24132
rect 25556 24120 25562 24132
rect 27430 24120 27436 24132
rect 25556 24092 27436 24120
rect 25556 24080 25562 24092
rect 27430 24080 27436 24092
rect 27488 24080 27494 24132
rect 27522 24080 27528 24132
rect 27580 24080 27586 24132
rect 27614 24080 27620 24132
rect 27672 24120 27678 24132
rect 28184 24120 28212 24160
rect 28276 24156 28488 24160
rect 28537 24157 28549 24160
rect 28583 24157 28595 24191
rect 28537 24151 28595 24157
rect 28552 24120 28580 24151
rect 28994 24148 29000 24200
rect 29052 24188 29058 24200
rect 29181 24191 29239 24197
rect 29181 24188 29193 24191
rect 29052 24160 29193 24188
rect 29052 24148 29058 24160
rect 29181 24157 29193 24160
rect 29227 24188 29239 24191
rect 30190 24188 30196 24200
rect 29227 24160 30196 24188
rect 29227 24157 29239 24160
rect 29181 24151 29239 24157
rect 30190 24148 30196 24160
rect 30248 24148 30254 24200
rect 30558 24148 30564 24200
rect 30616 24188 30622 24200
rect 31481 24191 31539 24197
rect 31481 24188 31493 24191
rect 30616 24160 31493 24188
rect 30616 24148 30622 24160
rect 31481 24157 31493 24160
rect 31527 24188 31539 24191
rect 31570 24188 31576 24200
rect 31527 24160 31576 24188
rect 31527 24157 31539 24160
rect 31481 24151 31539 24157
rect 31570 24148 31576 24160
rect 31628 24148 31634 24200
rect 31846 24148 31852 24200
rect 31904 24188 31910 24200
rect 32493 24191 32551 24197
rect 32493 24188 32505 24191
rect 31904 24160 32505 24188
rect 31904 24148 31910 24160
rect 32493 24157 32505 24160
rect 32539 24188 32551 24191
rect 32674 24188 32680 24200
rect 32539 24160 32680 24188
rect 32539 24157 32551 24160
rect 32493 24151 32551 24157
rect 32674 24148 32680 24160
rect 32732 24148 32738 24200
rect 33318 24148 33324 24200
rect 33376 24148 33382 24200
rect 34054 24148 34060 24200
rect 34112 24188 34118 24200
rect 34112 24160 35848 24188
rect 34112 24148 34118 24160
rect 32769 24123 32827 24129
rect 32769 24120 32781 24123
rect 27672 24092 28212 24120
rect 28276 24092 28488 24120
rect 28552 24092 32781 24120
rect 27672 24080 27678 24092
rect 16942 24052 16948 24064
rect 15488 24024 16948 24052
rect 16942 24012 16948 24024
rect 17000 24012 17006 24064
rect 17034 24012 17040 24064
rect 17092 24052 17098 24064
rect 18601 24055 18659 24061
rect 18601 24052 18613 24055
rect 17092 24024 18613 24052
rect 17092 24012 17098 24024
rect 18601 24021 18613 24024
rect 18647 24021 18659 24055
rect 18601 24015 18659 24021
rect 19429 24055 19487 24061
rect 19429 24021 19441 24055
rect 19475 24052 19487 24055
rect 20346 24052 20352 24064
rect 19475 24024 20352 24052
rect 19475 24021 19487 24024
rect 19429 24015 19487 24021
rect 20346 24012 20352 24024
rect 20404 24012 20410 24064
rect 24302 24012 24308 24064
rect 24360 24052 24366 24064
rect 24581 24055 24639 24061
rect 24581 24052 24593 24055
rect 24360 24024 24593 24052
rect 24360 24012 24366 24024
rect 24581 24021 24593 24024
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 24946 24012 24952 24064
rect 25004 24012 25010 24064
rect 25130 24012 25136 24064
rect 25188 24052 25194 24064
rect 28276 24052 28304 24092
rect 25188 24024 28304 24052
rect 25188 24012 25194 24024
rect 28350 24012 28356 24064
rect 28408 24012 28414 24064
rect 28460 24052 28488 24092
rect 32769 24089 32781 24092
rect 32815 24089 32827 24123
rect 32769 24083 32827 24089
rect 34514 24080 34520 24132
rect 34572 24120 34578 24132
rect 34974 24120 34980 24132
rect 34572 24092 34980 24120
rect 34572 24080 34578 24092
rect 34974 24080 34980 24092
rect 35032 24080 35038 24132
rect 35158 24080 35164 24132
rect 35216 24120 35222 24132
rect 35710 24120 35716 24132
rect 35216 24092 35716 24120
rect 35216 24080 35222 24092
rect 35710 24080 35716 24092
rect 35768 24080 35774 24132
rect 35820 24120 35848 24160
rect 35894 24148 35900 24200
rect 35952 24188 35958 24200
rect 36541 24191 36599 24197
rect 36541 24188 36553 24191
rect 35952 24160 36553 24188
rect 35952 24148 35958 24160
rect 36541 24157 36553 24160
rect 36587 24188 36599 24191
rect 36814 24188 36820 24200
rect 36587 24160 36820 24188
rect 36587 24157 36599 24160
rect 36541 24151 36599 24157
rect 36814 24148 36820 24160
rect 36872 24148 36878 24200
rect 37274 24148 37280 24200
rect 37332 24188 37338 24200
rect 37645 24191 37703 24197
rect 37645 24188 37657 24191
rect 37332 24160 37657 24188
rect 37332 24148 37338 24160
rect 37645 24157 37657 24160
rect 37691 24157 37703 24191
rect 37645 24151 37703 24157
rect 38470 24148 38476 24200
rect 38528 24148 38534 24200
rect 39206 24148 39212 24200
rect 39264 24148 39270 24200
rect 41417 24191 41475 24197
rect 41417 24157 41429 24191
rect 41463 24188 41475 24191
rect 41506 24188 41512 24200
rect 41463 24160 41512 24188
rect 41463 24157 41475 24160
rect 41417 24151 41475 24157
rect 41506 24148 41512 24160
rect 41564 24188 41570 24200
rect 42429 24191 42487 24197
rect 42429 24188 42441 24191
rect 41564 24160 42441 24188
rect 41564 24148 41570 24160
rect 42429 24157 42441 24160
rect 42475 24157 42487 24191
rect 42429 24151 42487 24157
rect 44358 24148 44364 24200
rect 44416 24148 44422 24200
rect 44726 24148 44732 24200
rect 44784 24188 44790 24200
rect 45189 24191 45247 24197
rect 45189 24188 45201 24191
rect 44784 24160 45201 24188
rect 44784 24148 44790 24160
rect 45189 24157 45201 24160
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 45554 24148 45560 24200
rect 45612 24188 45618 24200
rect 45922 24188 45928 24200
rect 45612 24160 45928 24188
rect 45612 24148 45618 24160
rect 45922 24148 45928 24160
rect 45980 24148 45986 24200
rect 46014 24148 46020 24200
rect 46072 24188 46078 24200
rect 46661 24191 46719 24197
rect 46661 24188 46673 24191
rect 46072 24160 46673 24188
rect 46072 24148 46078 24160
rect 46661 24157 46673 24160
rect 46707 24188 46719 24191
rect 47213 24191 47271 24197
rect 47213 24188 47225 24191
rect 46707 24160 47225 24188
rect 46707 24157 46719 24160
rect 46661 24151 46719 24157
rect 47213 24157 47225 24160
rect 47259 24157 47271 24191
rect 47213 24151 47271 24157
rect 47302 24148 47308 24200
rect 47360 24188 47366 24200
rect 47765 24191 47823 24197
rect 47765 24188 47777 24191
rect 47360 24160 47777 24188
rect 47360 24148 47366 24160
rect 47765 24157 47777 24160
rect 47811 24157 47823 24191
rect 47765 24151 47823 24157
rect 48590 24148 48596 24200
rect 48648 24148 48654 24200
rect 37921 24123 37979 24129
rect 37921 24120 37933 24123
rect 35820 24092 37933 24120
rect 37921 24089 37933 24092
rect 37967 24089 37979 24123
rect 37921 24083 37979 24089
rect 38286 24080 38292 24132
rect 38344 24120 38350 24132
rect 38344 24092 45554 24120
rect 38344 24080 38350 24092
rect 30374 24052 30380 24064
rect 28460 24024 30380 24052
rect 30374 24012 30380 24024
rect 30432 24012 30438 24064
rect 30929 24055 30987 24061
rect 30929 24021 30941 24055
rect 30975 24052 30987 24055
rect 31846 24052 31852 24064
rect 30975 24024 31852 24052
rect 30975 24021 30987 24024
rect 30929 24015 30987 24021
rect 31846 24012 31852 24024
rect 31904 24012 31910 24064
rect 32306 24012 32312 24064
rect 32364 24012 32370 24064
rect 33410 24012 33416 24064
rect 33468 24012 33474 24064
rect 35066 24012 35072 24064
rect 35124 24012 35130 24064
rect 35805 24055 35863 24061
rect 35805 24021 35817 24055
rect 35851 24052 35863 24055
rect 35986 24052 35992 24064
rect 35851 24024 35992 24052
rect 35851 24021 35863 24024
rect 35805 24015 35863 24021
rect 35986 24012 35992 24024
rect 36044 24012 36050 24064
rect 36446 24012 36452 24064
rect 36504 24052 36510 24064
rect 36817 24055 36875 24061
rect 36817 24052 36829 24055
rect 36504 24024 36829 24052
rect 36504 24012 36510 24024
rect 36817 24021 36829 24024
rect 36863 24021 36875 24055
rect 36817 24015 36875 24021
rect 42058 24012 42064 24064
rect 42116 24012 42122 24064
rect 43714 24012 43720 24064
rect 43772 24052 43778 24064
rect 44177 24055 44235 24061
rect 44177 24052 44189 24055
rect 43772 24024 44189 24052
rect 43772 24012 43778 24024
rect 44177 24021 44189 24024
rect 44223 24021 44235 24055
rect 44177 24015 44235 24021
rect 45370 24012 45376 24064
rect 45428 24012 45434 24064
rect 45526 24052 45554 24092
rect 46109 24055 46167 24061
rect 46109 24052 46121 24055
rect 45526 24024 46121 24052
rect 46109 24021 46121 24024
rect 46155 24021 46167 24055
rect 46109 24015 46167 24021
rect 46842 24012 46848 24064
rect 46900 24012 46906 24064
rect 47118 24012 47124 24064
rect 47176 24052 47182 24064
rect 47949 24055 48007 24061
rect 47949 24052 47961 24055
rect 47176 24024 47961 24052
rect 47176 24012 47182 24024
rect 47949 24021 47961 24024
rect 47995 24021 48007 24055
rect 47949 24015 48007 24021
rect 48682 24012 48688 24064
rect 48740 24052 48746 24064
rect 49237 24055 49295 24061
rect 49237 24052 49249 24055
rect 48740 24024 49249 24052
rect 48740 24012 48746 24024
rect 49237 24021 49249 24024
rect 49283 24021 49295 24055
rect 49237 24015 49295 24021
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 1765 23851 1823 23857
rect 1765 23817 1777 23851
rect 1811 23848 1823 23851
rect 3694 23848 3700 23860
rect 1811 23820 3700 23848
rect 1811 23817 1823 23820
rect 1765 23811 1823 23817
rect 3694 23808 3700 23820
rect 3752 23808 3758 23860
rect 5718 23848 5724 23860
rect 3896 23820 5724 23848
rect 1581 23783 1639 23789
rect 1581 23749 1593 23783
rect 1627 23780 1639 23783
rect 3896 23780 3924 23820
rect 5718 23808 5724 23820
rect 5776 23808 5782 23860
rect 7098 23808 7104 23860
rect 7156 23848 7162 23860
rect 11885 23851 11943 23857
rect 11885 23848 11897 23851
rect 7156 23820 11897 23848
rect 7156 23808 7162 23820
rect 11885 23817 11897 23820
rect 11931 23817 11943 23851
rect 11885 23811 11943 23817
rect 12250 23808 12256 23860
rect 12308 23808 12314 23860
rect 12345 23851 12403 23857
rect 12345 23817 12357 23851
rect 12391 23848 12403 23851
rect 15930 23848 15936 23860
rect 12391 23820 15936 23848
rect 12391 23817 12403 23820
rect 12345 23811 12403 23817
rect 15930 23808 15936 23820
rect 15988 23808 15994 23860
rect 17126 23848 17132 23860
rect 16040 23820 17132 23848
rect 1627 23752 3924 23780
rect 3973 23783 4031 23789
rect 1627 23749 1639 23752
rect 1581 23743 1639 23749
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 4154 23780 4160 23792
rect 4019 23752 4160 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 4154 23740 4160 23752
rect 4212 23740 4218 23792
rect 8478 23780 8484 23792
rect 4264 23752 8484 23780
rect 2130 23672 2136 23724
rect 2188 23672 2194 23724
rect 2682 23672 2688 23724
rect 2740 23712 2746 23724
rect 2777 23715 2835 23721
rect 2777 23712 2789 23715
rect 2740 23684 2789 23712
rect 2740 23672 2746 23684
rect 2777 23681 2789 23684
rect 2823 23681 2835 23715
rect 2777 23675 2835 23681
rect 3878 23672 3884 23724
rect 3936 23712 3942 23724
rect 4264 23712 4292 23752
rect 8478 23740 8484 23752
rect 8536 23740 8542 23792
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9950 23780 9956 23792
rect 9171 23752 9956 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 9950 23740 9956 23752
rect 10008 23740 10014 23792
rect 10965 23783 11023 23789
rect 10965 23749 10977 23783
rect 11011 23780 11023 23783
rect 12526 23780 12532 23792
rect 11011 23752 12532 23780
rect 11011 23749 11023 23752
rect 10965 23743 11023 23749
rect 12526 23740 12532 23752
rect 12584 23740 12590 23792
rect 14277 23783 14335 23789
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 15746 23780 15752 23792
rect 14323 23752 15752 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 15746 23740 15752 23752
rect 15804 23740 15810 23792
rect 3936 23684 4292 23712
rect 3936 23672 3942 23684
rect 4798 23672 4804 23724
rect 4856 23672 4862 23724
rect 6546 23672 6552 23724
rect 6604 23712 6610 23724
rect 7101 23715 7159 23721
rect 7101 23712 7113 23715
rect 6604 23684 7113 23712
rect 6604 23672 6610 23684
rect 7101 23681 7113 23684
rect 7147 23681 7159 23715
rect 7101 23675 7159 23681
rect 7193 23715 7251 23721
rect 7193 23681 7205 23715
rect 7239 23712 7251 23715
rect 7742 23712 7748 23724
rect 7239 23684 7748 23712
rect 7239 23681 7251 23684
rect 7193 23675 7251 23681
rect 7742 23672 7748 23684
rect 7800 23672 7806 23724
rect 7926 23672 7932 23724
rect 7984 23672 7990 23724
rect 9861 23715 9919 23721
rect 9861 23681 9873 23715
rect 9907 23712 9919 23715
rect 11422 23712 11428 23724
rect 9907 23684 11428 23712
rect 9907 23681 9919 23684
rect 9861 23675 9919 23681
rect 11422 23672 11428 23684
rect 11480 23672 11486 23724
rect 11514 23672 11520 23724
rect 11572 23712 11578 23724
rect 12250 23712 12256 23724
rect 11572 23684 12256 23712
rect 11572 23672 11578 23684
rect 12250 23672 12256 23684
rect 12308 23712 12314 23724
rect 12802 23712 12808 23724
rect 12308 23684 12808 23712
rect 12308 23672 12314 23684
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23712 13323 23715
rect 13538 23712 13544 23724
rect 13311 23684 13544 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 13538 23672 13544 23684
rect 13596 23672 13602 23724
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23712 15163 23715
rect 16040 23712 16068 23820
rect 17126 23808 17132 23820
rect 17184 23808 17190 23860
rect 17218 23808 17224 23860
rect 17276 23848 17282 23860
rect 18782 23848 18788 23860
rect 17276 23820 18788 23848
rect 17276 23808 17282 23820
rect 18782 23808 18788 23820
rect 18840 23808 18846 23860
rect 24213 23851 24271 23857
rect 18984 23820 24164 23848
rect 16117 23783 16175 23789
rect 16117 23749 16129 23783
rect 16163 23780 16175 23783
rect 18322 23780 18328 23792
rect 16163 23752 18328 23780
rect 16163 23749 16175 23752
rect 16117 23743 16175 23749
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 18874 23740 18880 23792
rect 18932 23780 18938 23792
rect 18984 23789 19012 23820
rect 18969 23783 19027 23789
rect 18969 23780 18981 23783
rect 18932 23752 18981 23780
rect 18932 23740 18938 23752
rect 18969 23749 18981 23752
rect 19015 23749 19027 23783
rect 18969 23743 19027 23749
rect 19058 23740 19064 23792
rect 19116 23780 19122 23792
rect 19116 23752 19458 23780
rect 19116 23740 19122 23752
rect 21174 23740 21180 23792
rect 21232 23740 21238 23792
rect 21818 23740 21824 23792
rect 21876 23780 21882 23792
rect 22281 23783 22339 23789
rect 22281 23780 22293 23783
rect 21876 23752 22293 23780
rect 21876 23740 21882 23752
rect 22281 23749 22293 23752
rect 22327 23749 22339 23783
rect 22281 23743 22339 23749
rect 23290 23740 23296 23792
rect 23348 23740 23354 23792
rect 24136 23780 24164 23820
rect 24213 23817 24225 23851
rect 24259 23848 24271 23851
rect 24946 23848 24952 23860
rect 24259 23820 24952 23848
rect 24259 23817 24271 23820
rect 24213 23811 24271 23817
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 26418 23848 26424 23860
rect 25056 23820 26424 23848
rect 25056 23780 25084 23820
rect 26418 23808 26424 23820
rect 26476 23808 26482 23860
rect 29365 23851 29423 23857
rect 29365 23848 29377 23851
rect 26620 23820 29377 23848
rect 24136 23752 25084 23780
rect 25133 23783 25191 23789
rect 25133 23749 25145 23783
rect 25179 23780 25191 23783
rect 25406 23780 25412 23792
rect 25179 23752 25412 23780
rect 25179 23749 25191 23752
rect 25133 23743 25191 23749
rect 25406 23740 25412 23752
rect 25464 23740 25470 23792
rect 26510 23780 26516 23792
rect 26358 23752 26516 23780
rect 26510 23740 26516 23752
rect 26568 23740 26574 23792
rect 15151 23684 16068 23712
rect 15151 23681 15163 23684
rect 15105 23675 15163 23681
rect 16850 23672 16856 23724
rect 16908 23672 16914 23724
rect 16942 23672 16948 23724
rect 17000 23712 17006 23724
rect 17000 23684 18000 23712
rect 17000 23672 17006 23684
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 6457 23647 6515 23653
rect 6457 23613 6469 23647
rect 6503 23644 6515 23647
rect 6503 23616 7328 23644
rect 6503 23613 6515 23616
rect 6457 23607 6515 23613
rect 1210 23536 1216 23588
rect 1268 23576 1274 23588
rect 6733 23579 6791 23585
rect 6733 23576 6745 23579
rect 1268 23548 2360 23576
rect 1268 23536 1274 23548
rect 1762 23468 1768 23520
rect 1820 23508 1826 23520
rect 2225 23511 2283 23517
rect 2225 23508 2237 23511
rect 1820 23480 2237 23508
rect 1820 23468 1826 23480
rect 2225 23477 2237 23480
rect 2271 23477 2283 23511
rect 2332 23508 2360 23548
rect 2746 23548 6745 23576
rect 2746 23508 2774 23548
rect 6733 23545 6745 23548
rect 6779 23545 6791 23579
rect 7300 23576 7328 23616
rect 7374 23604 7380 23656
rect 7432 23604 7438 23656
rect 12529 23647 12587 23653
rect 11532 23616 12434 23644
rect 11532 23576 11560 23616
rect 7300 23548 11560 23576
rect 12406 23576 12434 23616
rect 12529 23613 12541 23647
rect 12575 23644 12587 23647
rect 17034 23644 17040 23656
rect 12575 23616 17040 23644
rect 12575 23613 12587 23616
rect 12529 23607 12587 23613
rect 17034 23604 17040 23616
rect 17092 23604 17098 23656
rect 17862 23604 17868 23656
rect 17920 23604 17926 23656
rect 17972 23644 18000 23684
rect 18690 23672 18696 23724
rect 18748 23672 18754 23724
rect 20898 23672 20904 23724
rect 20956 23712 20962 23724
rect 20993 23715 21051 23721
rect 20993 23712 21005 23715
rect 20956 23684 21005 23712
rect 20956 23672 20962 23684
rect 20993 23681 21005 23684
rect 21039 23681 21051 23715
rect 26620 23712 26648 23820
rect 29365 23817 29377 23820
rect 29411 23817 29423 23851
rect 29365 23811 29423 23817
rect 29546 23808 29552 23860
rect 29604 23848 29610 23860
rect 33413 23851 33471 23857
rect 33413 23848 33425 23851
rect 29604 23820 33425 23848
rect 29604 23808 29610 23820
rect 33413 23817 33425 23820
rect 33459 23817 33471 23851
rect 33413 23811 33471 23817
rect 33594 23808 33600 23860
rect 33652 23848 33658 23860
rect 34057 23851 34115 23857
rect 34057 23848 34069 23851
rect 33652 23820 34069 23848
rect 33652 23808 33658 23820
rect 34057 23817 34069 23820
rect 34103 23817 34115 23851
rect 34057 23811 34115 23817
rect 34790 23808 34796 23860
rect 34848 23808 34854 23860
rect 38286 23848 38292 23860
rect 34900 23820 38292 23848
rect 27062 23740 27068 23792
rect 27120 23780 27126 23792
rect 27706 23780 27712 23792
rect 27120 23752 27712 23780
rect 27120 23740 27126 23752
rect 27706 23740 27712 23752
rect 27764 23740 27770 23792
rect 30098 23740 30104 23792
rect 30156 23740 30162 23792
rect 32858 23740 32864 23792
rect 32916 23780 32922 23792
rect 32953 23783 33011 23789
rect 32953 23780 32965 23783
rect 32916 23752 32965 23780
rect 32916 23740 32922 23752
rect 32953 23749 32965 23752
rect 32999 23749 33011 23783
rect 34900 23780 34928 23820
rect 38286 23808 38292 23820
rect 38344 23808 38350 23860
rect 38470 23808 38476 23860
rect 38528 23808 38534 23860
rect 39025 23851 39083 23857
rect 39025 23817 39037 23851
rect 39071 23848 39083 23851
rect 39206 23848 39212 23860
rect 39071 23820 39212 23848
rect 39071 23817 39083 23820
rect 39025 23811 39083 23817
rect 39206 23808 39212 23820
rect 39264 23808 39270 23860
rect 39574 23808 39580 23860
rect 39632 23848 39638 23860
rect 39853 23851 39911 23857
rect 39853 23848 39865 23851
rect 39632 23820 39865 23848
rect 39632 23808 39638 23820
rect 39853 23817 39865 23820
rect 39899 23817 39911 23851
rect 39853 23811 39911 23817
rect 40310 23808 40316 23860
rect 40368 23808 40374 23860
rect 40678 23808 40684 23860
rect 40736 23808 40742 23860
rect 45922 23808 45928 23860
rect 45980 23848 45986 23860
rect 46293 23851 46351 23857
rect 46293 23848 46305 23851
rect 45980 23820 46305 23848
rect 45980 23808 45986 23820
rect 46293 23817 46305 23820
rect 46339 23817 46351 23851
rect 46293 23811 46351 23817
rect 47302 23808 47308 23860
rect 47360 23848 47366 23860
rect 47581 23851 47639 23857
rect 47581 23848 47593 23851
rect 47360 23820 47593 23848
rect 47360 23808 47366 23820
rect 47581 23817 47593 23820
rect 47627 23817 47639 23851
rect 47581 23811 47639 23817
rect 32953 23743 33011 23749
rect 34440 23752 34928 23780
rect 34992 23752 35572 23780
rect 20993 23675 21051 23681
rect 26344 23684 26648 23712
rect 19518 23644 19524 23656
rect 17972 23616 19524 23644
rect 19518 23604 19524 23616
rect 19576 23604 19582 23656
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 20088 23616 22017 23644
rect 13722 23576 13728 23588
rect 12406 23548 13728 23576
rect 6733 23539 6791 23545
rect 13722 23536 13728 23548
rect 13780 23536 13786 23588
rect 20088 23520 20116 23616
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22370 23644 22376 23656
rect 22005 23607 22063 23613
rect 22112 23616 22376 23644
rect 21637 23579 21695 23585
rect 21637 23545 21649 23579
rect 21683 23576 21695 23579
rect 22112 23576 22140 23616
rect 22370 23604 22376 23616
rect 22428 23604 22434 23656
rect 22830 23604 22836 23656
rect 22888 23644 22894 23656
rect 24854 23644 24860 23656
rect 22888 23616 24860 23644
rect 22888 23604 22894 23616
rect 24854 23604 24860 23616
rect 24912 23604 24918 23656
rect 25130 23644 25136 23656
rect 24964 23616 25136 23644
rect 24964 23576 24992 23616
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 25774 23604 25780 23656
rect 25832 23644 25838 23656
rect 26344 23644 26372 23684
rect 28534 23672 28540 23724
rect 28592 23672 28598 23724
rect 29546 23672 29552 23724
rect 29604 23672 29610 23724
rect 30282 23672 30288 23724
rect 30340 23672 30346 23724
rect 30837 23715 30895 23721
rect 30837 23681 30849 23715
rect 30883 23712 30895 23715
rect 31021 23715 31079 23721
rect 31021 23712 31033 23715
rect 30883 23684 31033 23712
rect 30883 23681 30895 23684
rect 30837 23675 30895 23681
rect 31021 23681 31033 23684
rect 31067 23712 31079 23715
rect 31386 23712 31392 23724
rect 31067 23684 31392 23712
rect 31067 23681 31079 23684
rect 31021 23675 31079 23681
rect 31386 23672 31392 23684
rect 31444 23672 31450 23724
rect 31489 23719 31547 23725
rect 31489 23685 31501 23719
rect 31535 23716 31547 23719
rect 31535 23688 31616 23716
rect 31535 23685 31547 23688
rect 31489 23679 31547 23685
rect 27154 23644 27160 23656
rect 25832 23616 26372 23644
rect 26436 23616 27160 23644
rect 25832 23604 25838 23616
rect 21683 23548 22140 23576
rect 23308 23548 24992 23576
rect 21683 23545 21695 23548
rect 21637 23539 21695 23545
rect 2332 23480 2774 23508
rect 2225 23471 2283 23477
rect 6546 23468 6552 23520
rect 6604 23468 6610 23520
rect 9582 23468 9588 23520
rect 9640 23508 9646 23520
rect 11514 23508 11520 23520
rect 9640 23480 11520 23508
rect 9640 23468 9646 23480
rect 11514 23468 11520 23480
rect 11572 23468 11578 23520
rect 11606 23468 11612 23520
rect 11664 23508 11670 23520
rect 12710 23508 12716 23520
rect 11664 23480 12716 23508
rect 11664 23468 11670 23480
rect 12710 23468 12716 23480
rect 12768 23468 12774 23520
rect 13170 23468 13176 23520
rect 13228 23508 13234 23520
rect 17770 23508 17776 23520
rect 13228 23480 17776 23508
rect 13228 23468 13234 23480
rect 17770 23468 17776 23480
rect 17828 23468 17834 23520
rect 18690 23468 18696 23520
rect 18748 23508 18754 23520
rect 20070 23508 20076 23520
rect 18748 23480 20076 23508
rect 18748 23468 18754 23480
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 20438 23468 20444 23520
rect 20496 23468 20502 23520
rect 22278 23468 22284 23520
rect 22336 23508 22342 23520
rect 23308 23508 23336 23548
rect 22336 23480 23336 23508
rect 22336 23468 22342 23480
rect 23750 23468 23756 23520
rect 23808 23468 23814 23520
rect 24854 23468 24860 23520
rect 24912 23508 24918 23520
rect 26436 23508 26464 23616
rect 27154 23604 27160 23616
rect 27212 23604 27218 23656
rect 27433 23647 27491 23653
rect 27433 23644 27445 23647
rect 27264 23616 27445 23644
rect 27264 23576 27292 23616
rect 27433 23613 27445 23616
rect 27479 23613 27491 23647
rect 30558 23644 30564 23656
rect 27433 23607 27491 23613
rect 28460 23616 30564 23644
rect 26620 23548 27292 23576
rect 26620 23520 26648 23548
rect 24912 23480 26464 23508
rect 24912 23468 24918 23480
rect 26602 23468 26608 23520
rect 26660 23468 26666 23520
rect 27246 23468 27252 23520
rect 27304 23508 27310 23520
rect 28460 23508 28488 23616
rect 30558 23604 30564 23616
rect 30616 23604 30622 23656
rect 31588 23644 31616 23688
rect 32030 23672 32036 23724
rect 32088 23712 32094 23724
rect 33965 23715 34023 23721
rect 33965 23712 33977 23715
rect 32088 23684 33977 23712
rect 32088 23672 32094 23684
rect 33965 23681 33977 23684
rect 34011 23681 34023 23715
rect 33965 23675 34023 23681
rect 31662 23644 31668 23656
rect 31588 23616 31668 23644
rect 31662 23604 31668 23616
rect 31720 23604 31726 23656
rect 32214 23604 32220 23656
rect 32272 23644 32278 23656
rect 32309 23647 32367 23653
rect 32309 23644 32321 23647
rect 32272 23616 32321 23644
rect 32272 23604 32278 23616
rect 32309 23613 32321 23616
rect 32355 23613 32367 23647
rect 32309 23607 32367 23613
rect 30653 23579 30711 23585
rect 30653 23545 30665 23579
rect 30699 23576 30711 23579
rect 30834 23576 30840 23588
rect 30699 23548 30840 23576
rect 30699 23545 30711 23548
rect 30653 23539 30711 23545
rect 30834 23536 30840 23548
rect 30892 23536 30898 23588
rect 31018 23536 31024 23588
rect 31076 23576 31082 23588
rect 34440 23576 34468 23752
rect 34698 23672 34704 23724
rect 34756 23672 34762 23724
rect 34514 23604 34520 23656
rect 34572 23644 34578 23656
rect 34992 23644 35020 23752
rect 35437 23715 35495 23721
rect 35437 23681 35449 23715
rect 35483 23681 35495 23715
rect 35437 23675 35495 23681
rect 34572 23616 35020 23644
rect 34572 23604 34578 23616
rect 31076 23548 34468 23576
rect 31076 23536 31082 23548
rect 27304 23480 28488 23508
rect 27304 23468 27310 23480
rect 28810 23468 28816 23520
rect 28868 23508 28874 23520
rect 28905 23511 28963 23517
rect 28905 23508 28917 23511
rect 28868 23480 28917 23508
rect 28868 23468 28874 23480
rect 28905 23477 28917 23480
rect 28951 23477 28963 23511
rect 28905 23471 28963 23477
rect 31294 23468 31300 23520
rect 31352 23468 31358 23520
rect 31386 23468 31392 23520
rect 31444 23508 31450 23520
rect 31849 23511 31907 23517
rect 31849 23508 31861 23511
rect 31444 23480 31861 23508
rect 31444 23468 31450 23480
rect 31849 23477 31861 23480
rect 31895 23508 31907 23511
rect 32214 23508 32220 23520
rect 31895 23480 32220 23508
rect 31895 23477 31907 23480
rect 31849 23471 31907 23477
rect 32214 23468 32220 23480
rect 32272 23468 32278 23520
rect 32490 23468 32496 23520
rect 32548 23508 32554 23520
rect 35452 23508 35480 23675
rect 35544 23576 35572 23752
rect 35618 23740 35624 23792
rect 35676 23740 35682 23792
rect 35710 23740 35716 23792
rect 35768 23780 35774 23792
rect 38657 23783 38715 23789
rect 38657 23780 38669 23783
rect 35768 23752 38669 23780
rect 35768 23740 35774 23752
rect 38657 23749 38669 23752
rect 38703 23749 38715 23783
rect 38657 23743 38715 23749
rect 36262 23672 36268 23724
rect 36320 23672 36326 23724
rect 36354 23672 36360 23724
rect 36412 23712 36418 23724
rect 36909 23715 36967 23721
rect 36909 23712 36921 23715
rect 36412 23684 36921 23712
rect 36412 23672 36418 23684
rect 36909 23681 36921 23684
rect 36955 23712 36967 23715
rect 37277 23715 37335 23721
rect 37277 23712 37289 23715
rect 36955 23684 37289 23712
rect 36955 23681 36967 23684
rect 36909 23675 36967 23681
rect 37277 23681 37289 23684
rect 37323 23681 37335 23715
rect 37277 23675 37335 23681
rect 37642 23672 37648 23724
rect 37700 23712 37706 23724
rect 37921 23715 37979 23721
rect 37921 23712 37933 23715
rect 37700 23684 37933 23712
rect 37700 23672 37706 23684
rect 37921 23681 37933 23684
rect 37967 23712 37979 23715
rect 38197 23715 38255 23721
rect 38197 23712 38209 23715
rect 37967 23684 38209 23712
rect 37967 23681 37979 23684
rect 37921 23675 37979 23681
rect 38197 23681 38209 23684
rect 38243 23681 38255 23715
rect 40328 23712 40356 23808
rect 44174 23740 44180 23792
rect 44232 23780 44238 23792
rect 46201 23783 46259 23789
rect 46201 23780 46213 23783
rect 44232 23752 46213 23780
rect 44232 23740 44238 23752
rect 40865 23715 40923 23721
rect 40865 23712 40877 23715
rect 40328 23684 40877 23712
rect 38197 23675 38255 23681
rect 40865 23681 40877 23684
rect 40911 23681 40923 23715
rect 40865 23675 40923 23681
rect 40954 23672 40960 23724
rect 41012 23712 41018 23724
rect 41509 23715 41567 23721
rect 41509 23712 41521 23715
rect 41012 23684 41521 23712
rect 41012 23672 41018 23684
rect 41509 23681 41521 23684
rect 41555 23712 41567 23715
rect 41785 23715 41843 23721
rect 41785 23712 41797 23715
rect 41555 23684 41797 23712
rect 41555 23681 41567 23684
rect 41509 23675 41567 23681
rect 41785 23681 41797 23684
rect 41831 23681 41843 23715
rect 41785 23675 41843 23681
rect 42058 23672 42064 23724
rect 42116 23712 42122 23724
rect 42613 23715 42671 23721
rect 42613 23712 42625 23715
rect 42116 23684 42625 23712
rect 42116 23672 42122 23684
rect 42613 23681 42625 23684
rect 42659 23681 42671 23715
rect 42613 23675 42671 23681
rect 43714 23672 43720 23724
rect 43772 23672 43778 23724
rect 43806 23672 43812 23724
rect 43864 23712 43870 23724
rect 44634 23712 44640 23724
rect 43864 23684 44640 23712
rect 43864 23672 43870 23684
rect 44634 23672 44640 23684
rect 44692 23712 44698 23724
rect 45572 23721 45600 23752
rect 46201 23749 46213 23752
rect 46247 23749 46259 23783
rect 46201 23743 46259 23749
rect 44821 23715 44879 23721
rect 44821 23712 44833 23715
rect 44692 23684 44833 23712
rect 44692 23672 44698 23684
rect 44821 23681 44833 23684
rect 44867 23681 44879 23715
rect 44821 23675 44879 23681
rect 45557 23715 45615 23721
rect 45557 23681 45569 23715
rect 45603 23712 45615 23715
rect 45603 23684 45637 23712
rect 45603 23681 45615 23684
rect 45557 23675 45615 23681
rect 46658 23672 46664 23724
rect 46716 23712 46722 23724
rect 46753 23715 46811 23721
rect 46753 23712 46765 23715
rect 46716 23684 46765 23712
rect 46716 23672 46722 23684
rect 46753 23681 46765 23684
rect 46799 23712 46811 23715
rect 47305 23715 47363 23721
rect 47305 23712 47317 23715
rect 46799 23684 47317 23712
rect 46799 23681 46811 23684
rect 46753 23675 46811 23681
rect 47305 23681 47317 23684
rect 47351 23681 47363 23715
rect 47305 23675 47363 23681
rect 47762 23672 47768 23724
rect 47820 23712 47826 23724
rect 47949 23715 48007 23721
rect 47949 23712 47961 23715
rect 47820 23684 47961 23712
rect 47820 23672 47826 23684
rect 47949 23681 47961 23684
rect 47995 23712 48007 23715
rect 48314 23712 48320 23724
rect 47995 23684 48320 23712
rect 47995 23681 48007 23684
rect 47949 23675 48007 23681
rect 48314 23672 48320 23684
rect 48372 23672 48378 23724
rect 48682 23672 48688 23724
rect 48740 23672 48746 23724
rect 38562 23604 38568 23656
rect 38620 23644 38626 23656
rect 38620 23616 45048 23644
rect 38620 23604 38626 23616
rect 36725 23579 36783 23585
rect 36725 23576 36737 23579
rect 35544 23548 36737 23576
rect 36725 23545 36737 23548
rect 36771 23545 36783 23579
rect 36725 23539 36783 23545
rect 37182 23536 37188 23588
rect 37240 23576 37246 23588
rect 41325 23579 41383 23585
rect 41325 23576 41337 23579
rect 37240 23548 41337 23576
rect 37240 23536 37246 23548
rect 41325 23545 41337 23548
rect 41371 23545 41383 23579
rect 41325 23539 41383 23545
rect 41414 23536 41420 23588
rect 41472 23576 41478 23588
rect 45020 23585 45048 23616
rect 44361 23579 44419 23585
rect 44361 23576 44373 23579
rect 41472 23548 44373 23576
rect 41472 23536 41478 23548
rect 44361 23545 44373 23548
rect 44407 23545 44419 23579
rect 44361 23539 44419 23545
rect 45005 23579 45063 23585
rect 45005 23545 45017 23579
rect 45051 23545 45063 23579
rect 45005 23539 45063 23545
rect 32548 23480 35480 23508
rect 32548 23468 32554 23480
rect 36078 23468 36084 23520
rect 36136 23468 36142 23520
rect 37366 23468 37372 23520
rect 37424 23508 37430 23520
rect 37737 23511 37795 23517
rect 37737 23508 37749 23511
rect 37424 23480 37749 23508
rect 37424 23468 37430 23480
rect 37737 23477 37749 23480
rect 37783 23477 37795 23511
rect 37737 23471 37795 23477
rect 43257 23511 43315 23517
rect 43257 23477 43269 23511
rect 43303 23508 43315 23511
rect 43346 23508 43352 23520
rect 43303 23480 43352 23508
rect 43303 23477 43315 23480
rect 43257 23471 43315 23477
rect 43346 23468 43352 23480
rect 43404 23468 43410 23520
rect 45738 23468 45744 23520
rect 45796 23468 45802 23520
rect 46934 23468 46940 23520
rect 46992 23468 46998 23520
rect 47026 23468 47032 23520
rect 47084 23508 47090 23520
rect 48133 23511 48191 23517
rect 48133 23508 48145 23511
rect 47084 23480 48145 23508
rect 47084 23468 47090 23480
rect 48133 23477 48145 23480
rect 48179 23477 48191 23511
rect 48133 23471 48191 23477
rect 48682 23468 48688 23520
rect 48740 23508 48746 23520
rect 49329 23511 49387 23517
rect 49329 23508 49341 23511
rect 48740 23480 49341 23508
rect 48740 23468 48746 23480
rect 49329 23477 49341 23480
rect 49375 23477 49387 23511
rect 49329 23471 49387 23477
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 1854 23264 1860 23316
rect 1912 23304 1918 23316
rect 14461 23307 14519 23313
rect 14461 23304 14473 23307
rect 1912 23276 14473 23304
rect 1912 23264 1918 23276
rect 14461 23273 14473 23276
rect 14507 23273 14519 23307
rect 14461 23267 14519 23273
rect 17862 23264 17868 23316
rect 17920 23304 17926 23316
rect 19610 23304 19616 23316
rect 17920 23276 19616 23304
rect 17920 23264 17926 23276
rect 19610 23264 19616 23276
rect 19668 23264 19674 23316
rect 20336 23307 20394 23313
rect 20336 23273 20348 23307
rect 20382 23304 20394 23307
rect 21450 23304 21456 23316
rect 20382 23276 21456 23304
rect 20382 23273 20394 23276
rect 20336 23267 20394 23273
rect 21450 23264 21456 23276
rect 21508 23264 21514 23316
rect 22370 23264 22376 23316
rect 22428 23304 22434 23316
rect 23290 23304 23296 23316
rect 22428 23276 23296 23304
rect 22428 23264 22434 23276
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 23566 23264 23572 23316
rect 23624 23304 23630 23316
rect 25777 23307 25835 23313
rect 25777 23304 25789 23307
rect 23624 23276 25789 23304
rect 23624 23264 23630 23276
rect 25777 23273 25789 23276
rect 25823 23273 25835 23307
rect 25777 23267 25835 23273
rect 27512 23307 27570 23313
rect 27512 23273 27524 23307
rect 27558 23304 27570 23307
rect 28810 23304 28816 23316
rect 27558 23276 28816 23304
rect 27558 23273 27570 23276
rect 27512 23267 27570 23273
rect 28810 23264 28816 23276
rect 28868 23264 28874 23316
rect 28997 23307 29055 23313
rect 28997 23273 29009 23307
rect 29043 23304 29055 23307
rect 29086 23304 29092 23316
rect 29043 23276 29092 23304
rect 29043 23273 29055 23276
rect 28997 23267 29055 23273
rect 29086 23264 29092 23276
rect 29144 23304 29150 23316
rect 29990 23307 30048 23313
rect 29990 23304 30002 23307
rect 29144 23276 30002 23304
rect 29144 23264 29150 23276
rect 29990 23273 30002 23276
rect 30036 23273 30048 23307
rect 29990 23267 30048 23273
rect 31294 23264 31300 23316
rect 31352 23304 31358 23316
rect 33042 23304 33048 23316
rect 31352 23276 33048 23304
rect 31352 23264 31358 23276
rect 33042 23264 33048 23276
rect 33100 23264 33106 23316
rect 36262 23264 36268 23316
rect 36320 23304 36326 23316
rect 36633 23307 36691 23313
rect 36633 23304 36645 23307
rect 36320 23276 36645 23304
rect 36320 23264 36326 23276
rect 36633 23273 36645 23276
rect 36679 23273 36691 23307
rect 36633 23267 36691 23273
rect 36814 23264 36820 23316
rect 36872 23264 36878 23316
rect 37274 23264 37280 23316
rect 37332 23264 37338 23316
rect 43993 23307 44051 23313
rect 43993 23273 44005 23307
rect 44039 23304 44051 23307
rect 44358 23304 44364 23316
rect 44039 23276 44364 23304
rect 44039 23273 44051 23276
rect 43993 23267 44051 23273
rect 44358 23264 44364 23276
rect 44416 23264 44422 23316
rect 44634 23264 44640 23316
rect 44692 23264 44698 23316
rect 48590 23264 48596 23316
rect 48648 23304 48654 23316
rect 49329 23307 49387 23313
rect 49329 23304 49341 23307
rect 48648 23276 49341 23304
rect 48648 23264 48654 23276
rect 49329 23273 49341 23276
rect 49375 23273 49387 23307
rect 49329 23267 49387 23273
rect 2746 23208 7972 23236
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 2746 23100 2774 23208
rect 2866 23128 2872 23180
rect 2924 23168 2930 23180
rect 4338 23168 4344 23180
rect 2924 23140 4344 23168
rect 2924 23128 2930 23140
rect 4338 23128 4344 23140
rect 4396 23128 4402 23180
rect 4706 23128 4712 23180
rect 4764 23128 4770 23180
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 7944 23168 7972 23208
rect 12894 23196 12900 23248
rect 12952 23236 12958 23248
rect 13446 23236 13452 23248
rect 12952 23208 13452 23236
rect 12952 23196 12958 23208
rect 13446 23196 13452 23208
rect 13504 23196 13510 23248
rect 18874 23196 18880 23248
rect 18932 23196 18938 23248
rect 19334 23196 19340 23248
rect 19392 23236 19398 23248
rect 19392 23208 20208 23236
rect 19392 23196 19398 23208
rect 11422 23168 11428 23180
rect 7944 23140 11428 23168
rect 11422 23128 11428 23140
rect 11480 23128 11486 23180
rect 11517 23171 11575 23177
rect 11517 23137 11529 23171
rect 11563 23168 11575 23171
rect 12434 23168 12440 23180
rect 11563 23140 12440 23168
rect 11563 23137 11575 23140
rect 11517 23131 11575 23137
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 13265 23171 13323 23177
rect 13265 23137 13277 23171
rect 13311 23168 13323 23171
rect 13630 23168 13636 23180
rect 13311 23140 13636 23168
rect 13311 23137 13323 23140
rect 13265 23131 13323 23137
rect 13630 23128 13636 23140
rect 13688 23128 13694 23180
rect 16485 23171 16543 23177
rect 16485 23137 16497 23171
rect 16531 23168 16543 23171
rect 17402 23168 17408 23180
rect 16531 23140 17408 23168
rect 16531 23137 16543 23140
rect 16485 23131 16543 23137
rect 17402 23128 17408 23140
rect 17460 23128 17466 23180
rect 20070 23128 20076 23180
rect 20128 23128 20134 23180
rect 20180 23168 20208 23208
rect 23750 23196 23756 23248
rect 23808 23236 23814 23248
rect 23808 23208 25268 23236
rect 23808 23196 23814 23208
rect 21818 23168 21824 23180
rect 20180 23140 21824 23168
rect 21818 23128 21824 23140
rect 21876 23128 21882 23180
rect 22557 23171 22615 23177
rect 22557 23137 22569 23171
rect 22603 23168 22615 23171
rect 23768 23168 23796 23196
rect 22603 23140 23796 23168
rect 22603 23137 22615 23140
rect 22557 23131 22615 23137
rect 25130 23128 25136 23180
rect 25188 23128 25194 23180
rect 25240 23168 25268 23208
rect 25682 23196 25688 23248
rect 25740 23236 25746 23248
rect 26789 23239 26847 23245
rect 26789 23236 26801 23239
rect 25740 23208 26801 23236
rect 25740 23196 25746 23208
rect 26789 23205 26801 23208
rect 26835 23205 26847 23239
rect 26789 23199 26847 23205
rect 28626 23196 28632 23248
rect 28684 23196 28690 23248
rect 28718 23196 28724 23248
rect 28776 23236 28782 23248
rect 29730 23236 29736 23248
rect 28776 23208 29736 23236
rect 28776 23196 28782 23208
rect 29730 23196 29736 23208
rect 29788 23196 29794 23248
rect 32582 23196 32588 23248
rect 32640 23196 32646 23248
rect 33321 23239 33379 23245
rect 33321 23205 33333 23239
rect 33367 23236 33379 23239
rect 33502 23236 33508 23248
rect 33367 23208 33508 23236
rect 33367 23205 33379 23208
rect 33321 23199 33379 23205
rect 33502 23196 33508 23208
rect 33560 23196 33566 23248
rect 33686 23196 33692 23248
rect 33744 23236 33750 23248
rect 34057 23239 34115 23245
rect 34057 23236 34069 23239
rect 33744 23208 34069 23236
rect 33744 23196 33750 23208
rect 34057 23205 34069 23208
rect 34103 23205 34115 23239
rect 34057 23199 34115 23205
rect 34882 23196 34888 23248
rect 34940 23196 34946 23248
rect 34974 23196 34980 23248
rect 35032 23236 35038 23248
rect 37001 23239 37059 23245
rect 37001 23236 37013 23239
rect 35032 23208 37013 23236
rect 35032 23196 35038 23208
rect 37001 23205 37013 23208
rect 37047 23205 37059 23239
rect 37001 23199 37059 23205
rect 26329 23171 26387 23177
rect 26329 23168 26341 23171
rect 25240 23140 26341 23168
rect 26329 23137 26341 23140
rect 26375 23137 26387 23171
rect 26329 23131 26387 23137
rect 27154 23128 27160 23180
rect 27212 23168 27218 23180
rect 27249 23171 27307 23177
rect 27249 23168 27261 23171
rect 27212 23140 27261 23168
rect 27212 23128 27218 23140
rect 27249 23137 27261 23140
rect 27295 23168 27307 23171
rect 27614 23168 27620 23180
rect 27295 23140 27620 23168
rect 27295 23137 27307 23140
rect 27249 23131 27307 23137
rect 27614 23128 27620 23140
rect 27672 23128 27678 23180
rect 28644 23168 28672 23196
rect 31386 23168 31392 23180
rect 28644 23140 28856 23168
rect 1811 23072 2774 23100
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 3418 23060 3424 23112
rect 3476 23060 3482 23112
rect 3602 23060 3608 23112
rect 3660 23060 3666 23112
rect 4246 23060 4252 23112
rect 4304 23100 4310 23112
rect 5353 23103 5411 23109
rect 5353 23100 5365 23103
rect 4304 23072 5365 23100
rect 4304 23060 4310 23072
rect 5353 23069 5365 23072
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 7190 23060 7196 23112
rect 7248 23060 7254 23112
rect 8938 23060 8944 23112
rect 8996 23100 9002 23112
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 8996 23072 9321 23100
rect 8996 23060 9002 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 13906 23060 13912 23112
rect 13964 23060 13970 23112
rect 14366 23060 14372 23112
rect 14424 23060 14430 23112
rect 15470 23060 15476 23112
rect 15528 23060 15534 23112
rect 16850 23060 16856 23112
rect 16908 23100 16914 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 16908 23072 17141 23100
rect 16908 23060 16914 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23100 19671 23103
rect 19978 23100 19984 23112
rect 19659 23072 19984 23100
rect 19659 23069 19671 23072
rect 19613 23063 19671 23069
rect 19978 23060 19984 23072
rect 20036 23060 20042 23112
rect 21910 23060 21916 23112
rect 21968 23100 21974 23112
rect 22281 23103 22339 23109
rect 22281 23100 22293 23103
rect 21968 23072 22293 23100
rect 21968 23060 21974 23072
rect 22281 23069 22293 23072
rect 22327 23069 22339 23103
rect 22281 23063 22339 23069
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23100 25007 23103
rect 25038 23100 25044 23112
rect 24995 23072 25044 23100
rect 24995 23069 25007 23072
rect 24949 23063 25007 23069
rect 25038 23060 25044 23072
rect 25096 23060 25102 23112
rect 26160 23072 27016 23100
rect 2774 22992 2780 23044
rect 2832 22992 2838 23044
rect 3510 22992 3516 23044
rect 3568 23032 3574 23044
rect 3789 23035 3847 23041
rect 3789 23032 3801 23035
rect 3568 23004 3801 23032
rect 3568 22992 3574 23004
rect 3789 23001 3801 23004
rect 3835 23001 3847 23035
rect 3789 22995 3847 23001
rect 4065 23035 4123 23041
rect 4065 23001 4077 23035
rect 4111 23032 4123 23035
rect 4111 23004 4568 23032
rect 4111 23001 4123 23004
rect 4065 22995 4123 23001
rect 4540 22976 4568 23004
rect 8846 22992 8852 23044
rect 8904 23032 8910 23044
rect 8904 23004 9536 23032
rect 8904 22992 8910 23004
rect 4154 22924 4160 22976
rect 4212 22924 4218 22976
rect 4522 22924 4528 22976
rect 4580 22924 4586 22976
rect 4617 22967 4675 22973
rect 4617 22933 4629 22967
rect 4663 22964 4675 22967
rect 6270 22964 6276 22976
rect 4663 22936 6276 22964
rect 4663 22933 4675 22936
rect 4617 22927 4675 22933
rect 6270 22924 6276 22936
rect 6328 22924 6334 22976
rect 9030 22924 9036 22976
rect 9088 22964 9094 22976
rect 9398 22964 9404 22976
rect 9088 22936 9404 22964
rect 9088 22924 9094 22936
rect 9398 22924 9404 22936
rect 9456 22924 9462 22976
rect 9508 22964 9536 23004
rect 9582 22992 9588 23044
rect 9640 22992 9646 23044
rect 9674 22992 9680 23044
rect 9732 23032 9738 23044
rect 11793 23035 11851 23041
rect 11793 23032 11805 23035
rect 9732 23004 10074 23032
rect 11624 23004 11805 23032
rect 9732 22992 9738 23004
rect 11057 22967 11115 22973
rect 11057 22964 11069 22967
rect 9508 22936 11069 22964
rect 11057 22933 11069 22936
rect 11103 22964 11115 22967
rect 11624 22964 11652 23004
rect 11793 23001 11805 23004
rect 11839 23001 11851 23035
rect 11793 22995 11851 23001
rect 12250 22992 12256 23044
rect 12308 22992 12314 23044
rect 17034 22992 17040 23044
rect 17092 23032 17098 23044
rect 17405 23035 17463 23041
rect 17405 23032 17417 23035
rect 17092 23004 17417 23032
rect 17092 22992 17098 23004
rect 17405 23001 17417 23004
rect 17451 23001 17463 23035
rect 19058 23032 19064 23044
rect 18630 23004 19064 23032
rect 17405 22995 17463 23001
rect 19058 22992 19064 23004
rect 19116 22992 19122 23044
rect 21358 22992 21364 23044
rect 21416 22992 21422 23044
rect 23290 22992 23296 23044
rect 23348 22992 23354 23044
rect 26160 23032 26188 23072
rect 23860 23004 24624 23032
rect 11103 22936 11652 22964
rect 11103 22933 11115 22936
rect 11057 22927 11115 22933
rect 11698 22924 11704 22976
rect 11756 22964 11762 22976
rect 12618 22964 12624 22976
rect 11756 22936 12624 22964
rect 11756 22924 11762 22936
rect 12618 22924 12624 22936
rect 12676 22924 12682 22976
rect 12802 22924 12808 22976
rect 12860 22964 12866 22976
rect 13633 22967 13691 22973
rect 13633 22964 13645 22967
rect 12860 22936 13645 22964
rect 12860 22924 12866 22936
rect 13633 22933 13645 22936
rect 13679 22964 13691 22967
rect 14550 22964 14556 22976
rect 13679 22936 14556 22964
rect 13679 22933 13691 22936
rect 13633 22927 13691 22933
rect 14550 22924 14556 22936
rect 14608 22964 14614 22976
rect 14921 22967 14979 22973
rect 14921 22964 14933 22967
rect 14608 22936 14933 22964
rect 14608 22924 14614 22936
rect 14921 22933 14933 22936
rect 14967 22933 14979 22967
rect 14921 22927 14979 22933
rect 15470 22924 15476 22976
rect 15528 22964 15534 22976
rect 19334 22964 19340 22976
rect 15528 22936 19340 22964
rect 15528 22924 15534 22936
rect 19334 22924 19340 22936
rect 19392 22924 19398 22976
rect 19429 22967 19487 22973
rect 19429 22933 19441 22967
rect 19475 22964 19487 22967
rect 20622 22964 20628 22976
rect 19475 22936 20628 22964
rect 19475 22933 19487 22936
rect 19429 22927 19487 22933
rect 20622 22924 20628 22936
rect 20680 22924 20686 22976
rect 21082 22924 21088 22976
rect 21140 22964 21146 22976
rect 23860 22964 23888 23004
rect 21140 22936 23888 22964
rect 21140 22924 21146 22936
rect 23934 22924 23940 22976
rect 23992 22964 23998 22976
rect 24596 22973 24624 23004
rect 25056 23004 26188 23032
rect 26237 23035 26295 23041
rect 25056 22973 25084 23004
rect 26237 23001 26249 23035
rect 26283 23032 26295 23035
rect 26988 23032 27016 23072
rect 28534 23060 28540 23112
rect 28592 23100 28598 23112
rect 28592 23086 28658 23100
rect 28592 23072 28672 23086
rect 28592 23060 28598 23072
rect 27798 23032 27804 23044
rect 26283 23004 26924 23032
rect 26988 23004 27804 23032
rect 26283 23001 26295 23004
rect 26237 22995 26295 23001
rect 24029 22967 24087 22973
rect 24029 22964 24041 22967
rect 23992 22936 24041 22964
rect 23992 22924 23998 22936
rect 24029 22933 24041 22936
rect 24075 22933 24087 22967
rect 24029 22927 24087 22933
rect 24581 22967 24639 22973
rect 24581 22933 24593 22967
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 25041 22967 25099 22973
rect 25041 22933 25053 22967
rect 25087 22933 25099 22967
rect 25041 22927 25099 22933
rect 25958 22924 25964 22976
rect 26016 22964 26022 22976
rect 26145 22967 26203 22973
rect 26145 22964 26157 22967
rect 26016 22936 26157 22964
rect 26016 22924 26022 22936
rect 26145 22933 26157 22936
rect 26191 22933 26203 22967
rect 26896 22964 26924 23004
rect 27798 22992 27804 23004
rect 27856 22992 27862 23044
rect 28350 22964 28356 22976
rect 26896 22936 28356 22964
rect 26145 22927 26203 22933
rect 28350 22924 28356 22936
rect 28408 22924 28414 22976
rect 28644 22964 28672 23072
rect 28828 23032 28856 23140
rect 29748 23140 31392 23168
rect 28902 23060 28908 23112
rect 28960 23100 28966 23112
rect 29748 23109 29776 23140
rect 31386 23128 31392 23140
rect 31444 23128 31450 23180
rect 31938 23128 31944 23180
rect 31996 23168 32002 23180
rect 36078 23168 36084 23180
rect 31996 23140 36084 23168
rect 31996 23128 32002 23140
rect 36078 23128 36084 23140
rect 36136 23128 36142 23180
rect 47489 23171 47547 23177
rect 47489 23137 47501 23171
rect 47535 23168 47547 23171
rect 47535 23140 48544 23168
rect 47535 23137 47547 23140
rect 47489 23131 47547 23137
rect 31726 23112 31892 23116
rect 48516 23112 48544 23140
rect 29733 23103 29791 23109
rect 29733 23100 29745 23103
rect 28960 23072 29745 23100
rect 28960 23060 28966 23072
rect 29733 23069 29745 23072
rect 29779 23069 29791 23103
rect 31478 23100 31484 23112
rect 31142 23072 31484 23100
rect 29733 23063 29791 23069
rect 31478 23060 31484 23072
rect 31536 23100 31542 23112
rect 31726 23100 31852 23112
rect 31536 23088 31852 23100
rect 31536 23072 31754 23088
rect 31536 23060 31542 23072
rect 31846 23060 31852 23088
rect 31904 23100 31910 23112
rect 31904 23072 32996 23100
rect 31904 23060 31910 23072
rect 30282 23032 30288 23044
rect 28828 23004 30288 23032
rect 30282 22992 30288 23004
rect 30340 22992 30346 23044
rect 32398 22992 32404 23044
rect 32456 22992 32462 23044
rect 32968 22976 32996 23072
rect 35066 23060 35072 23112
rect 35124 23060 35130 23112
rect 35710 23060 35716 23112
rect 35768 23060 35774 23112
rect 41141 23103 41199 23109
rect 41141 23069 41153 23103
rect 41187 23100 41199 23103
rect 41414 23100 41420 23112
rect 41187 23072 41420 23100
rect 41187 23069 41199 23072
rect 41141 23063 41199 23069
rect 41414 23060 41420 23072
rect 41472 23060 41478 23112
rect 43346 23060 43352 23112
rect 43404 23060 43410 23112
rect 47673 23103 47731 23109
rect 47673 23069 47685 23103
rect 47719 23100 47731 23103
rect 47854 23100 47860 23112
rect 47719 23072 47860 23100
rect 47719 23069 47731 23072
rect 47673 23063 47731 23069
rect 47854 23060 47860 23072
rect 47912 23100 47918 23112
rect 47949 23103 48007 23109
rect 47949 23100 47961 23103
rect 47912 23072 47961 23100
rect 47912 23060 47918 23072
rect 47949 23069 47961 23072
rect 47995 23069 48007 23103
rect 47949 23063 48007 23069
rect 48498 23060 48504 23112
rect 48556 23100 48562 23112
rect 48685 23103 48743 23109
rect 48685 23100 48697 23103
rect 48556 23072 48697 23100
rect 48556 23060 48562 23072
rect 48685 23069 48697 23072
rect 48731 23069 48743 23103
rect 48685 23063 48743 23069
rect 33137 23035 33195 23041
rect 33137 23001 33149 23035
rect 33183 23032 33195 23035
rect 33318 23032 33324 23044
rect 33183 23004 33324 23032
rect 33183 23001 33195 23004
rect 33137 22995 33195 23001
rect 33318 22992 33324 23004
rect 33376 22992 33382 23044
rect 33502 22992 33508 23044
rect 33560 23032 33566 23044
rect 33873 23035 33931 23041
rect 33873 23032 33885 23035
rect 33560 23004 33885 23032
rect 33560 22992 33566 23004
rect 33873 23001 33885 23004
rect 33919 23001 33931 23035
rect 33873 22995 33931 23001
rect 34425 23035 34483 23041
rect 34425 23001 34437 23035
rect 34471 23032 34483 23035
rect 34471 23004 39988 23032
rect 34471 23001 34483 23004
rect 34425 22995 34483 23001
rect 29365 22967 29423 22973
rect 29365 22964 29377 22967
rect 28644 22936 29377 22964
rect 29365 22933 29377 22936
rect 29411 22964 29423 22967
rect 29822 22964 29828 22976
rect 29411 22936 29828 22964
rect 29411 22933 29423 22936
rect 29365 22927 29423 22933
rect 29822 22924 29828 22936
rect 29880 22924 29886 22976
rect 30834 22924 30840 22976
rect 30892 22964 30898 22976
rect 31481 22967 31539 22973
rect 31481 22964 31493 22967
rect 30892 22936 31493 22964
rect 30892 22924 30898 22936
rect 31481 22933 31493 22936
rect 31527 22933 31539 22967
rect 31481 22927 31539 22933
rect 31846 22924 31852 22976
rect 31904 22964 31910 22976
rect 31941 22967 31999 22973
rect 31941 22964 31953 22967
rect 31904 22936 31953 22964
rect 31904 22924 31910 22936
rect 31941 22933 31953 22936
rect 31987 22933 31999 22967
rect 31941 22927 31999 22933
rect 32950 22924 32956 22976
rect 33008 22964 33014 22976
rect 34440 22964 34468 22995
rect 39960 22976 39988 23004
rect 33008 22936 34468 22964
rect 33008 22924 33014 22936
rect 35526 22924 35532 22976
rect 35584 22924 35590 22976
rect 36170 22924 36176 22976
rect 36228 22924 36234 22976
rect 39942 22924 39948 22976
rect 40000 22964 40006 22976
rect 42429 22967 42487 22973
rect 42429 22964 42441 22967
rect 40000 22936 42441 22964
rect 40000 22924 40006 22936
rect 42429 22933 42441 22936
rect 42475 22933 42487 22967
rect 42429 22927 42487 22933
rect 47486 22924 47492 22976
rect 47544 22964 47550 22976
rect 48133 22967 48191 22973
rect 48133 22964 48145 22967
rect 47544 22936 48145 22964
rect 47544 22924 47550 22936
rect 48133 22933 48145 22936
rect 48179 22933 48191 22967
rect 48133 22927 48191 22933
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 1026 22720 1032 22772
rect 1084 22760 1090 22772
rect 3789 22763 3847 22769
rect 3789 22760 3801 22763
rect 1084 22732 3801 22760
rect 1084 22720 1090 22732
rect 3789 22729 3801 22732
rect 3835 22729 3847 22763
rect 3789 22723 3847 22729
rect 6457 22763 6515 22769
rect 6457 22729 6469 22763
rect 6503 22760 6515 22763
rect 11790 22760 11796 22772
rect 6503 22732 11796 22760
rect 6503 22729 6515 22732
rect 6457 22723 6515 22729
rect 11790 22720 11796 22732
rect 11848 22720 11854 22772
rect 11882 22720 11888 22772
rect 11940 22760 11946 22772
rect 12526 22760 12532 22772
rect 11940 22732 12532 22760
rect 11940 22720 11946 22732
rect 12526 22720 12532 22732
rect 12584 22720 12590 22772
rect 13630 22760 13636 22772
rect 12728 22732 13636 22760
rect 1946 22652 1952 22704
rect 2004 22692 2010 22704
rect 2004 22664 5212 22692
rect 2004 22652 2010 22664
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 1854 22624 1860 22636
rect 1811 22596 1860 22624
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 4246 22624 4252 22636
rect 1964 22596 4252 22624
rect 1118 22516 1124 22568
rect 1176 22556 1182 22568
rect 1964 22556 1992 22596
rect 4246 22584 4252 22596
rect 4304 22584 4310 22636
rect 4798 22584 4804 22636
rect 4856 22584 4862 22636
rect 1176 22528 1992 22556
rect 2777 22559 2835 22565
rect 1176 22516 1182 22528
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 2866 22556 2872 22568
rect 2823 22528 2872 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 3510 22516 3516 22568
rect 3568 22556 3574 22568
rect 3881 22559 3939 22565
rect 3881 22556 3893 22559
rect 3568 22528 3893 22556
rect 3568 22516 3574 22528
rect 3881 22525 3893 22528
rect 3927 22525 3939 22559
rect 3881 22519 3939 22525
rect 4065 22559 4123 22565
rect 4065 22525 4077 22559
rect 4111 22525 4123 22559
rect 4065 22519 4123 22525
rect 2590 22380 2596 22432
rect 2648 22420 2654 22432
rect 3421 22423 3479 22429
rect 3421 22420 3433 22423
rect 2648 22392 3433 22420
rect 2648 22380 2654 22392
rect 3421 22389 3433 22392
rect 3467 22389 3479 22423
rect 4080 22420 4108 22519
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 5184 22556 5212 22664
rect 6730 22652 6736 22704
rect 6788 22692 6794 22704
rect 7926 22692 7932 22704
rect 6788 22664 7932 22692
rect 6788 22652 6794 22664
rect 7926 22652 7932 22664
rect 7984 22652 7990 22704
rect 10686 22652 10692 22704
rect 10744 22652 10750 22704
rect 12728 22701 12756 22732
rect 13630 22720 13636 22732
rect 13688 22720 13694 22772
rect 14550 22720 14556 22772
rect 14608 22720 14614 22772
rect 18601 22763 18659 22769
rect 18601 22729 18613 22763
rect 18647 22760 18659 22763
rect 18782 22760 18788 22772
rect 18647 22732 18788 22760
rect 18647 22729 18659 22732
rect 18601 22723 18659 22729
rect 18782 22720 18788 22732
rect 18840 22720 18846 22772
rect 19058 22720 19064 22772
rect 19116 22760 19122 22772
rect 19116 22732 21312 22760
rect 19116 22720 19122 22732
rect 12713 22695 12771 22701
rect 12713 22661 12725 22695
rect 12759 22661 12771 22695
rect 12713 22655 12771 22661
rect 12802 22652 12808 22704
rect 12860 22692 12866 22704
rect 12860 22664 13202 22692
rect 12860 22652 12866 22664
rect 16114 22652 16120 22704
rect 16172 22652 16178 22704
rect 16758 22652 16764 22704
rect 16816 22692 16822 22704
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 16816 22664 17141 22692
rect 16816 22652 16822 22664
rect 17129 22661 17141 22664
rect 17175 22661 17187 22695
rect 20070 22692 20076 22704
rect 17129 22655 17187 22661
rect 19720 22664 20076 22692
rect 6822 22584 6828 22636
rect 6880 22624 6886 22636
rect 7101 22627 7159 22633
rect 7101 22624 7113 22627
rect 6880 22596 7113 22624
rect 6880 22584 6886 22596
rect 7101 22593 7113 22596
rect 7147 22593 7159 22627
rect 7101 22587 7159 22593
rect 7193 22627 7251 22633
rect 7193 22593 7205 22627
rect 7239 22624 7251 22627
rect 7834 22624 7840 22636
rect 7239 22596 7840 22624
rect 7239 22593 7251 22596
rect 7193 22587 7251 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 8113 22627 8171 22633
rect 8113 22593 8125 22627
rect 8159 22624 8171 22627
rect 8294 22624 8300 22636
rect 8159 22596 8300 22624
rect 8159 22593 8171 22596
rect 8113 22587 8171 22593
rect 8294 22584 8300 22596
rect 8352 22584 8358 22636
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22624 10011 22627
rect 10042 22624 10048 22636
rect 9999 22596 10048 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 10042 22584 10048 22596
rect 10100 22584 10106 22636
rect 11790 22584 11796 22636
rect 11848 22584 11854 22636
rect 15010 22584 15016 22636
rect 15068 22584 15074 22636
rect 5184 22528 6868 22556
rect 5994 22448 6000 22500
rect 6052 22488 6058 22500
rect 6733 22491 6791 22497
rect 6733 22488 6745 22491
rect 6052 22460 6745 22488
rect 6052 22448 6058 22460
rect 6733 22457 6745 22460
rect 6779 22457 6791 22491
rect 6840 22488 6868 22528
rect 7006 22516 7012 22568
rect 7064 22556 7070 22568
rect 7285 22559 7343 22565
rect 7285 22556 7297 22559
rect 7064 22528 7297 22556
rect 7064 22516 7070 22528
rect 7285 22525 7297 22528
rect 7331 22525 7343 22559
rect 7285 22519 7343 22525
rect 8662 22516 8668 22568
rect 8720 22516 8726 22568
rect 12437 22559 12495 22565
rect 12437 22525 12449 22559
rect 12483 22525 12495 22559
rect 12437 22519 12495 22525
rect 11977 22491 12035 22497
rect 11977 22488 11989 22491
rect 6840 22460 11989 22488
rect 6733 22451 6791 22457
rect 11977 22457 11989 22460
rect 12023 22457 12035 22491
rect 12452 22488 12480 22519
rect 16850 22516 16856 22568
rect 16908 22516 16914 22568
rect 18138 22516 18144 22568
rect 18196 22556 18202 22568
rect 18248 22556 18276 22610
rect 18506 22584 18512 22636
rect 18564 22624 18570 22636
rect 19245 22627 19303 22633
rect 19245 22624 19257 22627
rect 18564 22596 19257 22624
rect 18564 22584 18570 22596
rect 19245 22593 19257 22596
rect 19291 22593 19303 22627
rect 19245 22587 19303 22593
rect 19426 22584 19432 22636
rect 19484 22624 19490 22636
rect 19720 22633 19748 22664
rect 20070 22652 20076 22664
rect 20128 22652 20134 22704
rect 21284 22692 21312 22732
rect 21450 22720 21456 22772
rect 21508 22760 21514 22772
rect 25130 22760 25136 22772
rect 21508 22732 25136 22760
rect 21508 22720 21514 22732
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 25682 22720 25688 22772
rect 25740 22720 25746 22772
rect 25774 22720 25780 22772
rect 25832 22720 25838 22772
rect 27157 22763 27215 22769
rect 27157 22729 27169 22763
rect 27203 22729 27215 22763
rect 27157 22723 27215 22729
rect 21358 22692 21364 22704
rect 21206 22664 21364 22692
rect 21358 22652 21364 22664
rect 21416 22692 21422 22704
rect 22189 22695 22247 22701
rect 22189 22692 22201 22695
rect 21416 22664 22201 22692
rect 21416 22652 21422 22664
rect 22189 22661 22201 22664
rect 22235 22692 22247 22695
rect 22370 22692 22376 22704
rect 22235 22664 22376 22692
rect 22235 22661 22247 22664
rect 22189 22655 22247 22661
rect 22370 22652 22376 22664
rect 22428 22652 22434 22704
rect 22465 22695 22523 22701
rect 22465 22661 22477 22695
rect 22511 22692 22523 22695
rect 23658 22692 23664 22704
rect 22511 22664 23664 22692
rect 22511 22661 22523 22664
rect 22465 22655 22523 22661
rect 23658 22652 23664 22664
rect 23716 22652 23722 22704
rect 24394 22652 24400 22704
rect 24452 22652 24458 22704
rect 24762 22652 24768 22704
rect 24820 22692 24826 22704
rect 27172 22692 27200 22723
rect 28810 22720 28816 22772
rect 28868 22760 28874 22772
rect 28868 22732 29960 22760
rect 28868 22720 28874 22732
rect 24820 22664 27200 22692
rect 24820 22652 24826 22664
rect 27614 22652 27620 22704
rect 27672 22652 27678 22704
rect 28626 22652 28632 22704
rect 28684 22692 28690 22704
rect 29932 22692 29960 22732
rect 30558 22720 30564 22772
rect 30616 22720 30622 22772
rect 32950 22720 32956 22772
rect 33008 22720 33014 22772
rect 33042 22720 33048 22772
rect 33100 22760 33106 22772
rect 33229 22763 33287 22769
rect 33229 22760 33241 22763
rect 33100 22732 33241 22760
rect 33100 22720 33106 22732
rect 33229 22729 33241 22732
rect 33275 22729 33287 22763
rect 33229 22723 33287 22729
rect 34698 22720 34704 22772
rect 34756 22760 34762 22772
rect 35066 22760 35072 22772
rect 34756 22732 35072 22760
rect 34756 22720 34762 22732
rect 35066 22720 35072 22732
rect 35124 22720 35130 22772
rect 39942 22720 39948 22772
rect 40000 22720 40006 22772
rect 47762 22720 47768 22772
rect 47820 22720 47826 22772
rect 31665 22695 31723 22701
rect 28684 22664 29118 22692
rect 29932 22664 31156 22692
rect 28684 22652 28690 22664
rect 19705 22627 19763 22633
rect 19705 22624 19717 22627
rect 19484 22596 19717 22624
rect 19484 22584 19490 22596
rect 19705 22593 19717 22596
rect 19751 22593 19763 22627
rect 19705 22587 19763 22593
rect 21910 22584 21916 22636
rect 21968 22624 21974 22636
rect 22830 22624 22836 22636
rect 21968 22596 22836 22624
rect 21968 22584 21974 22596
rect 22830 22584 22836 22596
rect 22888 22624 22894 22636
rect 23109 22627 23167 22633
rect 23109 22624 23121 22627
rect 22888 22596 23121 22624
rect 22888 22584 22894 22596
rect 23109 22593 23121 22596
rect 23155 22593 23167 22627
rect 26602 22624 26608 22636
rect 23109 22587 23167 22593
rect 25792 22596 26608 22624
rect 19058 22556 19064 22568
rect 18196 22528 19064 22556
rect 18196 22516 18202 22528
rect 19058 22516 19064 22528
rect 19116 22516 19122 22568
rect 19981 22559 20039 22565
rect 19981 22525 19993 22559
rect 20027 22556 20039 22559
rect 20070 22556 20076 22568
rect 20027 22528 20076 22556
rect 20027 22525 20039 22528
rect 19981 22519 20039 22525
rect 20070 22516 20076 22528
rect 20128 22556 20134 22568
rect 20438 22556 20444 22568
rect 20128 22528 20444 22556
rect 20128 22516 20134 22528
rect 20438 22516 20444 22528
rect 20496 22516 20502 22568
rect 22646 22516 22652 22568
rect 22704 22556 22710 22568
rect 23385 22559 23443 22565
rect 23385 22556 23397 22559
rect 22704 22528 23397 22556
rect 22704 22516 22710 22528
rect 23385 22525 23397 22528
rect 23431 22556 23443 22559
rect 23934 22556 23940 22568
rect 23431 22528 23940 22556
rect 23431 22525 23443 22528
rect 23385 22519 23443 22525
rect 23934 22516 23940 22528
rect 23992 22516 23998 22568
rect 25130 22516 25136 22568
rect 25188 22556 25194 22568
rect 25792 22556 25820 22596
rect 26602 22584 26608 22596
rect 26660 22584 26666 22636
rect 27338 22624 27344 22636
rect 26712 22596 27344 22624
rect 25188 22528 25820 22556
rect 25869 22559 25927 22565
rect 25188 22516 25194 22528
rect 25869 22525 25881 22559
rect 25915 22525 25927 22559
rect 25869 22519 25927 22525
rect 25884 22488 25912 22519
rect 25958 22516 25964 22568
rect 26016 22556 26022 22568
rect 26418 22556 26424 22568
rect 26016 22528 26424 22556
rect 26016 22516 26022 22528
rect 26418 22516 26424 22528
rect 26476 22556 26482 22568
rect 26712 22565 26740 22596
rect 27338 22584 27344 22596
rect 27396 22624 27402 22636
rect 27525 22627 27583 22633
rect 27525 22624 27537 22627
rect 27396 22596 27537 22624
rect 27396 22584 27402 22596
rect 27525 22593 27537 22596
rect 27571 22593 27583 22627
rect 27632 22624 27660 22652
rect 28353 22627 28411 22633
rect 28353 22624 28365 22627
rect 27632 22596 28365 22624
rect 27525 22587 27583 22593
rect 28353 22593 28365 22596
rect 28399 22593 28411 22627
rect 28353 22587 28411 22593
rect 30926 22584 30932 22636
rect 30984 22584 30990 22636
rect 26513 22559 26571 22565
rect 26513 22556 26525 22559
rect 26476 22528 26525 22556
rect 26476 22516 26482 22528
rect 26513 22525 26525 22528
rect 26559 22556 26571 22559
rect 26697 22559 26755 22565
rect 26697 22556 26709 22559
rect 26559 22528 26709 22556
rect 26559 22525 26571 22528
rect 26513 22519 26571 22525
rect 26697 22525 26709 22528
rect 26743 22525 26755 22559
rect 26697 22519 26755 22525
rect 27246 22516 27252 22568
rect 27304 22556 27310 22568
rect 27617 22559 27675 22565
rect 27617 22556 27629 22559
rect 27304 22528 27629 22556
rect 27304 22516 27310 22528
rect 27617 22525 27629 22528
rect 27663 22525 27675 22559
rect 27617 22519 27675 22525
rect 27709 22559 27767 22565
rect 27709 22525 27721 22559
rect 27755 22525 27767 22559
rect 27709 22519 27767 22525
rect 28629 22559 28687 22565
rect 28629 22525 28641 22559
rect 28675 22556 28687 22559
rect 30834 22556 30840 22568
rect 28675 22528 30840 22556
rect 28675 22525 28687 22528
rect 28629 22519 28687 22525
rect 12452 22460 12572 22488
rect 11977 22451 12035 22457
rect 6362 22420 6368 22432
rect 4080 22392 6368 22420
rect 3421 22383 3479 22389
rect 6362 22380 6368 22392
rect 6420 22380 6426 22432
rect 7098 22380 7104 22432
rect 7156 22420 7162 22432
rect 10042 22420 10048 22432
rect 7156 22392 10048 22420
rect 7156 22380 7162 22392
rect 10042 22380 10048 22392
rect 10100 22380 10106 22432
rect 12434 22380 12440 22432
rect 12492 22420 12498 22432
rect 12544 22420 12572 22460
rect 21008 22460 22784 22488
rect 12492 22392 12572 22420
rect 12492 22380 12498 22392
rect 13446 22380 13452 22432
rect 13504 22420 13510 22432
rect 14185 22423 14243 22429
rect 14185 22420 14197 22423
rect 13504 22392 14197 22420
rect 13504 22380 13510 22392
rect 14185 22389 14197 22392
rect 14231 22389 14243 22423
rect 14185 22383 14243 22389
rect 18690 22380 18696 22432
rect 18748 22420 18754 22432
rect 19061 22423 19119 22429
rect 19061 22420 19073 22423
rect 18748 22392 19073 22420
rect 18748 22380 18754 22392
rect 19061 22389 19073 22392
rect 19107 22389 19119 22423
rect 19061 22383 19119 22389
rect 19242 22380 19248 22432
rect 19300 22420 19306 22432
rect 21008 22420 21036 22460
rect 19300 22392 21036 22420
rect 19300 22380 19306 22392
rect 21910 22380 21916 22432
rect 21968 22380 21974 22432
rect 22756 22420 22784 22460
rect 24872 22460 25912 22488
rect 26252 22460 27384 22488
rect 23474 22420 23480 22432
rect 22756 22392 23480 22420
rect 23474 22380 23480 22392
rect 23532 22380 23538 22432
rect 23934 22380 23940 22432
rect 23992 22420 23998 22432
rect 24872 22429 24900 22460
rect 26252 22432 26280 22460
rect 24857 22423 24915 22429
rect 24857 22420 24869 22423
rect 23992 22392 24869 22420
rect 23992 22380 23998 22392
rect 24857 22389 24869 22392
rect 24903 22389 24915 22423
rect 24857 22383 24915 22389
rect 25314 22380 25320 22432
rect 25372 22380 25378 22432
rect 25682 22380 25688 22432
rect 25740 22420 25746 22432
rect 26234 22420 26240 22432
rect 25740 22392 26240 22420
rect 25740 22380 25746 22392
rect 26234 22380 26240 22392
rect 26292 22380 26298 22432
rect 26421 22423 26479 22429
rect 26421 22389 26433 22423
rect 26467 22420 26479 22423
rect 26510 22420 26516 22432
rect 26467 22392 26516 22420
rect 26467 22389 26479 22392
rect 26421 22383 26479 22389
rect 26510 22380 26516 22392
rect 26568 22380 26574 22432
rect 27356 22420 27384 22460
rect 27430 22448 27436 22500
rect 27488 22488 27494 22500
rect 27724 22488 27752 22519
rect 30834 22516 30840 22528
rect 30892 22516 30898 22568
rect 31128 22565 31156 22664
rect 31665 22661 31677 22695
rect 31711 22692 31723 22695
rect 31849 22695 31907 22701
rect 31849 22692 31861 22695
rect 31711 22664 31861 22692
rect 31711 22661 31723 22664
rect 31665 22655 31723 22661
rect 31849 22661 31861 22664
rect 31895 22692 31907 22695
rect 32214 22692 32220 22704
rect 31895 22664 32220 22692
rect 31895 22661 31907 22664
rect 31849 22655 31907 22661
rect 32214 22652 32220 22664
rect 32272 22692 32278 22704
rect 39960 22692 39988 22720
rect 32272 22664 37596 22692
rect 39330 22664 39988 22692
rect 47673 22695 47731 22701
rect 32272 22652 32278 22664
rect 31294 22584 31300 22636
rect 31352 22624 31358 22636
rect 31352 22596 32260 22624
rect 31352 22584 31358 22596
rect 31021 22559 31079 22565
rect 31021 22525 31033 22559
rect 31067 22525 31079 22559
rect 31021 22519 31079 22525
rect 31113 22559 31171 22565
rect 31113 22525 31125 22559
rect 31159 22525 31171 22559
rect 31113 22519 31171 22525
rect 27488 22460 27752 22488
rect 31036 22488 31064 22519
rect 31202 22516 31208 22568
rect 31260 22556 31266 22568
rect 32232 22556 32260 22596
rect 32306 22584 32312 22636
rect 32364 22624 32370 22636
rect 32401 22627 32459 22633
rect 32401 22624 32413 22627
rect 32364 22596 32413 22624
rect 32364 22584 32370 22596
rect 32401 22593 32413 22596
rect 32447 22593 32459 22627
rect 32401 22587 32459 22593
rect 33870 22584 33876 22636
rect 33928 22584 33934 22636
rect 34974 22584 34980 22636
rect 35032 22584 35038 22636
rect 37568 22633 37596 22664
rect 47673 22661 47685 22695
rect 47719 22692 47731 22695
rect 47719 22664 49096 22692
rect 47719 22661 47731 22664
rect 47673 22655 47731 22661
rect 49068 22636 49096 22664
rect 37553 22627 37611 22633
rect 37553 22593 37565 22627
rect 37599 22624 37611 22627
rect 37829 22627 37887 22633
rect 37829 22624 37841 22627
rect 37599 22596 37841 22624
rect 37599 22593 37611 22596
rect 37553 22587 37611 22593
rect 37829 22593 37841 22596
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 43901 22627 43959 22633
rect 43901 22593 43913 22627
rect 43947 22624 43959 22627
rect 44726 22624 44732 22636
rect 43947 22596 44732 22624
rect 43947 22593 43959 22596
rect 43901 22587 43959 22593
rect 44726 22584 44732 22596
rect 44784 22584 44790 22636
rect 48041 22627 48099 22633
rect 48041 22593 48053 22627
rect 48087 22624 48099 22627
rect 48314 22624 48320 22636
rect 48087 22596 48320 22624
rect 48087 22593 48099 22596
rect 48041 22587 48099 22593
rect 48314 22584 48320 22596
rect 48372 22584 48378 22636
rect 49050 22584 49056 22636
rect 49108 22584 49114 22636
rect 33045 22559 33103 22565
rect 33045 22556 33057 22559
rect 31260 22528 32168 22556
rect 32232 22528 33057 22556
rect 31260 22516 31266 22528
rect 31938 22488 31944 22500
rect 31036 22460 31944 22488
rect 27488 22448 27494 22460
rect 31938 22448 31944 22460
rect 31996 22448 32002 22500
rect 32140 22488 32168 22528
rect 33045 22525 33057 22528
rect 33091 22525 33103 22559
rect 33045 22519 33103 22525
rect 33594 22516 33600 22568
rect 33652 22516 33658 22568
rect 38105 22559 38163 22565
rect 38105 22525 38117 22559
rect 38151 22556 38163 22559
rect 44545 22559 44603 22565
rect 44545 22556 44557 22559
rect 38151 22528 44557 22556
rect 38151 22525 38163 22528
rect 38105 22519 38163 22525
rect 44545 22525 44557 22528
rect 44591 22525 44603 22559
rect 44545 22519 44603 22525
rect 32140 22460 33364 22488
rect 28810 22420 28816 22432
rect 27356 22392 28816 22420
rect 28810 22380 28816 22392
rect 28868 22380 28874 22432
rect 28994 22380 29000 22432
rect 29052 22420 29058 22432
rect 30101 22423 30159 22429
rect 30101 22420 30113 22423
rect 29052 22392 30113 22420
rect 29052 22380 29058 22392
rect 30101 22389 30113 22392
rect 30147 22389 30159 22423
rect 30101 22383 30159 22389
rect 32490 22380 32496 22432
rect 32548 22380 32554 22432
rect 33336 22420 33364 22460
rect 33410 22448 33416 22500
rect 33468 22488 33474 22500
rect 34701 22491 34759 22497
rect 34701 22488 34713 22491
rect 33468 22460 34713 22488
rect 33468 22448 33474 22460
rect 34701 22457 34713 22460
rect 34747 22457 34759 22491
rect 34701 22451 34759 22457
rect 47394 22448 47400 22500
rect 47452 22488 47458 22500
rect 49237 22491 49295 22497
rect 49237 22488 49249 22491
rect 47452 22460 49249 22488
rect 47452 22448 47458 22460
rect 49237 22457 49249 22460
rect 49283 22457 49295 22491
rect 49237 22451 49295 22457
rect 35345 22423 35403 22429
rect 35345 22420 35357 22423
rect 33336 22392 35357 22420
rect 35345 22389 35357 22392
rect 35391 22420 35403 22423
rect 35710 22420 35716 22432
rect 35391 22392 35716 22420
rect 35391 22389 35403 22392
rect 35345 22383 35403 22389
rect 35710 22380 35716 22392
rect 35768 22380 35774 22432
rect 37734 22380 37740 22432
rect 37792 22420 37798 22432
rect 39577 22423 39635 22429
rect 39577 22420 39589 22423
rect 37792 22392 39589 22420
rect 37792 22380 37798 22392
rect 39577 22389 39589 22392
rect 39623 22389 39635 22423
rect 39577 22383 39635 22389
rect 48498 22380 48504 22432
rect 48556 22380 48562 22432
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 2774 22176 2780 22228
rect 2832 22216 2838 22228
rect 2958 22216 2964 22228
rect 2832 22188 2964 22216
rect 2832 22176 2838 22188
rect 2958 22176 2964 22188
rect 3016 22176 3022 22228
rect 4798 22176 4804 22228
rect 4856 22216 4862 22228
rect 16114 22216 16120 22228
rect 4856 22188 16120 22216
rect 4856 22176 4862 22188
rect 16114 22176 16120 22188
rect 16172 22176 16178 22228
rect 16390 22176 16396 22228
rect 16448 22216 16454 22228
rect 16448 22188 18460 22216
rect 16448 22176 16454 22188
rect 2222 22108 2228 22160
rect 2280 22148 2286 22160
rect 3786 22148 3792 22160
rect 2280 22120 3792 22148
rect 2280 22108 2286 22120
rect 3786 22108 3792 22120
rect 3844 22108 3850 22160
rect 8757 22151 8815 22157
rect 8757 22117 8769 22151
rect 8803 22148 8815 22151
rect 9490 22148 9496 22160
rect 8803 22120 9496 22148
rect 8803 22117 8815 22120
rect 8757 22111 8815 22117
rect 9490 22108 9496 22120
rect 9548 22108 9554 22160
rect 11790 22108 11796 22160
rect 11848 22148 11854 22160
rect 11974 22148 11980 22160
rect 11848 22120 11980 22148
rect 11848 22108 11854 22120
rect 11974 22108 11980 22120
rect 12032 22148 12038 22160
rect 14734 22148 14740 22160
rect 12032 22120 14740 22148
rect 12032 22108 12038 22120
rect 14734 22108 14740 22120
rect 14792 22108 14798 22160
rect 18432 22148 18460 22188
rect 19886 22176 19892 22228
rect 19944 22216 19950 22228
rect 20070 22216 20076 22228
rect 19944 22188 20076 22216
rect 19944 22176 19950 22188
rect 20070 22176 20076 22188
rect 20128 22176 20134 22228
rect 23293 22219 23351 22225
rect 23293 22216 23305 22219
rect 23216 22188 23305 22216
rect 23216 22160 23244 22188
rect 23293 22185 23305 22188
rect 23339 22185 23351 22219
rect 23293 22179 23351 22185
rect 24578 22176 24584 22228
rect 24636 22176 24642 22228
rect 26040 22219 26098 22225
rect 26040 22216 26052 22219
rect 25884 22188 26052 22216
rect 22646 22148 22652 22160
rect 18432 22120 22652 22148
rect 22646 22108 22652 22120
rect 22704 22108 22710 22160
rect 23198 22108 23204 22160
rect 23256 22108 23262 22160
rect 25130 22148 25136 22160
rect 23952 22120 25136 22148
rect 1302 22040 1308 22092
rect 1360 22080 1366 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1360 22052 2053 22080
rect 1360 22040 1366 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 4614 22040 4620 22092
rect 4672 22040 4678 22092
rect 5813 22083 5871 22089
rect 5813 22049 5825 22083
rect 5859 22080 5871 22083
rect 5859 22052 6868 22080
rect 5859 22049 5871 22052
rect 5813 22043 5871 22049
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 22012 1823 22015
rect 1946 22012 1952 22024
rect 1811 21984 1952 22012
rect 1811 21981 1823 21984
rect 1765 21975 1823 21981
rect 1946 21972 1952 21984
rect 2004 21972 2010 22024
rect 3970 21972 3976 22024
rect 4028 21972 4034 22024
rect 6273 22015 6331 22021
rect 5736 21984 6224 22012
rect 3421 21947 3479 21953
rect 3421 21913 3433 21947
rect 3467 21944 3479 21947
rect 5736 21944 5764 21984
rect 3467 21916 5764 21944
rect 3467 21913 3479 21916
rect 3421 21907 3479 21913
rect 3602 21836 3608 21888
rect 3660 21836 3666 21888
rect 6086 21836 6092 21888
rect 6144 21836 6150 21888
rect 6196 21876 6224 21984
rect 6273 21981 6285 22015
rect 6319 22012 6331 22015
rect 6454 22012 6460 22024
rect 6319 21984 6460 22012
rect 6319 21981 6331 21984
rect 6273 21975 6331 21981
rect 6454 21972 6460 21984
rect 6512 21972 6518 22024
rect 6840 21944 6868 22052
rect 7374 22040 7380 22092
rect 7432 22080 7438 22092
rect 7650 22080 7656 22092
rect 7432 22052 7656 22080
rect 7432 22040 7438 22052
rect 7650 22040 7656 22052
rect 7708 22040 7714 22092
rect 7926 22040 7932 22092
rect 7984 22040 7990 22092
rect 8386 22040 8392 22092
rect 8444 22080 8450 22092
rect 8941 22083 8999 22089
rect 8941 22080 8953 22083
rect 8444 22052 8953 22080
rect 8444 22040 8450 22052
rect 8941 22049 8953 22052
rect 8987 22080 8999 22083
rect 9030 22080 9036 22092
rect 8987 22052 9036 22080
rect 8987 22049 8999 22052
rect 8941 22043 8999 22049
rect 9030 22040 9036 22052
rect 9088 22040 9094 22092
rect 9140 22052 9674 22080
rect 6914 21972 6920 22024
rect 6972 21972 6978 22024
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 9140 22012 9168 22052
rect 8619 21984 9168 22012
rect 9646 22012 9674 22052
rect 9858 22040 9864 22092
rect 9916 22040 9922 22092
rect 10778 22080 10784 22092
rect 10520 22052 10784 22080
rect 10520 22024 10548 22052
rect 10778 22040 10784 22052
rect 10836 22040 10842 22092
rect 11238 22040 11244 22092
rect 11296 22040 11302 22092
rect 13354 22040 13360 22092
rect 13412 22040 13418 22092
rect 15102 22040 15108 22092
rect 15160 22080 15166 22092
rect 15657 22083 15715 22089
rect 15657 22080 15669 22083
rect 15160 22052 15669 22080
rect 15160 22040 15166 22052
rect 15657 22049 15669 22052
rect 15703 22049 15715 22083
rect 15657 22043 15715 22049
rect 17129 22083 17187 22089
rect 17129 22049 17141 22083
rect 17175 22080 17187 22083
rect 19426 22080 19432 22092
rect 17175 22052 19432 22080
rect 17175 22049 17187 22052
rect 17129 22043 17187 22049
rect 19426 22040 19432 22052
rect 19484 22040 19490 22092
rect 20073 22083 20131 22089
rect 20073 22049 20085 22083
rect 20119 22080 20131 22083
rect 21910 22080 21916 22092
rect 20119 22052 21916 22080
rect 20119 22049 20131 22052
rect 20073 22043 20131 22049
rect 21910 22040 21916 22052
rect 21968 22040 21974 22092
rect 23952 22089 23980 22120
rect 25130 22108 25136 22120
rect 25188 22108 25194 22160
rect 23937 22083 23995 22089
rect 23937 22049 23949 22083
rect 23983 22080 23995 22083
rect 25225 22083 25283 22089
rect 23983 22052 24017 22080
rect 23983 22049 23995 22052
rect 23937 22043 23995 22049
rect 25225 22049 25237 22083
rect 25271 22080 25283 22083
rect 25884 22080 25912 22188
rect 26040 22185 26052 22188
rect 26086 22216 26098 22219
rect 27798 22216 27804 22228
rect 26086 22188 27804 22216
rect 26086 22185 26098 22188
rect 26040 22179 26098 22185
rect 27798 22176 27804 22188
rect 27856 22176 27862 22228
rect 28442 22176 28448 22228
rect 28500 22216 28506 22228
rect 28902 22216 28908 22228
rect 28500 22188 28908 22216
rect 28500 22176 28506 22188
rect 28902 22176 28908 22188
rect 28960 22216 28966 22228
rect 29549 22219 29607 22225
rect 29549 22216 29561 22219
rect 28960 22188 29561 22216
rect 28960 22176 28966 22188
rect 29549 22185 29561 22188
rect 29595 22216 29607 22219
rect 29733 22219 29791 22225
rect 29733 22216 29745 22219
rect 29595 22188 29745 22216
rect 29595 22185 29607 22188
rect 29549 22179 29607 22185
rect 29733 22185 29745 22188
rect 29779 22185 29791 22219
rect 29733 22179 29791 22185
rect 31662 22176 31668 22228
rect 31720 22216 31726 22228
rect 33226 22216 33232 22228
rect 31720 22188 33232 22216
rect 31720 22176 31726 22188
rect 33226 22176 33232 22188
rect 33284 22176 33290 22228
rect 27430 22108 27436 22160
rect 27488 22148 27494 22160
rect 27525 22151 27583 22157
rect 27525 22148 27537 22151
rect 27488 22120 27537 22148
rect 27488 22108 27494 22120
rect 27525 22117 27537 22120
rect 27571 22117 27583 22151
rect 27525 22111 27583 22117
rect 30668 22120 30880 22148
rect 25271 22052 25912 22080
rect 25271 22049 25283 22052
rect 25225 22043 25283 22049
rect 26786 22040 26792 22092
rect 26844 22080 26850 22092
rect 29181 22083 29239 22089
rect 26844 22052 28994 22080
rect 26844 22040 26850 22052
rect 9646 21984 10456 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 10428 21944 10456 21984
rect 10502 21972 10508 22024
rect 10560 21972 10566 22024
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 10612 21984 12541 22012
rect 10612 21944 10640 21984
rect 12529 21981 12541 21984
rect 12575 22012 12587 22015
rect 12802 22012 12808 22024
rect 12575 21984 12808 22012
rect 12575 21981 12587 21984
rect 12529 21975 12587 21981
rect 12802 21972 12808 21984
rect 12860 21972 12866 22024
rect 15194 21972 15200 22024
rect 15252 21972 15258 22024
rect 19518 21972 19524 22024
rect 19576 21972 19582 22024
rect 20346 21972 20352 22024
rect 20404 21972 20410 22024
rect 22002 21972 22008 22024
rect 22060 22012 22066 22024
rect 22370 22012 22376 22024
rect 22060 21984 22376 22012
rect 22060 21972 22066 21984
rect 22370 21972 22376 21984
rect 22428 21972 22434 22024
rect 23658 21972 23664 22024
rect 23716 21972 23722 22024
rect 23753 22015 23811 22021
rect 23753 21981 23765 22015
rect 23799 22012 23811 22015
rect 24762 22012 24768 22024
rect 23799 21984 24768 22012
rect 23799 21981 23811 21984
rect 23753 21975 23811 21981
rect 24762 21972 24768 21984
rect 24820 21972 24826 22024
rect 25682 21972 25688 22024
rect 25740 22012 25746 22024
rect 25777 22015 25835 22021
rect 25777 22012 25789 22015
rect 25740 21984 25789 22012
rect 25740 21972 25746 21984
rect 25777 21981 25789 21984
rect 25823 21981 25835 22015
rect 25777 21975 25835 21981
rect 28813 22015 28871 22021
rect 28813 21981 28825 22015
rect 28859 22012 28871 22015
rect 28966 22012 28994 22052
rect 29181 22049 29193 22083
rect 29227 22080 29239 22083
rect 29822 22080 29828 22092
rect 29227 22052 29828 22080
rect 29227 22049 29239 22052
rect 29181 22043 29239 22049
rect 29822 22040 29828 22052
rect 29880 22040 29886 22092
rect 30561 22083 30619 22089
rect 30561 22049 30573 22083
rect 30607 22080 30619 22083
rect 30668 22080 30696 22120
rect 30607 22052 30696 22080
rect 30607 22049 30619 22052
rect 30561 22043 30619 22049
rect 30742 22040 30748 22092
rect 30800 22040 30806 22092
rect 30852 22080 30880 22120
rect 31846 22108 31852 22160
rect 31904 22148 31910 22160
rect 32398 22148 32404 22160
rect 31904 22120 32404 22148
rect 31904 22108 31910 22120
rect 32398 22108 32404 22120
rect 32456 22148 32462 22160
rect 33873 22151 33931 22157
rect 33873 22148 33885 22151
rect 32456 22120 33885 22148
rect 32456 22108 32462 22120
rect 33873 22117 33885 22120
rect 33919 22117 33931 22151
rect 33873 22111 33931 22117
rect 30852 22052 32720 22080
rect 31849 22015 31907 22021
rect 31849 22012 31861 22015
rect 28859 21984 31861 22012
rect 28859 21981 28871 21984
rect 28813 21975 28871 21981
rect 31849 21981 31861 21984
rect 31895 21981 31907 22015
rect 32217 22015 32275 22021
rect 32217 22012 32229 22015
rect 31849 21975 31907 21981
rect 31956 21984 32229 22012
rect 14090 21944 14096 21956
rect 6840 21916 10364 21944
rect 10428 21916 10640 21944
rect 12406 21916 14096 21944
rect 8478 21876 8484 21888
rect 6196 21848 8484 21876
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 9674 21836 9680 21888
rect 9732 21836 9738 21888
rect 9766 21836 9772 21888
rect 9824 21836 9830 21888
rect 10336 21876 10364 21916
rect 12250 21876 12256 21888
rect 10336 21848 12256 21876
rect 12250 21836 12256 21848
rect 12308 21876 12314 21888
rect 12406 21876 12434 21916
rect 14090 21904 14096 21916
rect 14148 21904 14154 21956
rect 14366 21904 14372 21956
rect 14424 21904 14430 21956
rect 14918 21904 14924 21956
rect 14976 21904 14982 21956
rect 17405 21947 17463 21953
rect 17405 21913 17417 21947
rect 17451 21944 17463 21947
rect 17494 21944 17500 21956
rect 17451 21916 17500 21944
rect 17451 21913 17463 21916
rect 17405 21907 17463 21913
rect 17494 21904 17500 21916
rect 17552 21904 17558 21956
rect 18138 21904 18144 21956
rect 18196 21904 18202 21956
rect 18966 21904 18972 21956
rect 19024 21944 19030 21956
rect 19024 21916 20208 21944
rect 19024 21904 19030 21916
rect 12308 21848 12434 21876
rect 12308 21836 12314 21848
rect 12618 21836 12624 21888
rect 12676 21876 12682 21888
rect 14461 21879 14519 21885
rect 14461 21876 14473 21879
rect 12676 21848 14473 21876
rect 12676 21836 12682 21848
rect 14461 21845 14473 21848
rect 14507 21845 14519 21879
rect 14461 21839 14519 21845
rect 16758 21836 16764 21888
rect 16816 21876 16822 21888
rect 18877 21879 18935 21885
rect 18877 21876 18889 21879
rect 16816 21848 18889 21876
rect 16816 21836 16822 21848
rect 18877 21845 18889 21848
rect 18923 21845 18935 21879
rect 18877 21839 18935 21845
rect 19334 21836 19340 21888
rect 19392 21876 19398 21888
rect 19613 21879 19671 21885
rect 19613 21876 19625 21879
rect 19392 21848 19625 21876
rect 19392 21836 19398 21848
rect 19613 21845 19625 21848
rect 19659 21845 19671 21879
rect 20180 21876 20208 21916
rect 20254 21904 20260 21956
rect 20312 21944 20318 21956
rect 21269 21947 21327 21953
rect 21269 21944 21281 21947
rect 20312 21916 21281 21944
rect 20312 21904 20318 21916
rect 21269 21913 21281 21916
rect 21315 21913 21327 21947
rect 22649 21947 22707 21953
rect 21269 21907 21327 21913
rect 22020 21916 22600 21944
rect 22020 21876 22048 21916
rect 20180 21848 22048 21876
rect 22097 21879 22155 21885
rect 19613 21839 19671 21845
rect 22097 21845 22109 21879
rect 22143 21876 22155 21879
rect 22186 21876 22192 21888
rect 22143 21848 22192 21876
rect 22143 21845 22155 21848
rect 22097 21839 22155 21845
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 22370 21836 22376 21888
rect 22428 21836 22434 21888
rect 22572 21876 22600 21916
rect 22649 21913 22661 21947
rect 22695 21944 22707 21947
rect 24949 21947 25007 21953
rect 24949 21944 24961 21947
rect 22695 21916 24961 21944
rect 22695 21913 22707 21916
rect 22649 21907 22707 21913
rect 24949 21913 24961 21916
rect 24995 21913 25007 21947
rect 24949 21907 25007 21913
rect 25041 21947 25099 21953
rect 25041 21913 25053 21947
rect 25087 21944 25099 21947
rect 26326 21944 26332 21956
rect 25087 21916 26332 21944
rect 25087 21913 25099 21916
rect 25041 21907 25099 21913
rect 26326 21904 26332 21916
rect 26384 21904 26390 21956
rect 26510 21904 26516 21956
rect 26568 21904 26574 21956
rect 27338 21904 27344 21956
rect 27396 21944 27402 21956
rect 27396 21916 28764 21944
rect 27396 21904 27402 21916
rect 25866 21876 25872 21888
rect 22572 21848 25872 21876
rect 25866 21836 25872 21848
rect 25924 21836 25930 21888
rect 25958 21836 25964 21888
rect 26016 21876 26022 21888
rect 27985 21879 28043 21885
rect 27985 21876 27997 21879
rect 26016 21848 27997 21876
rect 26016 21836 26022 21848
rect 27985 21845 27997 21848
rect 28031 21845 28043 21879
rect 27985 21839 28043 21845
rect 28626 21836 28632 21888
rect 28684 21836 28690 21888
rect 28736 21876 28764 21916
rect 29270 21904 29276 21956
rect 29328 21904 29334 21956
rect 29380 21916 30604 21944
rect 29380 21876 29408 21916
rect 28736 21848 29408 21876
rect 30098 21836 30104 21888
rect 30156 21836 30162 21888
rect 30466 21836 30472 21888
rect 30524 21836 30530 21888
rect 30576 21876 30604 21916
rect 30742 21904 30748 21956
rect 30800 21944 30806 21956
rect 31389 21947 31447 21953
rect 31389 21944 31401 21947
rect 30800 21916 31401 21944
rect 30800 21904 30806 21916
rect 31389 21913 31401 21916
rect 31435 21944 31447 21947
rect 31956 21944 31984 21984
rect 32217 21981 32229 21984
rect 32263 21981 32275 22015
rect 32217 21975 32275 21981
rect 32398 21972 32404 22024
rect 32456 22012 32462 22024
rect 32585 22015 32643 22021
rect 32585 22012 32597 22015
rect 32456 21984 32597 22012
rect 32456 21972 32462 21984
rect 32585 21981 32597 21984
rect 32631 21981 32643 22015
rect 32585 21975 32643 21981
rect 31435 21916 31984 21944
rect 32692 21944 32720 22052
rect 32766 22040 32772 22092
rect 32824 22080 32830 22092
rect 34241 22083 34299 22089
rect 34241 22080 34253 22083
rect 32824 22052 34253 22080
rect 32824 22040 32830 22052
rect 34241 22049 34253 22052
rect 34287 22049 34299 22083
rect 34241 22043 34299 22049
rect 32858 21972 32864 22024
rect 32916 21972 32922 22024
rect 33318 21972 33324 22024
rect 33376 22012 33382 22024
rect 34057 22015 34115 22021
rect 34057 22012 34069 22015
rect 33376 21984 34069 22012
rect 33376 21972 33382 21984
rect 34057 21981 34069 21984
rect 34103 21981 34115 22015
rect 34057 21975 34115 21981
rect 48593 22015 48651 22021
rect 48593 21981 48605 22015
rect 48639 22012 48651 22015
rect 48682 22012 48688 22024
rect 48639 21984 48688 22012
rect 48639 21981 48651 21984
rect 48593 21975 48651 21981
rect 48682 21972 48688 21984
rect 48740 21972 48746 22024
rect 49050 21972 49056 22024
rect 49108 21972 49114 22024
rect 35802 21944 35808 21956
rect 32692 21916 35808 21944
rect 31435 21913 31447 21916
rect 31389 21907 31447 21913
rect 35802 21904 35808 21916
rect 35860 21904 35866 21956
rect 31481 21879 31539 21885
rect 31481 21876 31493 21879
rect 30576 21848 31493 21876
rect 31481 21845 31493 21848
rect 31527 21845 31539 21879
rect 31481 21839 31539 21845
rect 31662 21836 31668 21888
rect 31720 21876 31726 21888
rect 32125 21879 32183 21885
rect 32125 21876 32137 21879
rect 31720 21848 32137 21876
rect 31720 21836 31726 21848
rect 32125 21845 32137 21848
rect 32171 21845 32183 21879
rect 32125 21839 32183 21845
rect 32306 21836 32312 21888
rect 32364 21876 32370 21888
rect 33689 21879 33747 21885
rect 33689 21876 33701 21879
rect 32364 21848 33701 21876
rect 32364 21836 32370 21848
rect 33689 21845 33701 21848
rect 33735 21845 33747 21879
rect 33689 21839 33747 21845
rect 44726 21836 44732 21888
rect 44784 21876 44790 21888
rect 48409 21879 48467 21885
rect 48409 21876 48421 21879
rect 44784 21848 48421 21876
rect 44784 21836 44790 21848
rect 48409 21845 48421 21848
rect 48455 21845 48467 21879
rect 48409 21839 48467 21845
rect 49234 21836 49240 21888
rect 49292 21836 49298 21888
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 6457 21675 6515 21681
rect 6457 21641 6469 21675
rect 6503 21672 6515 21675
rect 9306 21672 9312 21684
rect 6503 21644 9312 21672
rect 6503 21641 6515 21644
rect 6457 21635 6515 21641
rect 9306 21632 9312 21644
rect 9364 21632 9370 21684
rect 9401 21675 9459 21681
rect 9401 21641 9413 21675
rect 9447 21641 9459 21675
rect 9401 21635 9459 21641
rect 1780 21576 4292 21604
rect 1780 21545 1808 21576
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21505 1823 21539
rect 1765 21499 1823 21505
rect 2498 21496 2504 21548
rect 2556 21536 2562 21548
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 2556 21508 3433 21536
rect 2556 21496 2562 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 4264 21536 4292 21576
rect 4338 21564 4344 21616
rect 4396 21564 4402 21616
rect 5718 21564 5724 21616
rect 5776 21604 5782 21616
rect 6730 21604 6736 21616
rect 5776 21576 6736 21604
rect 5776 21564 5782 21576
rect 6730 21564 6736 21576
rect 6788 21564 6794 21616
rect 7558 21564 7564 21616
rect 7616 21604 7622 21616
rect 7929 21607 7987 21613
rect 7929 21604 7941 21607
rect 7616 21576 7941 21604
rect 7616 21564 7622 21576
rect 7929 21573 7941 21576
rect 7975 21573 7987 21607
rect 7929 21567 7987 21573
rect 8018 21564 8024 21616
rect 8076 21604 8082 21616
rect 8386 21604 8392 21616
rect 8076 21576 8392 21604
rect 8076 21564 8082 21576
rect 8386 21564 8392 21576
rect 8444 21564 8450 21616
rect 9416 21604 9444 21635
rect 10962 21632 10968 21684
rect 11020 21632 11026 21684
rect 11149 21675 11207 21681
rect 11149 21641 11161 21675
rect 11195 21672 11207 21675
rect 11195 21644 15976 21672
rect 11195 21641 11207 21644
rect 11149 21635 11207 21641
rect 15948 21616 15976 21644
rect 16022 21632 16028 21684
rect 16080 21632 16086 21684
rect 19886 21672 19892 21684
rect 17512 21644 19892 21672
rect 9582 21604 9588 21616
rect 9416 21576 9588 21604
rect 9582 21564 9588 21576
rect 9640 21604 9646 21616
rect 15102 21604 15108 21616
rect 9640 21576 12388 21604
rect 14582 21576 15108 21604
rect 9640 21564 9646 21576
rect 5534 21536 5540 21548
rect 4264 21508 5540 21536
rect 3421 21499 3479 21505
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 5626 21496 5632 21548
rect 5684 21496 5690 21548
rect 7009 21539 7067 21545
rect 7009 21505 7021 21539
rect 7055 21536 7067 21539
rect 7374 21536 7380 21548
rect 7055 21508 7380 21536
rect 7055 21505 7067 21508
rect 7009 21499 7067 21505
rect 7374 21496 7380 21508
rect 7432 21496 7438 21548
rect 9490 21496 9496 21548
rect 9548 21536 9554 21548
rect 10229 21539 10287 21545
rect 10229 21536 10241 21539
rect 9548 21508 10241 21536
rect 9548 21496 9554 21508
rect 10229 21505 10241 21508
rect 10275 21505 10287 21539
rect 11606 21536 11612 21548
rect 10229 21499 10287 21505
rect 10428 21508 11612 21536
rect 2038 21428 2044 21480
rect 2096 21428 2102 21480
rect 5074 21428 5080 21480
rect 5132 21468 5138 21480
rect 5721 21471 5779 21477
rect 5721 21468 5733 21471
rect 5132 21440 5733 21468
rect 5132 21428 5138 21440
rect 5721 21437 5733 21440
rect 5767 21437 5779 21471
rect 5721 21431 5779 21437
rect 5905 21471 5963 21477
rect 5905 21437 5917 21471
rect 5951 21468 5963 21471
rect 6546 21468 6552 21480
rect 5951 21440 6552 21468
rect 5951 21437 5963 21440
rect 5905 21431 5963 21437
rect 6546 21428 6552 21440
rect 6604 21428 6610 21480
rect 7653 21471 7711 21477
rect 7653 21437 7665 21471
rect 7699 21468 7711 21471
rect 7699 21440 7788 21468
rect 7699 21437 7711 21440
rect 7653 21431 7711 21437
rect 4890 21360 4896 21412
rect 4948 21400 4954 21412
rect 7193 21403 7251 21409
rect 7193 21400 7205 21403
rect 4948 21372 7205 21400
rect 4948 21360 4954 21372
rect 7193 21369 7205 21372
rect 7239 21369 7251 21403
rect 7193 21363 7251 21369
rect 5166 21292 5172 21344
rect 5224 21332 5230 21344
rect 5261 21335 5319 21341
rect 5261 21332 5273 21335
rect 5224 21304 5273 21332
rect 5224 21292 5230 21304
rect 5261 21301 5273 21304
rect 5307 21301 5319 21335
rect 5261 21295 5319 21301
rect 6178 21292 6184 21344
rect 6236 21332 6242 21344
rect 6549 21335 6607 21341
rect 6549 21332 6561 21335
rect 6236 21304 6561 21332
rect 6236 21292 6242 21304
rect 6549 21301 6561 21304
rect 6595 21301 6607 21335
rect 7760 21332 7788 21440
rect 8478 21428 8484 21480
rect 8536 21468 8542 21480
rect 8536 21440 10272 21468
rect 8536 21428 8542 21440
rect 10244 21400 10272 21440
rect 10318 21428 10324 21480
rect 10376 21428 10382 21480
rect 10428 21400 10456 21508
rect 11606 21496 11612 21508
rect 11664 21536 11670 21548
rect 11974 21536 11980 21548
rect 11664 21508 11980 21536
rect 11664 21496 11670 21508
rect 11974 21496 11980 21508
rect 12032 21496 12038 21548
rect 12161 21539 12219 21545
rect 12161 21505 12173 21539
rect 12207 21505 12219 21539
rect 12161 21499 12219 21505
rect 10505 21471 10563 21477
rect 10505 21437 10517 21471
rect 10551 21437 10563 21471
rect 10505 21431 10563 21437
rect 10244 21372 10456 21400
rect 10520 21400 10548 21431
rect 10594 21428 10600 21480
rect 10652 21468 10658 21480
rect 12176 21468 12204 21499
rect 12250 21496 12256 21548
rect 12308 21496 12314 21548
rect 12360 21477 12388 21576
rect 15102 21564 15108 21576
rect 15160 21564 15166 21616
rect 15930 21564 15936 21616
rect 15988 21564 15994 21616
rect 12434 21496 12440 21548
rect 12492 21536 12498 21548
rect 13081 21539 13139 21545
rect 13081 21536 13093 21539
rect 12492 21508 13093 21536
rect 12492 21496 12498 21508
rect 13081 21505 13093 21508
rect 13127 21505 13139 21539
rect 13081 21499 13139 21505
rect 14642 21496 14648 21548
rect 14700 21536 14706 21548
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 14700 21508 16865 21536
rect 14700 21496 14706 21508
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 17512 21536 17540 21644
rect 19886 21632 19892 21644
rect 19944 21632 19950 21684
rect 20809 21675 20867 21681
rect 20809 21672 20821 21675
rect 20088 21644 20821 21672
rect 17586 21564 17592 21616
rect 17644 21604 17650 21616
rect 18966 21604 18972 21616
rect 17644 21576 18972 21604
rect 17644 21564 17650 21576
rect 18966 21564 18972 21576
rect 19024 21564 19030 21616
rect 16853 21499 16911 21505
rect 17236 21508 17540 21536
rect 20088 21522 20116 21644
rect 20809 21641 20821 21644
rect 20855 21672 20867 21675
rect 20993 21675 21051 21681
rect 20993 21672 21005 21675
rect 20855 21644 21005 21672
rect 20855 21641 20867 21644
rect 20809 21635 20867 21641
rect 20993 21641 21005 21644
rect 21039 21672 21051 21675
rect 21358 21672 21364 21684
rect 21039 21644 21364 21672
rect 21039 21641 21051 21644
rect 20993 21635 21051 21641
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 22830 21632 22836 21684
rect 22888 21672 22894 21684
rect 23017 21675 23075 21681
rect 23017 21672 23029 21675
rect 22888 21644 23029 21672
rect 22888 21632 22894 21644
rect 23017 21641 23029 21644
rect 23063 21641 23075 21675
rect 23017 21635 23075 21641
rect 22922 21604 22928 21616
rect 20272 21576 22928 21604
rect 10652 21440 12204 21468
rect 12345 21471 12403 21477
rect 10652 21428 10658 21440
rect 12345 21437 12357 21471
rect 12391 21437 12403 21471
rect 12345 21431 12403 21437
rect 13354 21428 13360 21480
rect 13412 21428 13418 21480
rect 14090 21428 14096 21480
rect 14148 21468 14154 21480
rect 16209 21471 16267 21477
rect 14148 21440 16160 21468
rect 14148 21428 14154 21440
rect 10520 21372 12434 21400
rect 8938 21332 8944 21344
rect 7760 21304 8944 21332
rect 6549 21295 6607 21301
rect 8938 21292 8944 21304
rect 8996 21292 9002 21344
rect 9582 21292 9588 21344
rect 9640 21332 9646 21344
rect 9677 21335 9735 21341
rect 9677 21332 9689 21335
rect 9640 21304 9689 21332
rect 9640 21292 9646 21304
rect 9677 21301 9689 21304
rect 9723 21301 9735 21335
rect 9677 21295 9735 21301
rect 9861 21335 9919 21341
rect 9861 21301 9873 21335
rect 9907 21332 9919 21335
rect 11054 21332 11060 21344
rect 9907 21304 11060 21332
rect 9907 21301 9919 21304
rect 9861 21295 9919 21301
rect 11054 21292 11060 21304
rect 11112 21292 11118 21344
rect 11333 21335 11391 21341
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11514 21332 11520 21344
rect 11379 21304 11520 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11514 21292 11520 21304
rect 11572 21292 11578 21344
rect 11790 21292 11796 21344
rect 11848 21292 11854 21344
rect 12406 21332 12434 21372
rect 15562 21360 15568 21412
rect 15620 21360 15626 21412
rect 16132 21400 16160 21440
rect 16209 21437 16221 21471
rect 16255 21468 16267 21471
rect 17236 21468 17264 21508
rect 16255 21440 17264 21468
rect 16255 21437 16267 21440
rect 16209 21431 16267 21437
rect 17310 21428 17316 21480
rect 17368 21428 17374 21480
rect 18693 21471 18751 21477
rect 18693 21437 18705 21471
rect 18739 21468 18751 21471
rect 18739 21440 18828 21468
rect 18739 21437 18751 21440
rect 18693 21431 18751 21437
rect 17218 21400 17224 21412
rect 16132 21372 17224 21400
rect 17218 21360 17224 21372
rect 17276 21360 17282 21412
rect 13538 21332 13544 21344
rect 12406 21304 13544 21332
rect 13538 21292 13544 21304
rect 13596 21292 13602 21344
rect 14734 21292 14740 21344
rect 14792 21332 14798 21344
rect 14829 21335 14887 21341
rect 14829 21332 14841 21335
rect 14792 21304 14841 21332
rect 14792 21292 14798 21304
rect 14829 21301 14841 21304
rect 14875 21301 14887 21335
rect 14829 21295 14887 21301
rect 14918 21292 14924 21344
rect 14976 21332 14982 21344
rect 15289 21335 15347 21341
rect 15289 21332 15301 21335
rect 14976 21304 15301 21332
rect 14976 21292 14982 21304
rect 15289 21301 15301 21304
rect 15335 21332 15347 21335
rect 18598 21332 18604 21344
rect 15335 21304 18604 21332
rect 15335 21301 15347 21304
rect 15289 21295 15347 21301
rect 18598 21292 18604 21304
rect 18656 21292 18662 21344
rect 18800 21332 18828 21440
rect 18966 21428 18972 21480
rect 19024 21428 19030 21480
rect 19058 21428 19064 21480
rect 19116 21468 19122 21480
rect 20272 21468 20300 21576
rect 22922 21564 22928 21576
rect 22980 21564 22986 21616
rect 21269 21539 21327 21545
rect 21269 21505 21281 21539
rect 21315 21536 21327 21539
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 21315 21508 22385 21536
rect 21315 21505 21327 21508
rect 21269 21499 21327 21505
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 23032 21536 23060 21635
rect 25038 21632 25044 21684
rect 25096 21672 25102 21684
rect 25096 21644 25176 21672
rect 25096 21632 25102 21644
rect 23661 21607 23719 21613
rect 23661 21573 23673 21607
rect 23707 21604 23719 21607
rect 23934 21604 23940 21616
rect 23707 21576 23940 21604
rect 23707 21573 23719 21576
rect 23661 21567 23719 21573
rect 23934 21564 23940 21576
rect 23992 21564 23998 21616
rect 24394 21564 24400 21616
rect 24452 21564 24458 21616
rect 23382 21536 23388 21548
rect 23032 21508 23388 21536
rect 22373 21499 22431 21505
rect 23382 21496 23388 21508
rect 23440 21496 23446 21548
rect 25148 21536 25176 21644
rect 25958 21632 25964 21684
rect 26016 21632 26022 21684
rect 26326 21632 26332 21684
rect 26384 21672 26390 21684
rect 27249 21675 27307 21681
rect 27249 21672 27261 21675
rect 26384 21644 27261 21672
rect 26384 21632 26390 21644
rect 27249 21641 27261 21644
rect 27295 21641 27307 21675
rect 27249 21635 27307 21641
rect 27709 21675 27767 21681
rect 27709 21641 27721 21675
rect 27755 21672 27767 21675
rect 31113 21675 31171 21681
rect 27755 21644 30052 21672
rect 27755 21641 27767 21644
rect 27709 21635 27767 21641
rect 26053 21607 26111 21613
rect 26053 21573 26065 21607
rect 26099 21604 26111 21607
rect 26099 21576 28304 21604
rect 26099 21573 26111 21576
rect 26053 21567 26111 21573
rect 25148 21508 26740 21536
rect 19116 21440 20300 21468
rect 22465 21471 22523 21477
rect 19116 21428 19122 21440
rect 22465 21437 22477 21471
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 24670 21468 24676 21480
rect 22695 21440 24676 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 20254 21360 20260 21412
rect 20312 21400 20318 21412
rect 22005 21403 22063 21409
rect 22005 21400 22017 21403
rect 20312 21372 22017 21400
rect 20312 21360 20318 21372
rect 22005 21369 22017 21372
rect 22051 21369 22063 21403
rect 22005 21363 22063 21369
rect 19426 21332 19432 21344
rect 18800 21304 19432 21332
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 19702 21292 19708 21344
rect 19760 21332 19766 21344
rect 20441 21335 20499 21341
rect 20441 21332 20453 21335
rect 19760 21304 20453 21332
rect 19760 21292 19766 21304
rect 20441 21301 20453 21304
rect 20487 21301 20499 21335
rect 22480 21332 22508 21431
rect 24670 21428 24676 21440
rect 24728 21468 24734 21480
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24728 21440 25145 21468
rect 24728 21428 24734 21440
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 26237 21471 26295 21477
rect 26237 21437 26249 21471
rect 26283 21468 26295 21471
rect 26602 21468 26608 21480
rect 26283 21440 26608 21468
rect 26283 21437 26295 21440
rect 26237 21431 26295 21437
rect 26602 21428 26608 21440
rect 26660 21428 26666 21480
rect 26712 21477 26740 21508
rect 26878 21496 26884 21548
rect 26936 21536 26942 21548
rect 27338 21536 27344 21548
rect 26936 21508 27344 21536
rect 26936 21496 26942 21508
rect 27338 21496 27344 21508
rect 27396 21496 27402 21548
rect 27617 21539 27675 21545
rect 27617 21536 27629 21539
rect 27540 21508 27629 21536
rect 26697 21471 26755 21477
rect 26697 21437 26709 21471
rect 26743 21468 26755 21471
rect 27540 21468 27568 21508
rect 27617 21505 27629 21508
rect 27663 21536 27675 21539
rect 27890 21536 27896 21548
rect 27663 21508 27896 21536
rect 27663 21505 27675 21508
rect 27617 21499 27675 21505
rect 27890 21496 27896 21508
rect 27948 21496 27954 21548
rect 27801 21471 27859 21477
rect 27801 21468 27813 21471
rect 26743 21440 27568 21468
rect 27632 21440 27813 21468
rect 26743 21437 26755 21440
rect 26697 21431 26755 21437
rect 27632 21412 27660 21440
rect 27801 21437 27813 21440
rect 27847 21437 27859 21471
rect 27801 21431 27859 21437
rect 24762 21360 24768 21412
rect 24820 21400 24826 21412
rect 25593 21403 25651 21409
rect 25593 21400 25605 21403
rect 24820 21372 25605 21400
rect 24820 21360 24826 21372
rect 25593 21369 25605 21372
rect 25639 21369 25651 21403
rect 25593 21363 25651 21369
rect 27614 21360 27620 21412
rect 27672 21360 27678 21412
rect 28276 21400 28304 21576
rect 28718 21564 28724 21616
rect 28776 21604 28782 21616
rect 28994 21604 29000 21616
rect 28776 21576 29000 21604
rect 28776 21564 28782 21576
rect 28994 21564 29000 21576
rect 29052 21564 29058 21616
rect 30024 21604 30052 21644
rect 31113 21641 31125 21675
rect 31159 21672 31171 21675
rect 31159 21644 33180 21672
rect 31159 21641 31171 21644
rect 31113 21635 31171 21641
rect 33152 21604 33180 21644
rect 33226 21632 33232 21684
rect 33284 21632 33290 21684
rect 34514 21604 34520 21616
rect 30024 21576 33088 21604
rect 33152 21576 34520 21604
rect 29822 21496 29828 21548
rect 29880 21496 29886 21548
rect 31021 21539 31079 21545
rect 31021 21536 31033 21539
rect 30300 21508 31033 21536
rect 28442 21428 28448 21480
rect 28500 21428 28506 21480
rect 28718 21428 28724 21480
rect 28776 21428 28782 21480
rect 28810 21428 28816 21480
rect 28868 21468 28874 21480
rect 30300 21468 30328 21508
rect 31021 21505 31033 21508
rect 31067 21536 31079 21539
rect 31067 21508 31340 21536
rect 31067 21505 31079 21508
rect 31021 21499 31079 21505
rect 28868 21440 30328 21468
rect 31205 21471 31263 21477
rect 28868 21428 28874 21440
rect 31205 21437 31217 21471
rect 31251 21437 31263 21471
rect 31205 21431 31263 21437
rect 31220 21400 31248 21431
rect 28276 21372 28488 21400
rect 25314 21332 25320 21344
rect 22480 21304 25320 21332
rect 20441 21295 20499 21301
rect 25314 21292 25320 21304
rect 25372 21292 25378 21344
rect 28460 21332 28488 21372
rect 30208 21372 31248 21400
rect 30208 21344 30236 21372
rect 30098 21332 30104 21344
rect 28460 21304 30104 21332
rect 30098 21292 30104 21304
rect 30156 21292 30162 21344
rect 30190 21292 30196 21344
rect 30248 21292 30254 21344
rect 30650 21292 30656 21344
rect 30708 21292 30714 21344
rect 31312 21332 31340 21508
rect 31478 21496 31484 21548
rect 31536 21536 31542 21548
rect 31665 21539 31723 21545
rect 31665 21536 31677 21539
rect 31536 21508 31677 21536
rect 31536 21496 31542 21508
rect 31665 21505 31677 21508
rect 31711 21505 31723 21539
rect 31665 21499 31723 21505
rect 32214 21496 32220 21548
rect 32272 21536 32278 21548
rect 32401 21539 32459 21545
rect 32401 21536 32413 21539
rect 32272 21508 32413 21536
rect 32272 21496 32278 21508
rect 32401 21505 32413 21508
rect 32447 21536 32459 21539
rect 32861 21539 32919 21545
rect 32861 21536 32873 21539
rect 32447 21508 32873 21536
rect 32447 21505 32459 21508
rect 32401 21499 32459 21505
rect 32861 21505 32873 21508
rect 32907 21505 32919 21539
rect 33060 21536 33088 21576
rect 34514 21564 34520 21576
rect 34572 21564 34578 21616
rect 35526 21536 35532 21548
rect 33060 21508 35532 21536
rect 32861 21499 32919 21505
rect 35526 21496 35532 21508
rect 35584 21496 35590 21548
rect 47854 21496 47860 21548
rect 47912 21536 47918 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 47912 21508 47961 21536
rect 47912 21496 47918 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 31570 21428 31576 21480
rect 31628 21468 31634 21480
rect 33597 21471 33655 21477
rect 33597 21468 33609 21471
rect 31628 21440 33609 21468
rect 31628 21428 31634 21440
rect 33597 21437 33609 21440
rect 33643 21437 33655 21471
rect 33597 21431 33655 21437
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 31386 21360 31392 21412
rect 31444 21400 31450 21412
rect 32398 21400 32404 21412
rect 31444 21372 32404 21400
rect 31444 21360 31450 21372
rect 32398 21360 32404 21372
rect 32456 21400 32462 21412
rect 33045 21403 33103 21409
rect 33045 21400 33057 21403
rect 32456 21372 33057 21400
rect 32456 21360 32462 21372
rect 33045 21369 33057 21372
rect 33091 21369 33103 21403
rect 33045 21363 33103 21369
rect 31754 21332 31760 21344
rect 31312 21304 31760 21332
rect 31754 21292 31760 21304
rect 31812 21332 31818 21344
rect 31849 21335 31907 21341
rect 31849 21332 31861 21335
rect 31812 21304 31861 21332
rect 31812 21292 31818 21304
rect 31849 21301 31861 21304
rect 31895 21301 31907 21335
rect 31849 21295 31907 21301
rect 32490 21292 32496 21344
rect 32548 21292 32554 21344
rect 33410 21292 33416 21344
rect 33468 21292 33474 21344
rect 47673 21335 47731 21341
rect 47673 21301 47685 21335
rect 47719 21332 47731 21335
rect 47854 21332 47860 21344
rect 47719 21304 47860 21332
rect 47719 21301 47731 21304
rect 47673 21295 47731 21301
rect 47854 21292 47860 21304
rect 47912 21292 47918 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 3421 21131 3479 21137
rect 3421 21097 3433 21131
rect 3467 21128 3479 21131
rect 7098 21128 7104 21140
rect 3467 21100 7104 21128
rect 3467 21097 3479 21100
rect 3421 21091 3479 21097
rect 7098 21088 7104 21100
rect 7156 21088 7162 21140
rect 10318 21128 10324 21140
rect 7208 21100 10324 21128
rect 3326 21020 3332 21072
rect 3384 21060 3390 21072
rect 5077 21063 5135 21069
rect 5077 21060 5089 21063
rect 3384 21032 5089 21060
rect 3384 21020 3390 21032
rect 5077 21029 5089 21032
rect 5123 21029 5135 21063
rect 5077 21023 5135 21029
rect 6730 21020 6736 21072
rect 6788 21060 6794 21072
rect 7208 21060 7236 21100
rect 10318 21088 10324 21100
rect 10376 21088 10382 21140
rect 10965 21131 11023 21137
rect 10965 21097 10977 21131
rect 11011 21128 11023 21131
rect 15194 21128 15200 21140
rect 11011 21100 15200 21128
rect 11011 21097 11023 21100
rect 10965 21091 11023 21097
rect 15194 21088 15200 21100
rect 15252 21088 15258 21140
rect 23566 21128 23572 21140
rect 16224 21100 23572 21128
rect 6788 21032 7236 21060
rect 6788 21020 6794 21032
rect 7650 21020 7656 21072
rect 7708 21060 7714 21072
rect 7837 21063 7895 21069
rect 7837 21060 7849 21063
rect 7708 21032 7849 21060
rect 7708 21020 7714 21032
rect 7837 21029 7849 21032
rect 7883 21029 7895 21063
rect 11790 21060 11796 21072
rect 7837 21023 7895 21029
rect 8312 21032 11796 21060
rect 2130 20952 2136 21004
rect 2188 20992 2194 21004
rect 4154 20992 4160 21004
rect 2188 20964 4160 20992
rect 2188 20952 2194 20964
rect 4154 20952 4160 20964
rect 4212 20952 4218 21004
rect 4246 20952 4252 21004
rect 4304 20952 4310 21004
rect 5721 20995 5779 21001
rect 5721 20961 5733 20995
rect 5767 20992 5779 20995
rect 7006 20992 7012 21004
rect 5767 20964 7012 20992
rect 5767 20961 5779 20964
rect 5721 20955 5779 20961
rect 7006 20952 7012 20964
rect 7064 20992 7070 21004
rect 7374 20992 7380 21004
rect 7064 20964 7380 20992
rect 7064 20952 7070 20964
rect 7374 20952 7380 20964
rect 7432 20952 7438 21004
rect 8312 21001 8340 21032
rect 11790 21020 11796 21032
rect 11848 21020 11854 21072
rect 14642 21060 14648 21072
rect 12406 21032 14648 21060
rect 8297 20995 8355 21001
rect 8297 20961 8309 20995
rect 8343 20961 8355 20995
rect 8297 20955 8355 20961
rect 8481 20995 8539 21001
rect 8481 20961 8493 20995
rect 8527 20992 8539 20995
rect 8846 20992 8852 21004
rect 8527 20964 8852 20992
rect 8527 20961 8539 20964
rect 8481 20955 8539 20961
rect 8846 20952 8852 20964
rect 8904 20952 8910 21004
rect 9585 20995 9643 21001
rect 9585 20992 9597 20995
rect 8956 20964 9597 20992
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 1854 20924 1860 20936
rect 1811 20896 1860 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 3970 20884 3976 20936
rect 4028 20884 4034 20936
rect 5442 20884 5448 20936
rect 5500 20884 5506 20936
rect 7745 20927 7803 20933
rect 7745 20893 7757 20927
rect 7791 20924 7803 20927
rect 8202 20924 8208 20936
rect 7791 20896 8208 20924
rect 7791 20893 7803 20896
rect 7745 20887 7803 20893
rect 8202 20884 8208 20896
rect 8260 20884 8266 20936
rect 8570 20884 8576 20936
rect 8628 20924 8634 20936
rect 8956 20924 8984 20964
rect 9585 20961 9597 20964
rect 9631 20961 9643 20995
rect 9585 20955 9643 20961
rect 11514 20952 11520 21004
rect 11572 20992 11578 21004
rect 12406 20992 12434 21032
rect 14642 21020 14648 21032
rect 14700 21020 14706 21072
rect 11572 20964 12434 20992
rect 11572 20952 11578 20964
rect 12526 20952 12532 21004
rect 12584 20952 12590 21004
rect 14277 20995 14335 21001
rect 14277 20961 14289 20995
rect 14323 20992 14335 20995
rect 14918 20992 14924 21004
rect 14323 20964 14924 20992
rect 14323 20961 14335 20964
rect 14277 20955 14335 20961
rect 14918 20952 14924 20964
rect 14976 20952 14982 21004
rect 15105 20995 15163 21001
rect 15105 20961 15117 20995
rect 15151 20992 15163 20995
rect 15470 20992 15476 21004
rect 15151 20964 15476 20992
rect 15151 20961 15163 20964
rect 15105 20955 15163 20961
rect 15470 20952 15476 20964
rect 15528 20952 15534 21004
rect 16224 21001 16252 21100
rect 23566 21088 23572 21100
rect 23624 21088 23630 21140
rect 23658 21088 23664 21140
rect 23716 21128 23722 21140
rect 27706 21128 27712 21140
rect 23716 21100 24900 21128
rect 23716 21088 23722 21100
rect 17604 21032 18920 21060
rect 16209 20995 16267 21001
rect 16209 20961 16221 20995
rect 16255 20961 16267 20995
rect 16209 20955 16267 20961
rect 16390 20952 16396 21004
rect 16448 20952 16454 21004
rect 17604 21001 17632 21032
rect 17589 20995 17647 21001
rect 17589 20961 17601 20995
rect 17635 20961 17647 20995
rect 17589 20955 17647 20961
rect 18785 20995 18843 21001
rect 18785 20961 18797 20995
rect 18831 20961 18843 20995
rect 18892 20992 18920 21032
rect 21358 21020 21364 21072
rect 21416 21060 21422 21072
rect 22097 21063 22155 21069
rect 22097 21060 22109 21063
rect 21416 21032 22109 21060
rect 21416 21020 21422 21032
rect 22097 21029 22109 21032
rect 22143 21029 22155 21063
rect 22097 21023 22155 21029
rect 22370 21020 22376 21072
rect 22428 21060 22434 21072
rect 22428 21032 23796 21060
rect 22428 21020 22434 21032
rect 19702 20992 19708 21004
rect 18892 20964 19708 20992
rect 18785 20955 18843 20961
rect 8628 20896 8984 20924
rect 8628 20884 8634 20896
rect 9030 20884 9036 20936
rect 9088 20924 9094 20936
rect 9125 20927 9183 20933
rect 9125 20924 9137 20927
rect 9088 20896 9137 20924
rect 9088 20884 9094 20896
rect 9125 20893 9137 20896
rect 9171 20893 9183 20927
rect 9125 20887 9183 20893
rect 11698 20884 11704 20936
rect 11756 20924 11762 20936
rect 11977 20927 12035 20933
rect 11977 20924 11989 20927
rect 11756 20896 11989 20924
rect 11756 20884 11762 20896
rect 11977 20893 11989 20896
rect 12023 20924 12035 20927
rect 12066 20924 12072 20936
rect 12023 20896 12072 20924
rect 12023 20893 12035 20896
rect 11977 20887 12035 20893
rect 12066 20884 12072 20896
rect 12124 20884 12130 20936
rect 16574 20924 16580 20936
rect 14936 20896 16580 20924
rect 2774 20816 2780 20868
rect 2832 20816 2838 20868
rect 3510 20816 3516 20868
rect 3568 20856 3574 20868
rect 3605 20859 3663 20865
rect 3605 20856 3617 20859
rect 3568 20828 3617 20856
rect 3568 20816 3574 20828
rect 3605 20825 3617 20828
rect 3651 20856 3663 20859
rect 5626 20856 5632 20868
rect 3651 20828 5632 20856
rect 3651 20825 3663 20828
rect 3605 20819 3663 20825
rect 5626 20816 5632 20828
rect 5684 20816 5690 20868
rect 6178 20856 6184 20868
rect 5828 20828 6184 20856
rect 5258 20748 5264 20800
rect 5316 20788 5322 20800
rect 5828 20788 5856 20828
rect 6178 20816 6184 20828
rect 6236 20816 6242 20868
rect 7098 20816 7104 20868
rect 7156 20856 7162 20868
rect 10594 20856 10600 20868
rect 7156 20828 10600 20856
rect 7156 20816 7162 20828
rect 10594 20816 10600 20828
rect 10652 20816 10658 20868
rect 11330 20816 11336 20868
rect 11388 20816 11394 20868
rect 13725 20859 13783 20865
rect 13725 20825 13737 20859
rect 13771 20856 13783 20859
rect 14090 20856 14096 20868
rect 13771 20828 14096 20856
rect 13771 20825 13783 20828
rect 13725 20819 13783 20825
rect 14090 20816 14096 20828
rect 14148 20816 14154 20868
rect 14936 20856 14964 20896
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 17402 20884 17408 20936
rect 17460 20884 17466 20936
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20924 18567 20927
rect 18598 20924 18604 20936
rect 18555 20896 18604 20924
rect 18555 20893 18567 20896
rect 18509 20887 18567 20893
rect 18598 20884 18604 20896
rect 18656 20884 18662 20936
rect 18800 20924 18828 20955
rect 19702 20952 19708 20964
rect 19760 20952 19766 21004
rect 21450 20952 21456 21004
rect 21508 20992 21514 21004
rect 21545 20995 21603 21001
rect 21545 20992 21557 20995
rect 21508 20964 21557 20992
rect 21508 20952 21514 20964
rect 21545 20961 21557 20964
rect 21591 20961 21603 20995
rect 21545 20955 21603 20961
rect 22741 20995 22799 21001
rect 22741 20961 22753 20995
rect 22787 20992 22799 20995
rect 23566 20992 23572 21004
rect 22787 20964 23572 20992
rect 22787 20961 22799 20964
rect 22741 20955 22799 20961
rect 23566 20952 23572 20964
rect 23624 20952 23630 21004
rect 23768 21001 23796 21032
rect 23753 20995 23811 21001
rect 23753 20961 23765 20995
rect 23799 20961 23811 20995
rect 23753 20955 23811 20961
rect 23842 20952 23848 21004
rect 23900 20952 23906 21004
rect 18874 20924 18880 20936
rect 18800 20896 18880 20924
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 19426 20884 19432 20936
rect 19484 20884 19490 20936
rect 21468 20924 21496 20952
rect 20838 20896 21496 20924
rect 21821 20927 21879 20933
rect 21821 20893 21833 20927
rect 21867 20924 21879 20927
rect 22278 20924 22284 20936
rect 21867 20896 22284 20924
rect 21867 20893 21879 20896
rect 21821 20887 21879 20893
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 24118 20884 24124 20936
rect 24176 20924 24182 20936
rect 24762 20924 24768 20936
rect 24176 20896 24768 20924
rect 24176 20884 24182 20896
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 24872 20924 24900 21100
rect 25240 21100 27712 21128
rect 25240 21001 25268 21100
rect 27706 21088 27712 21100
rect 27764 21088 27770 21140
rect 27798 21088 27804 21140
rect 27856 21088 27862 21140
rect 27890 21088 27896 21140
rect 27948 21128 27954 21140
rect 28902 21128 28908 21140
rect 27948 21100 28908 21128
rect 27948 21088 27954 21100
rect 28902 21088 28908 21100
rect 28960 21088 28966 21140
rect 30006 21088 30012 21140
rect 30064 21088 30070 21140
rect 30098 21088 30104 21140
rect 30156 21128 30162 21140
rect 31386 21128 31392 21140
rect 30156 21100 31392 21128
rect 30156 21088 30162 21100
rect 31386 21088 31392 21100
rect 31444 21088 31450 21140
rect 32493 21131 32551 21137
rect 32493 21097 32505 21131
rect 32539 21128 32551 21131
rect 32582 21128 32588 21140
rect 32539 21100 32588 21128
rect 32539 21097 32551 21100
rect 32493 21091 32551 21097
rect 32582 21088 32588 21100
rect 32640 21088 32646 21140
rect 44818 21088 44824 21140
rect 44876 21128 44882 21140
rect 47486 21128 47492 21140
rect 44876 21100 47492 21128
rect 44876 21088 44882 21100
rect 47486 21088 47492 21100
rect 47544 21088 47550 21140
rect 49050 21088 49056 21140
rect 49108 21128 49114 21140
rect 49421 21131 49479 21137
rect 49421 21128 49433 21131
rect 49108 21100 49433 21128
rect 49108 21088 49114 21100
rect 49421 21097 49433 21100
rect 49467 21097 49479 21131
rect 49421 21091 49479 21097
rect 28258 21020 28264 21072
rect 28316 21060 28322 21072
rect 30024 21060 30052 21088
rect 33410 21060 33416 21072
rect 28316 21032 28580 21060
rect 30024 21032 33416 21060
rect 28316 21020 28322 21032
rect 25225 20995 25283 21001
rect 25225 20961 25237 20995
rect 25271 20961 25283 20995
rect 25225 20955 25283 20961
rect 25682 20952 25688 21004
rect 25740 20992 25746 21004
rect 26050 20992 26056 21004
rect 25740 20964 26056 20992
rect 25740 20952 25746 20964
rect 26050 20952 26056 20964
rect 26108 20952 26114 21004
rect 26329 20995 26387 21001
rect 26329 20961 26341 20995
rect 26375 20992 26387 20995
rect 27614 20992 27620 21004
rect 26375 20964 27620 20992
rect 26375 20961 26387 20964
rect 26329 20955 26387 20961
rect 27614 20952 27620 20964
rect 27672 20952 27678 21004
rect 28552 21001 28580 21032
rect 33410 21020 33416 21032
rect 33468 21020 33474 21072
rect 28537 20995 28595 21001
rect 28537 20961 28549 20995
rect 28583 20961 28595 20995
rect 28537 20955 28595 20961
rect 29086 20952 29092 21004
rect 29144 20992 29150 21004
rect 30009 20995 30067 21001
rect 30009 20992 30021 20995
rect 29144 20964 30021 20992
rect 29144 20952 29150 20964
rect 30009 20961 30021 20964
rect 30055 20961 30067 20995
rect 30009 20955 30067 20961
rect 30466 20952 30472 21004
rect 30524 20992 30530 21004
rect 31662 20992 31668 21004
rect 30524 20964 31668 20992
rect 30524 20952 30530 20964
rect 31662 20952 31668 20964
rect 31720 20992 31726 21004
rect 36446 20992 36452 21004
rect 31720 20964 36452 20992
rect 31720 20952 31726 20964
rect 36446 20952 36452 20964
rect 36504 20952 36510 21004
rect 25866 20924 25872 20936
rect 24872 20896 25872 20924
rect 25866 20884 25872 20896
rect 25924 20884 25930 20936
rect 28261 20927 28319 20933
rect 28261 20893 28273 20927
rect 28307 20924 28319 20927
rect 28442 20924 28448 20936
rect 28307 20896 28448 20924
rect 28307 20893 28319 20896
rect 28261 20887 28319 20893
rect 28442 20884 28448 20896
rect 28500 20924 28506 20936
rect 29270 20924 29276 20936
rect 28500 20896 29276 20924
rect 28500 20884 28506 20896
rect 29270 20884 29276 20896
rect 29328 20884 29334 20936
rect 29546 20884 29552 20936
rect 29604 20924 29610 20936
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 29604 20896 29745 20924
rect 29604 20884 29610 20896
rect 29733 20893 29745 20896
rect 29779 20893 29791 20927
rect 29733 20887 29791 20893
rect 31110 20884 31116 20936
rect 31168 20884 31174 20936
rect 32674 20884 32680 20936
rect 32732 20924 32738 20936
rect 32953 20927 33011 20933
rect 32953 20924 32965 20927
rect 32732 20896 32965 20924
rect 32732 20884 32738 20896
rect 32953 20893 32965 20896
rect 32999 20893 33011 20927
rect 32953 20887 33011 20893
rect 14568 20828 14964 20856
rect 15013 20859 15071 20865
rect 5316 20760 5856 20788
rect 5316 20748 5322 20760
rect 5902 20748 5908 20800
rect 5960 20788 5966 20800
rect 7193 20791 7251 20797
rect 7193 20788 7205 20791
rect 5960 20760 7205 20788
rect 5960 20748 5966 20760
rect 7193 20757 7205 20760
rect 7239 20757 7251 20791
rect 7193 20751 7251 20757
rect 7561 20791 7619 20797
rect 7561 20757 7573 20791
rect 7607 20788 7619 20791
rect 9214 20788 9220 20800
rect 7607 20760 9220 20788
rect 7607 20757 7619 20760
rect 7561 20751 7619 20757
rect 9214 20748 9220 20760
rect 9272 20748 9278 20800
rect 11422 20748 11428 20800
rect 11480 20748 11486 20800
rect 13906 20748 13912 20800
rect 13964 20748 13970 20800
rect 14568 20797 14596 20828
rect 15013 20825 15025 20859
rect 15059 20856 15071 20859
rect 25041 20859 25099 20865
rect 15059 20828 18736 20856
rect 15059 20825 15071 20828
rect 15013 20819 15071 20825
rect 14553 20791 14611 20797
rect 14553 20757 14565 20791
rect 14599 20757 14611 20791
rect 14553 20751 14611 20757
rect 14918 20748 14924 20800
rect 14976 20748 14982 20800
rect 15746 20748 15752 20800
rect 15804 20748 15810 20800
rect 16117 20791 16175 20797
rect 16117 20757 16129 20791
rect 16163 20788 16175 20791
rect 16666 20788 16672 20800
rect 16163 20760 16672 20788
rect 16163 20757 16175 20760
rect 16117 20751 16175 20757
rect 16666 20748 16672 20760
rect 16724 20748 16730 20800
rect 16942 20748 16948 20800
rect 17000 20748 17006 20800
rect 17034 20748 17040 20800
rect 17092 20788 17098 20800
rect 17313 20791 17371 20797
rect 17313 20788 17325 20791
rect 17092 20760 17325 20788
rect 17092 20748 17098 20760
rect 17313 20757 17325 20760
rect 17359 20788 17371 20791
rect 17586 20788 17592 20800
rect 17359 20760 17592 20788
rect 17359 20757 17371 20760
rect 17313 20751 17371 20757
rect 17586 20748 17592 20760
rect 17644 20748 17650 20800
rect 17678 20748 17684 20800
rect 17736 20788 17742 20800
rect 18141 20791 18199 20797
rect 18141 20788 18153 20791
rect 17736 20760 18153 20788
rect 17736 20748 17742 20760
rect 18141 20757 18153 20760
rect 18187 20757 18199 20791
rect 18141 20751 18199 20757
rect 18414 20748 18420 20800
rect 18472 20788 18478 20800
rect 18601 20791 18659 20797
rect 18601 20788 18613 20791
rect 18472 20760 18613 20788
rect 18472 20748 18478 20760
rect 18601 20757 18613 20760
rect 18647 20757 18659 20791
rect 18708 20788 18736 20828
rect 25041 20825 25053 20859
rect 25087 20856 25099 20859
rect 26234 20856 26240 20868
rect 25087 20828 26240 20856
rect 25087 20825 25099 20828
rect 25041 20819 25099 20825
rect 26234 20816 26240 20828
rect 26292 20816 26298 20868
rect 26602 20816 26608 20868
rect 26660 20856 26666 20868
rect 26660 20828 26818 20856
rect 26660 20816 26666 20828
rect 31846 20816 31852 20868
rect 31904 20816 31910 20868
rect 21082 20788 21088 20800
rect 18708 20760 21088 20788
rect 18601 20751 18659 20757
rect 21082 20748 21088 20760
rect 21140 20748 21146 20800
rect 21174 20748 21180 20800
rect 21232 20748 21238 20800
rect 22462 20748 22468 20800
rect 22520 20748 22526 20800
rect 22554 20748 22560 20800
rect 22612 20748 22618 20800
rect 22646 20748 22652 20800
rect 22704 20788 22710 20800
rect 23293 20791 23351 20797
rect 23293 20788 23305 20791
rect 22704 20760 23305 20788
rect 22704 20748 22710 20760
rect 23293 20757 23305 20760
rect 23339 20757 23351 20791
rect 23293 20751 23351 20757
rect 23658 20748 23664 20800
rect 23716 20748 23722 20800
rect 23934 20748 23940 20800
rect 23992 20788 23998 20800
rect 24673 20791 24731 20797
rect 24673 20788 24685 20791
rect 23992 20760 24685 20788
rect 23992 20748 23998 20760
rect 24673 20757 24685 20760
rect 24719 20757 24731 20791
rect 24673 20751 24731 20757
rect 25133 20791 25191 20797
rect 25133 20757 25145 20791
rect 25179 20788 25191 20791
rect 30650 20788 30656 20800
rect 25179 20760 30656 20788
rect 25179 20757 25191 20760
rect 25133 20751 25191 20757
rect 30650 20748 30656 20760
rect 30708 20748 30714 20800
rect 31202 20748 31208 20800
rect 31260 20748 31266 20800
rect 31938 20748 31944 20800
rect 31996 20748 32002 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 5629 20587 5687 20593
rect 5629 20553 5641 20587
rect 5675 20584 5687 20587
rect 7006 20584 7012 20596
rect 5675 20556 7012 20584
rect 5675 20553 5687 20556
rect 5629 20547 5687 20553
rect 7006 20544 7012 20556
rect 7064 20544 7070 20596
rect 8386 20544 8392 20596
rect 8444 20584 8450 20596
rect 9490 20584 9496 20596
rect 8444 20556 9496 20584
rect 8444 20544 8450 20556
rect 9490 20544 9496 20556
rect 9548 20584 9554 20596
rect 11330 20584 11336 20596
rect 9548 20556 9674 20584
rect 9548 20544 9554 20556
rect 3878 20476 3884 20528
rect 3936 20516 3942 20528
rect 4246 20516 4252 20528
rect 3936 20488 4252 20516
rect 3936 20476 3942 20488
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 5718 20476 5724 20528
rect 5776 20516 5782 20528
rect 7098 20516 7104 20528
rect 5776 20488 7104 20516
rect 5776 20476 5782 20488
rect 7098 20476 7104 20488
rect 7156 20476 7162 20528
rect 8754 20476 8760 20528
rect 8812 20476 8818 20528
rect 9646 20516 9674 20556
rect 10060 20556 11336 20584
rect 10060 20516 10088 20556
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 12989 20587 13047 20593
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 13035 20556 15792 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 9646 20488 10166 20516
rect 11790 20476 11796 20528
rect 11848 20476 11854 20528
rect 12434 20476 12440 20528
rect 12492 20516 12498 20528
rect 13538 20516 13544 20528
rect 12492 20488 13544 20516
rect 12492 20476 12498 20488
rect 13538 20476 13544 20488
rect 13596 20516 13602 20528
rect 15286 20516 15292 20528
rect 13596 20488 13768 20516
rect 15226 20488 15292 20516
rect 13596 20476 13602 20488
rect 1762 20408 1768 20460
rect 1820 20408 1826 20460
rect 3418 20408 3424 20460
rect 3476 20408 3482 20460
rect 4982 20408 4988 20460
rect 5040 20448 5046 20460
rect 5040 20420 5948 20448
rect 5040 20408 5046 20420
rect 2777 20383 2835 20389
rect 2777 20349 2789 20383
rect 2823 20380 2835 20383
rect 2866 20380 2872 20392
rect 2823 20352 2872 20380
rect 2823 20349 2835 20352
rect 2777 20343 2835 20349
rect 2866 20340 2872 20352
rect 2924 20340 2930 20392
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 5718 20340 5724 20392
rect 5776 20340 5782 20392
rect 5810 20340 5816 20392
rect 5868 20340 5874 20392
rect 5920 20380 5948 20420
rect 6086 20408 6092 20460
rect 6144 20448 6150 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6144 20420 6561 20448
rect 6144 20408 6150 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 7374 20408 7380 20460
rect 7432 20448 7438 20460
rect 9122 20448 9128 20460
rect 7432 20420 9128 20448
rect 7432 20408 7438 20420
rect 9122 20408 9128 20420
rect 9180 20408 9186 20460
rect 13740 20457 13768 20488
rect 15286 20476 15292 20488
rect 15344 20516 15350 20528
rect 15562 20516 15568 20528
rect 15344 20488 15568 20516
rect 15344 20476 15350 20488
rect 15562 20476 15568 20488
rect 15620 20476 15626 20528
rect 15764 20516 15792 20556
rect 16114 20544 16120 20596
rect 16172 20544 16178 20596
rect 16574 20544 16580 20596
rect 16632 20584 16638 20596
rect 16758 20584 16764 20596
rect 16632 20556 16764 20584
rect 16632 20544 16638 20556
rect 16758 20544 16764 20556
rect 16816 20544 16822 20596
rect 16942 20544 16948 20596
rect 17000 20584 17006 20596
rect 17497 20587 17555 20593
rect 17497 20584 17509 20587
rect 17000 20556 17509 20584
rect 17000 20544 17006 20556
rect 17497 20553 17509 20556
rect 17543 20553 17555 20587
rect 17497 20547 17555 20553
rect 18233 20587 18291 20593
rect 18233 20553 18245 20587
rect 18279 20584 18291 20587
rect 18322 20584 18328 20596
rect 18279 20556 18328 20584
rect 18279 20553 18291 20556
rect 18233 20547 18291 20553
rect 18322 20544 18328 20556
rect 18380 20544 18386 20596
rect 18509 20587 18567 20593
rect 18509 20553 18521 20587
rect 18555 20553 18567 20587
rect 18509 20547 18567 20553
rect 18524 20516 18552 20547
rect 18598 20544 18604 20596
rect 18656 20584 18662 20596
rect 18877 20587 18935 20593
rect 18877 20584 18889 20587
rect 18656 20556 18889 20584
rect 18656 20544 18662 20556
rect 18877 20553 18889 20556
rect 18923 20584 18935 20587
rect 19058 20584 19064 20596
rect 18923 20556 19064 20584
rect 18923 20553 18935 20556
rect 18877 20547 18935 20553
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19484 20556 22094 20584
rect 19484 20544 19490 20556
rect 15764 20488 18552 20516
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20417 12955 20451
rect 12897 20411 12955 20417
rect 13725 20451 13783 20457
rect 13725 20417 13737 20451
rect 13771 20417 13783 20451
rect 13725 20411 13783 20417
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 5920 20352 7021 20380
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 7009 20343 7067 20349
rect 8938 20340 8944 20392
rect 8996 20380 9002 20392
rect 9401 20383 9459 20389
rect 9401 20380 9413 20383
rect 8996 20352 9413 20380
rect 8996 20340 9002 20352
rect 9401 20349 9413 20352
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 9677 20383 9735 20389
rect 9677 20349 9689 20383
rect 9723 20380 9735 20383
rect 10962 20380 10968 20392
rect 9723 20352 10968 20380
rect 9723 20349 9735 20352
rect 9677 20343 9735 20349
rect 5626 20272 5632 20324
rect 5684 20312 5690 20324
rect 5684 20284 8892 20312
rect 5684 20272 5690 20284
rect 5261 20247 5319 20253
rect 5261 20213 5273 20247
rect 5307 20244 5319 20247
rect 7098 20244 7104 20256
rect 5307 20216 7104 20244
rect 5307 20213 5319 20216
rect 5261 20207 5319 20213
rect 7098 20204 7104 20216
rect 7156 20204 7162 20256
rect 7374 20204 7380 20256
rect 7432 20244 7438 20256
rect 8018 20244 8024 20256
rect 7432 20216 8024 20244
rect 7432 20204 7438 20216
rect 8018 20204 8024 20216
rect 8076 20204 8082 20256
rect 8386 20204 8392 20256
rect 8444 20204 8450 20256
rect 8864 20253 8892 20284
rect 8849 20247 8907 20253
rect 8849 20213 8861 20247
rect 8895 20213 8907 20247
rect 9416 20244 9444 20343
rect 10962 20340 10968 20352
rect 11020 20340 11026 20392
rect 12437 20383 12495 20389
rect 12437 20349 12449 20383
rect 12483 20380 12495 20383
rect 12526 20380 12532 20392
rect 12483 20352 12532 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 12526 20340 12532 20352
rect 12584 20380 12590 20392
rect 12912 20380 12940 20411
rect 16022 20408 16028 20460
rect 16080 20408 16086 20460
rect 17405 20451 17463 20457
rect 17405 20417 17417 20451
rect 17451 20417 17463 20451
rect 17405 20411 17463 20417
rect 12584 20352 12940 20380
rect 13173 20383 13231 20389
rect 12584 20340 12590 20352
rect 13173 20349 13185 20383
rect 13219 20349 13231 20383
rect 13173 20343 13231 20349
rect 9674 20244 9680 20256
rect 9416 20216 9680 20244
rect 8849 20207 8907 20213
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 11146 20204 11152 20256
rect 11204 20204 11210 20256
rect 11238 20204 11244 20256
rect 11296 20244 11302 20256
rect 11885 20247 11943 20253
rect 11885 20244 11897 20247
rect 11296 20216 11897 20244
rect 11296 20204 11302 20216
rect 11885 20213 11897 20216
rect 11931 20213 11943 20247
rect 11885 20207 11943 20213
rect 12529 20247 12587 20253
rect 12529 20213 12541 20247
rect 12575 20244 12587 20247
rect 12710 20244 12716 20256
rect 12575 20216 12716 20244
rect 12575 20213 12587 20216
rect 12529 20207 12587 20213
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 13188 20244 13216 20343
rect 13998 20340 14004 20392
rect 14056 20380 14062 20392
rect 14734 20380 14740 20392
rect 14056 20352 14740 20380
rect 14056 20340 14062 20352
rect 14734 20340 14740 20352
rect 14792 20380 14798 20392
rect 14792 20352 15148 20380
rect 14792 20340 14798 20352
rect 15120 20324 15148 20352
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 16853 20383 16911 20389
rect 16853 20380 16865 20383
rect 15252 20352 16865 20380
rect 15252 20340 15258 20352
rect 16853 20349 16865 20352
rect 16899 20380 16911 20383
rect 17420 20380 17448 20411
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 19720 20457 19748 20556
rect 21450 20516 21456 20528
rect 21206 20488 21456 20516
rect 21450 20476 21456 20488
rect 21508 20476 21514 20528
rect 22066 20516 22094 20556
rect 22462 20544 22468 20596
rect 22520 20584 22526 20596
rect 23385 20587 23443 20593
rect 23385 20584 23397 20587
rect 22520 20556 23397 20584
rect 22520 20544 22526 20556
rect 23385 20553 23397 20556
rect 23431 20553 23443 20587
rect 23385 20547 23443 20553
rect 23750 20544 23756 20596
rect 23808 20584 23814 20596
rect 24029 20587 24087 20593
rect 24029 20584 24041 20587
rect 23808 20556 24041 20584
rect 23808 20544 23814 20556
rect 24029 20553 24041 20556
rect 24075 20584 24087 20587
rect 24075 20556 25912 20584
rect 24075 20553 24087 20556
rect 24029 20547 24087 20553
rect 22741 20519 22799 20525
rect 22741 20516 22753 20519
rect 22066 20488 22753 20516
rect 22741 20485 22753 20488
rect 22787 20485 22799 20519
rect 22741 20479 22799 20485
rect 24486 20476 24492 20528
rect 24544 20516 24550 20528
rect 25884 20516 25912 20556
rect 26050 20544 26056 20596
rect 26108 20584 26114 20596
rect 26513 20587 26571 20593
rect 26513 20584 26525 20587
rect 26108 20556 26525 20584
rect 26108 20544 26114 20556
rect 26513 20553 26525 20556
rect 26559 20584 26571 20587
rect 27154 20584 27160 20596
rect 26559 20556 27160 20584
rect 26559 20553 26571 20556
rect 26513 20547 26571 20553
rect 27154 20544 27160 20556
rect 27212 20544 27218 20596
rect 27246 20544 27252 20596
rect 27304 20584 27310 20596
rect 27617 20587 27675 20593
rect 27617 20584 27629 20587
rect 27304 20556 27629 20584
rect 27304 20544 27310 20556
rect 27617 20553 27629 20556
rect 27663 20553 27675 20587
rect 27617 20547 27675 20553
rect 29546 20544 29552 20596
rect 29604 20584 29610 20596
rect 29604 20556 29960 20584
rect 29604 20544 29610 20556
rect 26142 20516 26148 20528
rect 24544 20488 25070 20516
rect 25884 20488 26148 20516
rect 24544 20476 24550 20488
rect 26142 20476 26148 20488
rect 26200 20476 26206 20528
rect 27172 20516 27200 20544
rect 29932 20516 29960 20556
rect 30926 20544 30932 20596
rect 30984 20584 30990 20596
rect 30984 20556 31754 20584
rect 30984 20544 30990 20556
rect 31573 20519 31631 20525
rect 31573 20516 31585 20519
rect 27172 20488 27660 20516
rect 29932 20488 31585 20516
rect 18969 20451 19027 20457
rect 18969 20448 18981 20451
rect 17644 20420 18981 20448
rect 17644 20408 17650 20420
rect 18969 20417 18981 20420
rect 19015 20417 19027 20451
rect 18969 20411 19027 20417
rect 19705 20451 19763 20457
rect 19705 20417 19717 20451
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 22002 20408 22008 20460
rect 22060 20408 22066 20460
rect 23382 20408 23388 20460
rect 23440 20448 23446 20460
rect 24210 20448 24216 20460
rect 23440 20420 24216 20448
rect 23440 20408 23446 20420
rect 24210 20408 24216 20420
rect 24268 20448 24274 20460
rect 24305 20451 24363 20457
rect 24305 20448 24317 20451
rect 24268 20420 24317 20448
rect 24268 20408 24274 20420
rect 24305 20417 24317 20420
rect 24351 20417 24363 20451
rect 24305 20411 24363 20417
rect 25866 20408 25872 20460
rect 25924 20448 25930 20460
rect 26789 20451 26847 20457
rect 26789 20448 26801 20451
rect 25924 20420 26801 20448
rect 25924 20408 25930 20420
rect 26789 20417 26801 20420
rect 26835 20448 26847 20451
rect 27522 20448 27528 20460
rect 26835 20420 27528 20448
rect 26835 20417 26847 20420
rect 26789 20411 26847 20417
rect 27522 20408 27528 20420
rect 27580 20408 27586 20460
rect 27632 20448 27660 20488
rect 31573 20485 31585 20488
rect 31619 20485 31631 20519
rect 31726 20516 31754 20556
rect 32125 20519 32183 20525
rect 32125 20516 32137 20519
rect 31726 20488 32137 20516
rect 31573 20479 31631 20485
rect 32125 20485 32137 20488
rect 32171 20485 32183 20519
rect 32125 20479 32183 20485
rect 27632 20420 27844 20448
rect 16899 20352 17448 20380
rect 17681 20383 17739 20389
rect 16899 20349 16911 20352
rect 16853 20343 16911 20349
rect 17681 20349 17693 20383
rect 17727 20380 17739 20383
rect 18782 20380 18788 20392
rect 17727 20352 18788 20380
rect 17727 20349 17739 20352
rect 17681 20343 17739 20349
rect 18782 20340 18788 20352
rect 18840 20340 18846 20392
rect 19061 20383 19119 20389
rect 19061 20349 19073 20383
rect 19107 20349 19119 20383
rect 19061 20343 19119 20349
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 20622 20380 20628 20392
rect 20027 20352 20628 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 15102 20272 15108 20324
rect 15160 20272 15166 20324
rect 16574 20312 16580 20324
rect 15396 20284 16580 20312
rect 15396 20244 15424 20284
rect 16574 20272 16580 20284
rect 16632 20272 16638 20324
rect 16758 20272 16764 20324
rect 16816 20312 16822 20324
rect 17037 20315 17095 20321
rect 17037 20312 17049 20315
rect 16816 20284 17049 20312
rect 16816 20272 16822 20284
rect 17037 20281 17049 20284
rect 17083 20281 17095 20315
rect 17037 20275 17095 20281
rect 17494 20272 17500 20324
rect 17552 20312 17558 20324
rect 19076 20312 19104 20343
rect 20622 20340 20628 20352
rect 20680 20340 20686 20392
rect 24581 20383 24639 20389
rect 24581 20349 24593 20383
rect 24627 20380 24639 20383
rect 24670 20380 24676 20392
rect 24627 20352 24676 20380
rect 24627 20349 24639 20352
rect 24581 20343 24639 20349
rect 24670 20340 24676 20352
rect 24728 20340 24734 20392
rect 25958 20340 25964 20392
rect 26016 20380 26022 20392
rect 26053 20383 26111 20389
rect 26053 20380 26065 20383
rect 26016 20352 26065 20380
rect 26016 20340 26022 20352
rect 26053 20349 26065 20352
rect 26099 20380 26111 20383
rect 27709 20383 27767 20389
rect 27709 20380 27721 20383
rect 26099 20352 27721 20380
rect 26099 20349 26111 20352
rect 26053 20343 26111 20349
rect 27709 20349 27721 20352
rect 27755 20349 27767 20383
rect 27816 20380 27844 20420
rect 29730 20408 29736 20460
rect 29788 20408 29794 20460
rect 31021 20451 31079 20457
rect 31021 20417 31033 20451
rect 31067 20448 31079 20451
rect 36906 20448 36912 20460
rect 31067 20420 36912 20448
rect 31067 20417 31079 20420
rect 31021 20411 31079 20417
rect 36906 20408 36912 20420
rect 36964 20408 36970 20460
rect 28350 20380 28356 20392
rect 27816 20352 28356 20380
rect 27709 20343 27767 20349
rect 28350 20340 28356 20352
rect 28408 20340 28414 20392
rect 28629 20383 28687 20389
rect 28629 20349 28641 20383
rect 28675 20380 28687 20383
rect 30190 20380 30196 20392
rect 28675 20352 30196 20380
rect 28675 20349 28687 20352
rect 28629 20343 28687 20349
rect 30190 20340 30196 20352
rect 30248 20340 30254 20392
rect 30282 20340 30288 20392
rect 30340 20380 30346 20392
rect 31113 20383 31171 20389
rect 31113 20380 31125 20383
rect 30340 20352 31125 20380
rect 30340 20340 30346 20352
rect 31113 20349 31125 20352
rect 31159 20349 31171 20383
rect 31113 20343 31171 20349
rect 31478 20340 31484 20392
rect 31536 20380 31542 20392
rect 31757 20383 31815 20389
rect 31757 20380 31769 20383
rect 31536 20352 31769 20380
rect 31536 20340 31542 20352
rect 31757 20349 31769 20352
rect 31803 20349 31815 20383
rect 31757 20343 31815 20349
rect 17552 20284 19104 20312
rect 17552 20272 17558 20284
rect 13188 20216 15424 20244
rect 15470 20204 15476 20256
rect 15528 20204 15534 20256
rect 15562 20204 15568 20256
rect 15620 20244 15626 20256
rect 16114 20244 16120 20256
rect 15620 20216 16120 20244
rect 15620 20204 15626 20216
rect 16114 20204 16120 20216
rect 16172 20244 16178 20256
rect 16669 20247 16727 20253
rect 16669 20244 16681 20247
rect 16172 20216 16681 20244
rect 16172 20204 16178 20216
rect 16669 20213 16681 20216
rect 16715 20244 16727 20247
rect 18322 20244 18328 20256
rect 16715 20216 18328 20244
rect 16715 20213 16727 20216
rect 16669 20207 16727 20213
rect 18322 20204 18328 20216
rect 18380 20204 18386 20256
rect 19076 20244 19104 20284
rect 22554 20272 22560 20324
rect 22612 20312 22618 20324
rect 27157 20315 27215 20321
rect 27157 20312 27169 20315
rect 22612 20284 24440 20312
rect 22612 20272 22618 20284
rect 21453 20247 21511 20253
rect 21453 20244 21465 20247
rect 19076 20216 21465 20244
rect 21453 20213 21465 20216
rect 21499 20213 21511 20247
rect 24412 20244 24440 20284
rect 25608 20284 27169 20312
rect 25608 20244 25636 20284
rect 27157 20281 27169 20284
rect 27203 20281 27215 20315
rect 27157 20275 27215 20281
rect 27614 20272 27620 20324
rect 27672 20312 27678 20324
rect 27890 20312 27896 20324
rect 27672 20284 27896 20312
rect 27672 20272 27678 20284
rect 27890 20272 27896 20284
rect 27948 20272 27954 20324
rect 24412 20216 25636 20244
rect 21453 20207 21511 20213
rect 25682 20204 25688 20256
rect 25740 20244 25746 20256
rect 26421 20247 26479 20253
rect 26421 20244 26433 20247
rect 25740 20216 26433 20244
rect 25740 20204 25746 20216
rect 26421 20213 26433 20216
rect 26467 20244 26479 20247
rect 26510 20244 26516 20256
rect 26467 20216 26516 20244
rect 26467 20213 26479 20216
rect 26421 20207 26479 20213
rect 26510 20204 26516 20216
rect 26568 20204 26574 20256
rect 27706 20204 27712 20256
rect 27764 20244 27770 20256
rect 28626 20244 28632 20256
rect 27764 20216 28632 20244
rect 27764 20204 27770 20216
rect 28626 20204 28632 20216
rect 28684 20244 28690 20256
rect 30101 20247 30159 20253
rect 30101 20244 30113 20247
rect 28684 20216 30113 20244
rect 28684 20204 28690 20216
rect 30101 20213 30113 20216
rect 30147 20213 30159 20247
rect 30101 20207 30159 20213
rect 30190 20204 30196 20256
rect 30248 20244 30254 20256
rect 30561 20247 30619 20253
rect 30561 20244 30573 20247
rect 30248 20216 30573 20244
rect 30248 20204 30254 20216
rect 30561 20213 30573 20216
rect 30607 20213 30619 20247
rect 30561 20207 30619 20213
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 3326 20000 3332 20052
rect 3384 20040 3390 20052
rect 3789 20043 3847 20049
rect 3789 20040 3801 20043
rect 3384 20012 3801 20040
rect 3384 20000 3390 20012
rect 3789 20009 3801 20012
rect 3835 20040 3847 20043
rect 3973 20043 4031 20049
rect 3973 20040 3985 20043
rect 3835 20012 3985 20040
rect 3835 20009 3847 20012
rect 3789 20003 3847 20009
rect 3973 20009 3985 20012
rect 4019 20040 4031 20043
rect 4157 20043 4215 20049
rect 4157 20040 4169 20043
rect 4019 20012 4169 20040
rect 4019 20009 4031 20012
rect 3973 20003 4031 20009
rect 4157 20009 4169 20012
rect 4203 20040 4215 20043
rect 5258 20040 5264 20052
rect 4203 20012 5264 20040
rect 4203 20009 4215 20012
rect 4157 20003 4215 20009
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 6273 20043 6331 20049
rect 6273 20009 6285 20043
rect 6319 20040 6331 20043
rect 7558 20040 7564 20052
rect 6319 20012 7564 20040
rect 6319 20009 6331 20012
rect 6273 20003 6331 20009
rect 7558 20000 7564 20012
rect 7616 20000 7622 20052
rect 8018 20000 8024 20052
rect 8076 20040 8082 20052
rect 8481 20043 8539 20049
rect 8481 20040 8493 20043
rect 8076 20012 8493 20040
rect 8076 20000 8082 20012
rect 8481 20009 8493 20012
rect 8527 20009 8539 20043
rect 8481 20003 8539 20009
rect 8570 20000 8576 20052
rect 8628 20040 8634 20052
rect 9858 20040 9864 20052
rect 8628 20012 9864 20040
rect 8628 20000 8634 20012
rect 9858 20000 9864 20012
rect 9916 20040 9922 20052
rect 10873 20043 10931 20049
rect 10873 20040 10885 20043
rect 9916 20012 10885 20040
rect 9916 20000 9922 20012
rect 10873 20009 10885 20012
rect 10919 20009 10931 20043
rect 10873 20003 10931 20009
rect 11330 20000 11336 20052
rect 11388 20040 11394 20052
rect 11425 20043 11483 20049
rect 11425 20040 11437 20043
rect 11388 20012 11437 20040
rect 11388 20000 11394 20012
rect 11425 20009 11437 20012
rect 11471 20040 11483 20043
rect 11882 20040 11888 20052
rect 11471 20012 11888 20040
rect 11471 20009 11483 20012
rect 11425 20003 11483 20009
rect 11882 20000 11888 20012
rect 11940 20000 11946 20052
rect 12989 20043 13047 20049
rect 12989 20009 13001 20043
rect 13035 20040 13047 20043
rect 13814 20040 13820 20052
rect 13035 20012 13820 20040
rect 13035 20009 13047 20012
rect 12989 20003 13047 20009
rect 13814 20000 13820 20012
rect 13872 20000 13878 20052
rect 14182 20000 14188 20052
rect 14240 20040 14246 20052
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 14240 20012 14289 20040
rect 14240 20000 14246 20012
rect 14277 20009 14289 20012
rect 14323 20040 14335 20043
rect 17586 20040 17592 20052
rect 14323 20012 17592 20040
rect 14323 20009 14335 20012
rect 14277 20003 14335 20009
rect 17586 20000 17592 20012
rect 17644 20000 17650 20052
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 19794 20040 19800 20052
rect 18739 20012 19800 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 19794 20000 19800 20012
rect 19852 20000 19858 20052
rect 21266 20000 21272 20052
rect 21324 20040 21330 20052
rect 24578 20040 24584 20052
rect 21324 20012 24584 20040
rect 21324 20000 21330 20012
rect 24578 20000 24584 20012
rect 24636 20000 24642 20052
rect 30745 20043 30803 20049
rect 30745 20040 30757 20043
rect 25148 20012 30757 20040
rect 12434 19972 12440 19984
rect 10796 19944 12440 19972
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 3326 19904 3332 19916
rect 2823 19876 3332 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 3326 19864 3332 19876
rect 3384 19864 3390 19916
rect 4525 19907 4583 19913
rect 4525 19873 4537 19907
rect 4571 19904 4583 19907
rect 5442 19904 5448 19916
rect 4571 19876 5448 19904
rect 4571 19873 4583 19876
rect 4525 19867 4583 19873
rect 5442 19864 5448 19876
rect 5500 19904 5506 19916
rect 6733 19907 6791 19913
rect 6733 19904 6745 19907
rect 5500 19876 6745 19904
rect 5500 19864 5506 19876
rect 6733 19873 6745 19876
rect 6779 19904 6791 19907
rect 8938 19904 8944 19916
rect 6779 19876 8944 19904
rect 6779 19873 6791 19876
rect 6733 19867 6791 19873
rect 8938 19864 8944 19876
rect 8996 19864 9002 19916
rect 9125 19907 9183 19913
rect 9125 19873 9137 19907
rect 9171 19904 9183 19907
rect 10796 19904 10824 19944
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 16761 19975 16819 19981
rect 16761 19941 16773 19975
rect 16807 19972 16819 19975
rect 17034 19972 17040 19984
rect 16807 19944 17040 19972
rect 16807 19941 16819 19944
rect 16761 19935 16819 19941
rect 17034 19932 17040 19944
rect 17092 19932 17098 19984
rect 17218 19932 17224 19984
rect 17276 19932 17282 19984
rect 18966 19972 18972 19984
rect 17880 19944 18972 19972
rect 9171 19876 10824 19904
rect 12345 19907 12403 19913
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 12345 19873 12357 19907
rect 12391 19904 12403 19907
rect 13354 19904 13360 19916
rect 12391 19876 13360 19904
rect 12391 19873 12403 19876
rect 12345 19867 12403 19873
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 13633 19907 13691 19913
rect 13633 19873 13645 19907
rect 13679 19904 13691 19907
rect 14829 19907 14887 19913
rect 14829 19904 14841 19907
rect 13679 19876 14841 19904
rect 13679 19873 13691 19876
rect 13633 19867 13691 19873
rect 14829 19873 14841 19876
rect 14875 19904 14887 19907
rect 15470 19904 15476 19916
rect 14875 19876 15476 19904
rect 14875 19873 14887 19876
rect 14829 19867 14887 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 16942 19864 16948 19916
rect 17000 19864 17006 19916
rect 17678 19864 17684 19916
rect 17736 19864 17742 19916
rect 17880 19913 17908 19944
rect 18966 19932 18972 19944
rect 19024 19972 19030 19984
rect 19242 19972 19248 19984
rect 19024 19944 19248 19972
rect 19024 19932 19030 19944
rect 19242 19932 19248 19944
rect 19300 19932 19306 19984
rect 22830 19932 22836 19984
rect 22888 19972 22894 19984
rect 24673 19975 24731 19981
rect 24673 19972 24685 19975
rect 22888 19944 24685 19972
rect 22888 19932 22894 19944
rect 24673 19941 24685 19944
rect 24719 19941 24731 19975
rect 24673 19935 24731 19941
rect 17865 19907 17923 19913
rect 17865 19873 17877 19907
rect 17911 19873 17923 19907
rect 17865 19867 17923 19873
rect 18782 19864 18788 19916
rect 18840 19904 18846 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 18840 19876 20545 19904
rect 18840 19864 18846 19876
rect 20533 19873 20545 19876
rect 20579 19904 20591 19907
rect 21174 19904 21180 19916
rect 20579 19876 21180 19904
rect 20579 19873 20591 19876
rect 20533 19867 20591 19873
rect 21174 19864 21180 19876
rect 21232 19864 21238 19916
rect 23842 19904 23848 19916
rect 22020 19876 23848 19904
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19836 1823 19839
rect 4062 19836 4068 19848
rect 1811 19808 4068 19836
rect 1811 19805 1823 19808
rect 1765 19799 1823 19805
rect 4062 19796 4068 19808
rect 4120 19796 4126 19848
rect 11054 19796 11060 19848
rect 11112 19836 11118 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 11112 19808 12173 19836
rect 11112 19796 11118 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12253 19839 12311 19845
rect 12253 19805 12265 19839
rect 12299 19836 12311 19839
rect 14458 19836 14464 19848
rect 12299 19808 14464 19836
rect 12299 19805 12311 19808
rect 12253 19799 12311 19805
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 17589 19839 17647 19845
rect 17589 19805 17601 19839
rect 17635 19836 17647 19839
rect 18877 19839 18935 19845
rect 17635 19808 18828 19836
rect 17635 19805 17647 19808
rect 17589 19799 17647 19805
rect 3605 19771 3663 19777
rect 3605 19737 3617 19771
rect 3651 19768 3663 19771
rect 3878 19768 3884 19780
rect 3651 19740 3884 19768
rect 3651 19737 3663 19740
rect 3605 19731 3663 19737
rect 3878 19728 3884 19740
rect 3936 19728 3942 19780
rect 4798 19728 4804 19780
rect 4856 19728 4862 19780
rect 5258 19728 5264 19780
rect 5316 19728 5322 19780
rect 6730 19728 6736 19780
rect 6788 19768 6794 19780
rect 7009 19771 7067 19777
rect 7009 19768 7021 19771
rect 6788 19740 7021 19768
rect 6788 19728 6794 19740
rect 7009 19737 7021 19740
rect 7055 19737 7067 19771
rect 7009 19731 7067 19737
rect 7466 19728 7472 19780
rect 7524 19728 7530 19780
rect 9401 19771 9459 19777
rect 9401 19737 9413 19771
rect 9447 19737 9459 19771
rect 9401 19731 9459 19737
rect 3694 19660 3700 19712
rect 3752 19700 3758 19712
rect 6914 19700 6920 19712
rect 3752 19672 6920 19700
rect 3752 19660 3758 19672
rect 6914 19660 6920 19672
rect 6972 19660 6978 19712
rect 9416 19700 9444 19731
rect 9490 19728 9496 19780
rect 9548 19768 9554 19780
rect 11146 19768 11152 19780
rect 9548 19740 9890 19768
rect 10704 19740 11152 19768
rect 9548 19728 9554 19740
rect 10704 19700 10732 19740
rect 11146 19728 11152 19740
rect 11204 19728 11210 19780
rect 13262 19768 13268 19780
rect 11256 19740 13268 19768
rect 9416 19672 10732 19700
rect 10962 19660 10968 19712
rect 11020 19700 11026 19712
rect 11256 19700 11284 19740
rect 13262 19728 13268 19740
rect 13320 19728 13326 19780
rect 13449 19771 13507 19777
rect 13449 19737 13461 19771
rect 13495 19768 13507 19771
rect 16114 19768 16120 19780
rect 13495 19740 15240 19768
rect 16054 19740 16120 19768
rect 13495 19737 13507 19740
rect 13449 19731 13507 19737
rect 11020 19672 11284 19700
rect 11020 19660 11026 19672
rect 11790 19660 11796 19712
rect 11848 19660 11854 19712
rect 11882 19660 11888 19712
rect 11940 19700 11946 19712
rect 13170 19700 13176 19712
rect 11940 19672 13176 19700
rect 11940 19660 11946 19672
rect 13170 19660 13176 19672
rect 13228 19660 13234 19712
rect 13354 19660 13360 19712
rect 13412 19660 13418 19712
rect 14182 19660 14188 19712
rect 14240 19700 14246 19712
rect 15010 19700 15016 19712
rect 14240 19672 15016 19700
rect 14240 19660 14246 19672
rect 15010 19660 15016 19672
rect 15068 19660 15074 19712
rect 15212 19700 15240 19740
rect 16114 19728 16120 19740
rect 16172 19728 16178 19780
rect 18322 19768 18328 19780
rect 16224 19740 18328 19768
rect 16224 19700 16252 19740
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 18800 19768 18828 19808
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19058 19836 19064 19848
rect 18923 19808 19064 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19058 19796 19064 19808
rect 19116 19796 19122 19848
rect 19702 19796 19708 19848
rect 19760 19836 19766 19848
rect 20257 19839 20315 19845
rect 20257 19836 20269 19839
rect 19760 19808 20269 19836
rect 19760 19796 19766 19808
rect 20257 19805 20269 19808
rect 20303 19805 20315 19839
rect 20257 19799 20315 19805
rect 19426 19768 19432 19780
rect 18800 19740 19432 19768
rect 19426 19728 19432 19740
rect 19484 19728 19490 19780
rect 19518 19728 19524 19780
rect 19576 19768 19582 19780
rect 19613 19771 19671 19777
rect 19613 19768 19625 19771
rect 19576 19740 19625 19768
rect 19576 19728 19582 19740
rect 19613 19737 19625 19740
rect 19659 19768 19671 19771
rect 20438 19768 20444 19780
rect 19659 19740 20444 19768
rect 19659 19737 19671 19740
rect 19613 19731 19671 19737
rect 20438 19728 20444 19740
rect 20496 19728 20502 19780
rect 21542 19728 21548 19780
rect 21600 19728 21606 19780
rect 15212 19672 16252 19700
rect 16301 19703 16359 19709
rect 16301 19669 16313 19703
rect 16347 19700 16359 19703
rect 16390 19700 16396 19712
rect 16347 19672 16396 19700
rect 16347 19669 16359 19672
rect 16301 19663 16359 19669
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 18414 19660 18420 19712
rect 18472 19660 18478 19712
rect 19705 19703 19763 19709
rect 19705 19669 19717 19703
rect 19751 19700 19763 19703
rect 19886 19700 19892 19712
rect 19751 19672 19892 19700
rect 19751 19669 19763 19672
rect 19705 19663 19763 19669
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 21450 19660 21456 19712
rect 21508 19700 21514 19712
rect 22020 19709 22048 19876
rect 23842 19864 23848 19876
rect 23900 19864 23906 19916
rect 25148 19913 25176 20012
rect 30745 20009 30757 20012
rect 30791 20009 30803 20043
rect 30745 20003 30803 20009
rect 30834 20000 30840 20052
rect 30892 20040 30898 20052
rect 49234 20040 49240 20052
rect 30892 20012 49240 20040
rect 30892 20000 30898 20012
rect 49234 20000 49240 20012
rect 49292 20000 49298 20052
rect 27982 19932 27988 19984
rect 28040 19972 28046 19984
rect 29638 19972 29644 19984
rect 28040 19944 29644 19972
rect 28040 19932 28046 19944
rect 29638 19932 29644 19944
rect 29696 19932 29702 19984
rect 29733 19975 29791 19981
rect 29733 19941 29745 19975
rect 29779 19972 29791 19975
rect 33502 19972 33508 19984
rect 29779 19944 33508 19972
rect 29779 19941 29791 19944
rect 29733 19935 29791 19941
rect 33502 19932 33508 19944
rect 33560 19932 33566 19984
rect 25133 19907 25191 19913
rect 25133 19873 25145 19907
rect 25179 19873 25191 19907
rect 25133 19867 25191 19873
rect 25222 19864 25228 19916
rect 25280 19864 25286 19916
rect 28629 19907 28687 19913
rect 28629 19904 28641 19907
rect 25332 19876 28641 19904
rect 22278 19796 22284 19848
rect 22336 19836 22342 19848
rect 22557 19839 22615 19845
rect 22557 19836 22569 19839
rect 22336 19808 22569 19836
rect 22336 19796 22342 19808
rect 22557 19805 22569 19808
rect 22603 19805 22615 19839
rect 22557 19799 22615 19805
rect 23750 19796 23756 19848
rect 23808 19796 23814 19848
rect 24762 19796 24768 19848
rect 24820 19836 24826 19848
rect 25332 19836 25360 19876
rect 28629 19873 28641 19876
rect 28675 19873 28687 19907
rect 28629 19867 28687 19873
rect 28718 19864 28724 19916
rect 28776 19904 28782 19916
rect 31297 19907 31355 19913
rect 31297 19904 31309 19907
rect 28776 19876 31309 19904
rect 28776 19864 28782 19876
rect 31297 19873 31309 19876
rect 31343 19873 31355 19907
rect 31297 19867 31355 19873
rect 24820 19808 25360 19836
rect 24820 19796 24826 19808
rect 25774 19796 25780 19848
rect 25832 19836 25838 19848
rect 25869 19839 25927 19845
rect 25869 19836 25881 19839
rect 25832 19808 25881 19836
rect 25832 19796 25838 19808
rect 25869 19805 25881 19808
rect 25915 19805 25927 19839
rect 25869 19799 25927 19805
rect 27246 19796 27252 19848
rect 27304 19836 27310 19848
rect 27893 19839 27951 19845
rect 27893 19836 27905 19839
rect 27304 19808 27905 19836
rect 27304 19796 27310 19808
rect 27893 19805 27905 19808
rect 27939 19836 27951 19839
rect 27982 19836 27988 19848
rect 27939 19808 27988 19836
rect 27939 19805 27951 19808
rect 27893 19799 27951 19805
rect 27982 19796 27988 19808
rect 28040 19796 28046 19848
rect 28353 19839 28411 19845
rect 28353 19805 28365 19839
rect 28399 19836 28411 19839
rect 28534 19836 28540 19848
rect 28399 19808 28540 19836
rect 28399 19805 28411 19808
rect 28353 19799 28411 19805
rect 28534 19796 28540 19808
rect 28592 19796 28598 19848
rect 29914 19796 29920 19848
rect 29972 19836 29978 19848
rect 30193 19839 30251 19845
rect 30193 19836 30205 19839
rect 29972 19808 30205 19836
rect 29972 19796 29978 19808
rect 30193 19805 30205 19808
rect 30239 19805 30251 19839
rect 30193 19799 30251 19805
rect 31205 19839 31263 19845
rect 31205 19805 31217 19839
rect 31251 19836 31263 19839
rect 37182 19836 37188 19848
rect 31251 19808 37188 19836
rect 31251 19805 31263 19808
rect 31205 19799 31263 19805
rect 37182 19796 37188 19808
rect 37240 19796 37246 19848
rect 22738 19728 22744 19780
rect 22796 19728 22802 19780
rect 23566 19728 23572 19780
rect 23624 19768 23630 19780
rect 26142 19768 26148 19780
rect 23624 19740 26148 19768
rect 23624 19728 23630 19740
rect 26142 19728 26148 19740
rect 26200 19728 26206 19780
rect 26602 19728 26608 19780
rect 26660 19728 26666 19780
rect 30834 19768 30840 19780
rect 27448 19740 30840 19768
rect 22005 19703 22063 19709
rect 22005 19700 22017 19703
rect 21508 19672 22017 19700
rect 21508 19660 21514 19672
rect 22005 19669 22017 19672
rect 22051 19669 22063 19703
rect 22005 19663 22063 19669
rect 23290 19660 23296 19712
rect 23348 19660 23354 19712
rect 23658 19660 23664 19712
rect 23716 19660 23722 19712
rect 25038 19660 25044 19712
rect 25096 19660 25102 19712
rect 25866 19660 25872 19712
rect 25924 19700 25930 19712
rect 27448 19700 27476 19740
rect 30834 19728 30840 19740
rect 30892 19728 30898 19780
rect 25924 19672 27476 19700
rect 27617 19703 27675 19709
rect 25924 19660 25930 19672
rect 27617 19669 27629 19703
rect 27663 19700 27675 19703
rect 27890 19700 27896 19712
rect 27663 19672 27896 19700
rect 27663 19669 27675 19672
rect 27617 19663 27675 19669
rect 27890 19660 27896 19672
rect 27948 19660 27954 19712
rect 28350 19660 28356 19712
rect 28408 19700 28414 19712
rect 30377 19703 30435 19709
rect 30377 19700 30389 19703
rect 28408 19672 30389 19700
rect 28408 19660 28414 19672
rect 30377 19669 30389 19672
rect 30423 19700 30435 19703
rect 30466 19700 30472 19712
rect 30423 19672 30472 19700
rect 30423 19669 30435 19672
rect 30377 19663 30435 19669
rect 30466 19660 30472 19672
rect 30524 19700 30530 19712
rect 31113 19703 31171 19709
rect 31113 19700 31125 19703
rect 30524 19672 31125 19700
rect 30524 19660 30530 19672
rect 31113 19669 31125 19672
rect 31159 19669 31171 19703
rect 31113 19663 31171 19669
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 4890 19496 4896 19508
rect 2746 19468 4896 19496
rect 2746 19428 2774 19468
rect 4890 19456 4896 19468
rect 4948 19456 4954 19508
rect 4982 19456 4988 19508
rect 5040 19496 5046 19508
rect 5261 19499 5319 19505
rect 5261 19496 5273 19499
rect 5040 19468 5273 19496
rect 5040 19456 5046 19468
rect 5261 19465 5273 19468
rect 5307 19465 5319 19499
rect 5261 19459 5319 19465
rect 5721 19499 5779 19505
rect 5721 19465 5733 19499
rect 5767 19496 5779 19499
rect 5994 19496 6000 19508
rect 5767 19468 6000 19496
rect 5767 19465 5779 19468
rect 5721 19459 5779 19465
rect 5994 19456 6000 19468
rect 6052 19456 6058 19508
rect 10318 19496 10324 19508
rect 7484 19468 10324 19496
rect 1780 19400 2774 19428
rect 1780 19369 1808 19400
rect 4154 19388 4160 19440
rect 4212 19428 4218 19440
rect 4341 19431 4399 19437
rect 4341 19428 4353 19431
rect 4212 19400 4353 19428
rect 4212 19388 4218 19400
rect 4341 19397 4353 19400
rect 4387 19397 4399 19431
rect 4341 19391 4399 19397
rect 5629 19431 5687 19437
rect 5629 19397 5641 19431
rect 5675 19428 5687 19431
rect 7484 19428 7512 19468
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 10413 19499 10471 19505
rect 10413 19465 10425 19499
rect 10459 19465 10471 19499
rect 10413 19459 10471 19465
rect 5675 19400 7512 19428
rect 5675 19397 5687 19400
rect 5629 19391 5687 19397
rect 7558 19388 7564 19440
rect 7616 19428 7622 19440
rect 9309 19431 9367 19437
rect 9309 19428 9321 19431
rect 7616 19400 9321 19428
rect 7616 19388 7622 19400
rect 9309 19397 9321 19400
rect 9355 19397 9367 19431
rect 10428 19428 10456 19459
rect 10870 19456 10876 19508
rect 10928 19456 10934 19508
rect 12158 19456 12164 19508
rect 12216 19496 12222 19508
rect 14550 19496 14556 19508
rect 12216 19468 14556 19496
rect 12216 19456 12222 19468
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 14826 19456 14832 19508
rect 14884 19456 14890 19508
rect 17221 19499 17279 19505
rect 17221 19465 17233 19499
rect 17267 19496 17279 19499
rect 17402 19496 17408 19508
rect 17267 19468 17408 19496
rect 17267 19465 17279 19468
rect 17221 19459 17279 19465
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 17865 19499 17923 19505
rect 17865 19496 17877 19499
rect 17512 19468 17877 19496
rect 11422 19428 11428 19440
rect 10428 19400 11428 19428
rect 9309 19391 9367 19397
rect 11422 19388 11428 19400
rect 11480 19388 11486 19440
rect 11882 19428 11888 19440
rect 11716 19400 11888 19428
rect 1765 19363 1823 19369
rect 1765 19329 1777 19363
rect 1811 19329 1823 19363
rect 1765 19323 1823 19329
rect 2777 19363 2835 19369
rect 2777 19329 2789 19363
rect 2823 19360 2835 19363
rect 2866 19360 2872 19372
rect 2823 19332 2872 19360
rect 2823 19329 2835 19332
rect 2777 19323 2835 19329
rect 2866 19320 2872 19332
rect 2924 19320 2930 19372
rect 3602 19320 3608 19372
rect 3660 19320 3666 19372
rect 5258 19320 5264 19372
rect 5316 19360 5322 19372
rect 6641 19363 6699 19369
rect 5316 19346 5488 19360
rect 5316 19332 5448 19346
rect 5316 19320 5322 19332
rect 5442 19294 5448 19332
rect 5500 19294 5506 19346
rect 6641 19334 6653 19363
rect 6564 19329 6653 19334
rect 6687 19329 6699 19363
rect 6564 19323 6699 19329
rect 6564 19306 6684 19323
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 7469 19363 7527 19369
rect 7469 19360 7481 19363
rect 6972 19332 7481 19360
rect 6972 19320 6978 19332
rect 7469 19329 7481 19332
rect 7515 19329 7527 19363
rect 7469 19323 7527 19329
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19360 8631 19363
rect 8662 19360 8668 19372
rect 8619 19332 8668 19360
rect 8619 19329 8631 19332
rect 8573 19323 8631 19329
rect 8662 19320 8668 19332
rect 8720 19320 8726 19372
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19360 10379 19363
rect 10778 19360 10784 19372
rect 10367 19332 10784 19360
rect 10367 19329 10379 19332
rect 10321 19323 10379 19329
rect 10778 19320 10784 19332
rect 10836 19320 10842 19372
rect 11716 19369 11744 19400
rect 11882 19388 11888 19400
rect 11940 19388 11946 19440
rect 14458 19388 14464 19440
rect 14516 19428 14522 19440
rect 17512 19428 17540 19468
rect 17865 19465 17877 19468
rect 17911 19465 17923 19499
rect 18966 19496 18972 19508
rect 17865 19459 17923 19465
rect 17972 19468 18972 19496
rect 14516 19400 17540 19428
rect 14516 19388 14522 19400
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 5902 19252 5908 19304
rect 5960 19252 5966 19304
rect 5350 19184 5356 19236
rect 5408 19224 5414 19236
rect 6564 19224 6592 19306
rect 10962 19252 10968 19304
rect 11020 19252 11026 19304
rect 11977 19295 12035 19301
rect 11977 19261 11989 19295
rect 12023 19292 12035 19295
rect 12342 19292 12348 19304
rect 12023 19264 12348 19292
rect 12023 19261 12035 19264
rect 11977 19255 12035 19261
rect 12342 19252 12348 19264
rect 12400 19252 12406 19304
rect 13096 19292 13124 19346
rect 13262 19320 13268 19372
rect 13320 19360 13326 19372
rect 13320 19332 13492 19360
rect 13320 19320 13326 19332
rect 13170 19292 13176 19304
rect 13096 19264 13176 19292
rect 13170 19252 13176 19264
rect 13228 19252 13234 19304
rect 13464 19301 13492 19332
rect 14090 19320 14096 19372
rect 14148 19360 14154 19372
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 14148 19332 14749 19360
rect 14148 19320 14154 19332
rect 14737 19329 14749 19332
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 15654 19320 15660 19372
rect 15712 19320 15718 19372
rect 17310 19320 17316 19372
rect 17368 19360 17374 19372
rect 17405 19363 17463 19369
rect 17405 19360 17417 19363
rect 17368 19332 17417 19360
rect 17368 19320 17374 19332
rect 17405 19329 17417 19332
rect 17451 19329 17463 19363
rect 17405 19323 17463 19329
rect 17494 19320 17500 19372
rect 17552 19360 17558 19372
rect 17972 19360 18000 19468
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 19058 19456 19064 19508
rect 19116 19456 19122 19508
rect 19242 19456 19248 19508
rect 19300 19496 19306 19508
rect 21453 19499 21511 19505
rect 21453 19496 21465 19499
rect 19300 19468 21465 19496
rect 19300 19456 19306 19468
rect 21453 19465 21465 19468
rect 21499 19465 21511 19499
rect 21453 19459 21511 19465
rect 22373 19499 22431 19505
rect 22373 19465 22385 19499
rect 22419 19496 22431 19499
rect 23290 19496 23296 19508
rect 22419 19468 23296 19496
rect 22419 19465 22431 19468
rect 22373 19459 22431 19465
rect 23290 19456 23296 19468
rect 23348 19456 23354 19508
rect 23566 19456 23572 19508
rect 23624 19496 23630 19508
rect 23661 19499 23719 19505
rect 23661 19496 23673 19499
rect 23624 19468 23673 19496
rect 23624 19456 23630 19468
rect 23661 19465 23673 19468
rect 23707 19465 23719 19499
rect 25866 19496 25872 19508
rect 23661 19459 23719 19465
rect 23952 19468 25872 19496
rect 18046 19388 18052 19440
rect 18104 19428 18110 19440
rect 18325 19431 18383 19437
rect 18325 19428 18337 19431
rect 18104 19400 18337 19428
rect 18104 19388 18110 19400
rect 18325 19397 18337 19400
rect 18371 19397 18383 19431
rect 18325 19391 18383 19397
rect 18506 19388 18512 19440
rect 18564 19428 18570 19440
rect 18782 19428 18788 19440
rect 18564 19400 18788 19428
rect 18564 19388 18570 19400
rect 18782 19388 18788 19400
rect 18840 19388 18846 19440
rect 21542 19428 21548 19440
rect 21206 19400 21548 19428
rect 21542 19388 21548 19400
rect 21600 19428 21606 19440
rect 21818 19428 21824 19440
rect 21600 19400 21824 19428
rect 21600 19388 21606 19400
rect 21818 19388 21824 19400
rect 21876 19388 21882 19440
rect 22465 19431 22523 19437
rect 22465 19397 22477 19431
rect 22511 19428 22523 19431
rect 22646 19428 22652 19440
rect 22511 19400 22652 19428
rect 22511 19397 22523 19400
rect 22465 19391 22523 19397
rect 22646 19388 22652 19400
rect 22704 19388 22710 19440
rect 17552 19332 18000 19360
rect 17552 19320 17558 19332
rect 18138 19320 18144 19372
rect 18196 19360 18202 19372
rect 18233 19363 18291 19369
rect 18233 19360 18245 19363
rect 18196 19332 18245 19360
rect 18196 19320 18202 19332
rect 18233 19329 18245 19332
rect 18279 19329 18291 19363
rect 18233 19323 18291 19329
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19245 19363 19303 19369
rect 19245 19360 19257 19363
rect 19116 19332 19257 19360
rect 19116 19320 19122 19332
rect 19245 19329 19257 19332
rect 19291 19329 19303 19363
rect 19245 19323 19303 19329
rect 21910 19320 21916 19372
rect 21968 19360 21974 19372
rect 23952 19360 23980 19468
rect 25866 19456 25872 19468
rect 25924 19456 25930 19508
rect 26234 19456 26240 19508
rect 26292 19496 26298 19508
rect 26421 19499 26479 19505
rect 26421 19496 26433 19499
rect 26292 19468 26433 19496
rect 26292 19456 26298 19468
rect 26421 19465 26433 19468
rect 26467 19465 26479 19499
rect 26421 19459 26479 19465
rect 27154 19456 27160 19508
rect 27212 19496 27218 19508
rect 27709 19499 27767 19505
rect 27709 19496 27721 19499
rect 27212 19468 27721 19496
rect 27212 19456 27218 19468
rect 27709 19465 27721 19468
rect 27755 19465 27767 19499
rect 27709 19459 27767 19465
rect 30469 19499 30527 19505
rect 30469 19465 30481 19499
rect 30515 19496 30527 19499
rect 30515 19468 31754 19496
rect 30515 19465 30527 19468
rect 30469 19459 30527 19465
rect 24121 19431 24179 19437
rect 24121 19397 24133 19431
rect 24167 19428 24179 19431
rect 25498 19428 25504 19440
rect 24167 19400 25504 19428
rect 24167 19397 24179 19400
rect 24121 19391 24179 19397
rect 25498 19388 25504 19400
rect 25556 19388 25562 19440
rect 26602 19388 26608 19440
rect 26660 19428 26666 19440
rect 26970 19428 26976 19440
rect 26660 19400 26976 19428
rect 26660 19388 26666 19400
rect 26970 19388 26976 19400
rect 27028 19428 27034 19440
rect 27246 19428 27252 19440
rect 27028 19400 27252 19428
rect 27028 19388 27034 19400
rect 27246 19388 27252 19400
rect 27304 19388 27310 19440
rect 28537 19431 28595 19437
rect 28537 19397 28549 19431
rect 28583 19428 28595 19431
rect 28626 19428 28632 19440
rect 28583 19400 28632 19428
rect 28583 19397 28595 19400
rect 28537 19391 28595 19397
rect 28626 19388 28632 19400
rect 28684 19388 28690 19440
rect 31726 19428 31754 19468
rect 32030 19428 32036 19440
rect 31726 19400 32036 19428
rect 32030 19388 32036 19400
rect 32088 19388 32094 19440
rect 21968 19332 23980 19360
rect 24029 19363 24087 19369
rect 21968 19320 21974 19332
rect 24029 19329 24041 19363
rect 24075 19329 24087 19363
rect 24029 19323 24087 19329
rect 24949 19363 25007 19369
rect 24949 19329 24961 19363
rect 24995 19329 25007 19363
rect 24949 19323 25007 19329
rect 13449 19295 13507 19301
rect 13449 19261 13461 19295
rect 13495 19261 13507 19295
rect 13449 19255 13507 19261
rect 13909 19295 13967 19301
rect 13909 19261 13921 19295
rect 13955 19292 13967 19295
rect 14642 19292 14648 19304
rect 13955 19264 14648 19292
rect 13955 19261 13967 19264
rect 13909 19255 13967 19261
rect 14642 19252 14648 19264
rect 14700 19252 14706 19304
rect 14918 19252 14924 19304
rect 14976 19252 14982 19304
rect 15102 19252 15108 19304
rect 15160 19292 15166 19304
rect 15160 19264 15976 19292
rect 15160 19252 15166 19264
rect 5408 19196 6592 19224
rect 5408 19184 5414 19196
rect 6638 19184 6644 19236
rect 6696 19224 6702 19236
rect 8386 19224 8392 19236
rect 6696 19196 8392 19224
rect 6696 19184 6702 19196
rect 8386 19184 8392 19196
rect 8444 19224 8450 19236
rect 9490 19224 9496 19236
rect 8444 19196 9496 19224
rect 8444 19184 8450 19196
rect 9490 19184 9496 19196
rect 9548 19184 9554 19236
rect 10137 19227 10195 19233
rect 10137 19193 10149 19227
rect 10183 19224 10195 19227
rect 11698 19224 11704 19236
rect 10183 19196 11704 19224
rect 10183 19193 10195 19196
rect 10137 19187 10195 19193
rect 11698 19184 11704 19196
rect 11756 19184 11762 19236
rect 15841 19227 15899 19233
rect 15841 19224 15853 19227
rect 13096 19196 15853 19224
rect 4798 19116 4804 19168
rect 4856 19156 4862 19168
rect 6362 19156 6368 19168
rect 4856 19128 6368 19156
rect 4856 19116 4862 19128
rect 6362 19116 6368 19128
rect 6420 19116 6426 19168
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 13096 19156 13124 19196
rect 15841 19193 15853 19196
rect 15887 19193 15899 19227
rect 15948 19224 15976 19264
rect 16298 19252 16304 19304
rect 16356 19292 16362 19304
rect 16850 19292 16856 19304
rect 16356 19264 16856 19292
rect 16356 19252 16362 19264
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 16945 19295 17003 19301
rect 16945 19261 16957 19295
rect 16991 19292 17003 19295
rect 17586 19292 17592 19304
rect 16991 19264 17592 19292
rect 16991 19261 17003 19264
rect 16945 19255 17003 19261
rect 17586 19252 17592 19264
rect 17644 19252 17650 19304
rect 18046 19252 18052 19304
rect 18104 19292 18110 19304
rect 18417 19295 18475 19301
rect 18417 19292 18429 19295
rect 18104 19264 18429 19292
rect 18104 19252 18110 19264
rect 18417 19261 18429 19264
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 19702 19252 19708 19304
rect 19760 19252 19766 19304
rect 20622 19252 20628 19304
rect 20680 19292 20686 19304
rect 22646 19292 22652 19304
rect 20680 19264 22652 19292
rect 20680 19252 20686 19264
rect 22646 19252 22652 19264
rect 22704 19252 22710 19304
rect 23382 19252 23388 19304
rect 23440 19292 23446 19304
rect 24044 19292 24072 19323
rect 23440 19264 24072 19292
rect 24305 19295 24363 19301
rect 23440 19252 23446 19264
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 24854 19292 24860 19304
rect 24351 19264 24860 19292
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 16482 19224 16488 19236
rect 15948 19196 16488 19224
rect 15841 19187 15899 19193
rect 16482 19184 16488 19196
rect 16540 19184 16546 19236
rect 16868 19224 16896 19252
rect 19720 19224 19748 19252
rect 16868 19196 19748 19224
rect 21818 19184 21824 19236
rect 21876 19224 21882 19236
rect 21876 19196 22140 19224
rect 21876 19184 21882 19196
rect 11112 19128 13124 19156
rect 11112 19116 11118 19128
rect 13170 19116 13176 19168
rect 13228 19156 13234 19168
rect 14093 19159 14151 19165
rect 14093 19156 14105 19159
rect 13228 19128 14105 19156
rect 13228 19116 13234 19128
rect 14093 19125 14105 19128
rect 14139 19156 14151 19159
rect 14182 19156 14188 19168
rect 14139 19128 14188 19156
rect 14139 19125 14151 19128
rect 14093 19119 14151 19125
rect 14182 19116 14188 19128
rect 14240 19116 14246 19168
rect 14366 19116 14372 19168
rect 14424 19116 14430 19168
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 16022 19156 16028 19168
rect 14516 19128 16028 19156
rect 14516 19116 14522 19128
rect 16022 19116 16028 19128
rect 16080 19116 16086 19168
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 16209 19159 16267 19165
rect 16209 19156 16221 19159
rect 16172 19128 16221 19156
rect 16172 19116 16178 19128
rect 16209 19125 16221 19128
rect 16255 19125 16267 19159
rect 16209 19119 16267 19125
rect 16393 19159 16451 19165
rect 16393 19125 16405 19159
rect 16439 19156 16451 19159
rect 16574 19156 16580 19168
rect 16439 19128 16580 19156
rect 16439 19125 16451 19128
rect 16393 19119 16451 19125
rect 16574 19116 16580 19128
rect 16632 19116 16638 19168
rect 16761 19159 16819 19165
rect 16761 19125 16773 19159
rect 16807 19156 16819 19159
rect 16850 19156 16856 19168
rect 16807 19128 16856 19156
rect 16807 19125 16819 19128
rect 16761 19119 16819 19125
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 17402 19116 17408 19168
rect 17460 19156 17466 19168
rect 17681 19159 17739 19165
rect 17681 19156 17693 19159
rect 17460 19128 17693 19156
rect 17460 19116 17466 19128
rect 17681 19125 17693 19128
rect 17727 19156 17739 19159
rect 18138 19156 18144 19168
rect 17727 19128 18144 19156
rect 17727 19125 17739 19128
rect 17681 19119 17739 19125
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 18874 19116 18880 19168
rect 18932 19156 18938 19168
rect 19968 19159 20026 19165
rect 19968 19156 19980 19159
rect 18932 19128 19980 19156
rect 18932 19116 18938 19128
rect 19968 19125 19980 19128
rect 20014 19156 20026 19159
rect 20990 19156 20996 19168
rect 20014 19128 20996 19156
rect 20014 19125 20026 19128
rect 19968 19119 20026 19125
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 22002 19116 22008 19168
rect 22060 19116 22066 19168
rect 22112 19156 22140 19196
rect 22186 19184 22192 19236
rect 22244 19224 22250 19236
rect 23293 19227 23351 19233
rect 23293 19224 23305 19227
rect 22244 19196 23305 19224
rect 22244 19184 22250 19196
rect 23293 19193 23305 19196
rect 23339 19224 23351 19227
rect 24964 19224 24992 19323
rect 29638 19320 29644 19372
rect 29696 19320 29702 19372
rect 30650 19320 30656 19372
rect 30708 19360 30714 19372
rect 31113 19363 31171 19369
rect 31113 19360 31125 19363
rect 30708 19332 31125 19360
rect 30708 19320 30714 19332
rect 31113 19329 31125 19332
rect 31159 19329 31171 19363
rect 31113 19323 31171 19329
rect 25774 19252 25780 19304
rect 25832 19252 25838 19304
rect 26878 19252 26884 19304
rect 26936 19292 26942 19304
rect 26973 19295 27031 19301
rect 26973 19292 26985 19295
rect 26936 19264 26985 19292
rect 26936 19252 26942 19264
rect 26973 19261 26985 19264
rect 27019 19261 27031 19295
rect 26973 19255 27031 19261
rect 27798 19252 27804 19304
rect 27856 19292 27862 19304
rect 28261 19295 28319 19301
rect 28261 19292 28273 19295
rect 27856 19264 28273 19292
rect 27856 19252 27862 19264
rect 28261 19261 28273 19264
rect 28307 19261 28319 19295
rect 29656 19292 29684 19320
rect 30834 19292 30840 19304
rect 29656 19264 30840 19292
rect 28261 19255 28319 19261
rect 30834 19252 30840 19264
rect 30892 19292 30898 19304
rect 30929 19295 30987 19301
rect 30929 19292 30941 19295
rect 30892 19264 30941 19292
rect 30892 19252 30898 19264
rect 30929 19261 30941 19264
rect 30975 19261 30987 19295
rect 30929 19255 30987 19261
rect 25314 19224 25320 19236
rect 23339 19196 25320 19224
rect 23339 19193 23351 19196
rect 23293 19187 23351 19193
rect 25314 19184 25320 19196
rect 25372 19184 25378 19236
rect 27430 19184 27436 19236
rect 27488 19184 27494 19236
rect 22554 19156 22560 19168
rect 22112 19128 22560 19156
rect 22554 19116 22560 19128
rect 22612 19156 22618 19168
rect 23109 19159 23167 19165
rect 23109 19156 23121 19159
rect 22612 19128 23121 19156
rect 22612 19116 22618 19128
rect 23109 19125 23121 19128
rect 23155 19156 23167 19159
rect 23750 19156 23756 19168
rect 23155 19128 23756 19156
rect 23155 19125 23167 19128
rect 23109 19119 23167 19125
rect 23750 19116 23756 19128
rect 23808 19116 23814 19168
rect 25222 19116 25228 19168
rect 25280 19156 25286 19168
rect 26602 19156 26608 19168
rect 25280 19128 26608 19156
rect 25280 19116 25286 19128
rect 26602 19116 26608 19128
rect 26660 19116 26666 19168
rect 27614 19116 27620 19168
rect 27672 19156 27678 19168
rect 27893 19159 27951 19165
rect 27893 19156 27905 19159
rect 27672 19128 27905 19156
rect 27672 19116 27678 19128
rect 27893 19125 27905 19128
rect 27939 19156 27951 19159
rect 28350 19156 28356 19168
rect 27939 19128 28356 19156
rect 27939 19125 27951 19128
rect 27893 19119 27951 19125
rect 28350 19116 28356 19128
rect 28408 19116 28414 19168
rect 28626 19116 28632 19168
rect 28684 19156 28690 19168
rect 30009 19159 30067 19165
rect 30009 19156 30021 19159
rect 28684 19128 30021 19156
rect 28684 19116 28690 19128
rect 30009 19125 30021 19128
rect 30055 19156 30067 19159
rect 30282 19156 30288 19168
rect 30055 19128 30288 19156
rect 30055 19125 30067 19128
rect 30009 19119 30067 19125
rect 30282 19116 30288 19128
rect 30340 19116 30346 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 3927 18924 8156 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 3988 18825 4016 18924
rect 8128 18884 8156 18924
rect 9398 18912 9404 18964
rect 9456 18912 9462 18964
rect 9766 18912 9772 18964
rect 9824 18952 9830 18964
rect 11609 18955 11667 18961
rect 11609 18952 11621 18955
rect 9824 18924 11621 18952
rect 9824 18912 9830 18924
rect 11609 18921 11621 18924
rect 11655 18921 11667 18955
rect 11609 18915 11667 18921
rect 12250 18912 12256 18964
rect 12308 18952 12314 18964
rect 14366 18952 14372 18964
rect 12308 18924 14372 18952
rect 12308 18912 12314 18924
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 14826 18912 14832 18964
rect 14884 18952 14890 18964
rect 22002 18952 22008 18964
rect 14884 18924 22008 18952
rect 14884 18912 14890 18924
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 22646 18912 22652 18964
rect 22704 18952 22710 18964
rect 22925 18955 22983 18961
rect 22925 18952 22937 18955
rect 22704 18924 22937 18952
rect 22704 18912 22710 18924
rect 22925 18921 22937 18924
rect 22971 18921 22983 18955
rect 25682 18952 25688 18964
rect 22925 18915 22983 18921
rect 25516 18924 25688 18952
rect 14185 18887 14243 18893
rect 8128 18856 14136 18884
rect 3973 18819 4031 18825
rect 3973 18785 3985 18819
rect 4019 18785 4031 18819
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 3973 18779 4031 18785
rect 4632 18788 6837 18816
rect 4632 18760 4660 18788
rect 6825 18785 6837 18788
rect 6871 18816 6883 18819
rect 8478 18816 8484 18828
rect 6871 18788 8484 18816
rect 6871 18785 6883 18788
rect 6825 18779 6883 18785
rect 8478 18776 8484 18788
rect 8536 18776 8542 18828
rect 8573 18819 8631 18825
rect 8573 18785 8585 18819
rect 8619 18785 8631 18819
rect 8573 18779 8631 18785
rect 9033 18819 9091 18825
rect 9033 18785 9045 18819
rect 9079 18816 9091 18819
rect 9306 18816 9312 18828
rect 9079 18788 9312 18816
rect 9079 18785 9091 18788
rect 9033 18779 9091 18785
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18748 1823 18751
rect 4430 18748 4436 18760
rect 1811 18720 4436 18748
rect 1811 18717 1823 18720
rect 1765 18711 1823 18717
rect 4430 18708 4436 18720
rect 4488 18708 4494 18760
rect 4614 18708 4620 18760
rect 4672 18708 4678 18760
rect 8588 18748 8616 18779
rect 9306 18776 9312 18788
rect 9364 18776 9370 18828
rect 9766 18776 9772 18828
rect 9824 18816 9830 18828
rect 9861 18819 9919 18825
rect 9861 18816 9873 18819
rect 9824 18788 9873 18816
rect 9824 18776 9830 18788
rect 9861 18785 9873 18788
rect 9907 18785 9919 18819
rect 9861 18779 9919 18785
rect 9950 18776 9956 18828
rect 10008 18776 10014 18828
rect 10226 18776 10232 18828
rect 10284 18816 10290 18828
rect 10962 18816 10968 18828
rect 10284 18788 10968 18816
rect 10284 18776 10290 18788
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 11146 18776 11152 18828
rect 11204 18816 11210 18828
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 11204 18788 12173 18816
rect 11204 18776 11210 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 14108 18816 14136 18856
rect 14185 18853 14197 18887
rect 14231 18884 14243 18887
rect 14458 18884 14464 18896
rect 14231 18856 14464 18884
rect 14231 18853 14243 18856
rect 14185 18847 14243 18853
rect 14458 18844 14464 18856
rect 14516 18844 14522 18896
rect 16482 18844 16488 18896
rect 16540 18884 16546 18896
rect 18141 18887 18199 18893
rect 16540 18856 17632 18884
rect 16540 18844 16546 18856
rect 15102 18816 15108 18828
rect 14108 18788 15108 18816
rect 12161 18779 12219 18785
rect 15102 18776 15108 18788
rect 15160 18776 15166 18828
rect 15197 18819 15255 18825
rect 15197 18785 15209 18819
rect 15243 18816 15255 18819
rect 16206 18816 16212 18828
rect 15243 18788 16212 18816
rect 15243 18785 15255 18788
rect 15197 18779 15255 18785
rect 16206 18776 16212 18788
rect 16264 18776 16270 18828
rect 16666 18776 16672 18828
rect 16724 18816 16730 18828
rect 17497 18819 17555 18825
rect 17497 18816 17509 18819
rect 16724 18788 17509 18816
rect 16724 18776 16730 18788
rect 17497 18785 17509 18788
rect 17543 18785 17555 18819
rect 17604 18816 17632 18856
rect 18141 18853 18153 18887
rect 18187 18884 18199 18887
rect 18322 18884 18328 18896
rect 18187 18856 18328 18884
rect 18187 18853 18199 18856
rect 18141 18847 18199 18853
rect 18322 18844 18328 18856
rect 18380 18844 18386 18896
rect 19334 18844 19340 18896
rect 19392 18884 19398 18896
rect 20714 18884 20720 18896
rect 19392 18856 20720 18884
rect 19392 18844 19398 18856
rect 20714 18844 20720 18856
rect 20772 18844 20778 18896
rect 25130 18844 25136 18896
rect 25188 18884 25194 18896
rect 25516 18884 25544 18924
rect 25682 18912 25688 18924
rect 25740 18912 25746 18964
rect 26142 18912 26148 18964
rect 26200 18952 26206 18964
rect 27157 18955 27215 18961
rect 27157 18952 27169 18955
rect 26200 18924 27169 18952
rect 26200 18912 26206 18924
rect 27157 18921 27169 18924
rect 27203 18921 27215 18955
rect 27157 18915 27215 18921
rect 27246 18912 27252 18964
rect 27304 18952 27310 18964
rect 47026 18952 47032 18964
rect 27304 18924 47032 18952
rect 27304 18912 27310 18924
rect 47026 18912 47032 18924
rect 47084 18912 47090 18964
rect 25188 18856 25544 18884
rect 25188 18844 25194 18856
rect 26786 18844 26792 18896
rect 26844 18884 26850 18896
rect 26844 18856 31754 18884
rect 26844 18844 26850 18856
rect 18693 18819 18751 18825
rect 18693 18816 18705 18819
rect 17604 18788 18705 18816
rect 17497 18779 17555 18785
rect 18693 18785 18705 18788
rect 18739 18785 18751 18819
rect 18693 18779 18751 18785
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 20349 18819 20407 18825
rect 20349 18816 20361 18819
rect 19760 18788 20361 18816
rect 19760 18776 19766 18788
rect 20349 18785 20361 18788
rect 20395 18816 20407 18819
rect 21177 18819 21235 18825
rect 21177 18816 21189 18819
rect 20395 18788 21189 18816
rect 20395 18785 20407 18788
rect 20349 18779 20407 18785
rect 21177 18785 21189 18788
rect 21223 18785 21235 18819
rect 21177 18779 21235 18785
rect 21450 18776 21456 18828
rect 21508 18776 21514 18828
rect 21542 18776 21548 18828
rect 21600 18816 21606 18828
rect 21600 18788 23520 18816
rect 21600 18776 21606 18788
rect 9122 18748 9128 18760
rect 8588 18720 9128 18748
rect 9122 18708 9128 18720
rect 9180 18748 9186 18760
rect 10042 18748 10048 18760
rect 9180 18720 10048 18748
rect 9180 18708 9186 18720
rect 10042 18708 10048 18720
rect 10100 18708 10106 18760
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18748 10655 18751
rect 11330 18748 11336 18760
rect 10643 18720 11336 18748
rect 10643 18717 10655 18720
rect 10597 18711 10655 18717
rect 11330 18708 11336 18720
rect 11388 18708 11394 18760
rect 11882 18708 11888 18760
rect 11940 18748 11946 18760
rect 13354 18748 13360 18760
rect 11940 18720 13360 18748
rect 11940 18708 11946 18720
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18748 14611 18751
rect 14826 18748 14832 18760
rect 14599 18720 14832 18748
rect 14599 18717 14611 18720
rect 14553 18711 14611 18717
rect 14826 18708 14832 18720
rect 14884 18708 14890 18760
rect 17034 18708 17040 18760
rect 17092 18748 17098 18760
rect 18046 18748 18052 18760
rect 17092 18720 18052 18748
rect 17092 18708 17098 18720
rect 18046 18708 18052 18720
rect 18104 18708 18110 18760
rect 18598 18708 18604 18760
rect 18656 18748 18662 18760
rect 18874 18748 18880 18760
rect 18656 18720 18880 18748
rect 18656 18708 18662 18720
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 19659 18720 20944 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 2774 18640 2780 18692
rect 2832 18640 2838 18692
rect 3050 18640 3056 18692
rect 3108 18680 3114 18692
rect 3605 18683 3663 18689
rect 3605 18680 3617 18683
rect 3108 18652 3617 18680
rect 3108 18640 3114 18652
rect 3605 18649 3617 18652
rect 3651 18680 3663 18683
rect 4062 18680 4068 18692
rect 3651 18652 4068 18680
rect 3651 18649 3663 18652
rect 3605 18643 3663 18649
rect 4062 18640 4068 18652
rect 4120 18640 4126 18692
rect 4798 18640 4804 18692
rect 4856 18680 4862 18692
rect 4893 18683 4951 18689
rect 4893 18680 4905 18683
rect 4856 18652 4905 18680
rect 4856 18640 4862 18652
rect 4893 18649 4905 18652
rect 4939 18649 4951 18683
rect 4893 18643 4951 18649
rect 3326 18572 3332 18624
rect 3384 18572 3390 18624
rect 4908 18612 4936 18643
rect 5442 18640 5448 18692
rect 5500 18640 5506 18692
rect 7101 18683 7159 18689
rect 7101 18649 7113 18683
rect 7147 18680 7159 18683
rect 7190 18680 7196 18692
rect 7147 18652 7196 18680
rect 7147 18649 7159 18652
rect 7101 18643 7159 18649
rect 7190 18640 7196 18652
rect 7248 18640 7254 18692
rect 7558 18640 7564 18692
rect 7616 18640 7622 18692
rect 8570 18640 8576 18692
rect 8628 18680 8634 18692
rect 8628 18652 8892 18680
rect 8628 18640 8634 18652
rect 6178 18612 6184 18624
rect 4908 18584 6184 18612
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 6362 18572 6368 18624
rect 6420 18612 6426 18624
rect 8754 18612 8760 18624
rect 6420 18584 8760 18612
rect 6420 18572 6426 18584
rect 8754 18572 8760 18584
rect 8812 18572 8818 18624
rect 8864 18612 8892 18652
rect 8938 18640 8944 18692
rect 8996 18680 9002 18692
rect 8996 18652 10640 18680
rect 8996 18640 9002 18652
rect 9769 18615 9827 18621
rect 9769 18612 9781 18615
rect 8864 18584 9781 18612
rect 9769 18581 9781 18584
rect 9815 18612 9827 18615
rect 9858 18612 9864 18624
rect 9815 18584 9864 18612
rect 9815 18581 9827 18584
rect 9769 18575 9827 18581
rect 9858 18572 9864 18584
rect 9916 18572 9922 18624
rect 10612 18612 10640 18652
rect 10686 18640 10692 18692
rect 10744 18680 10750 18692
rect 10965 18683 11023 18689
rect 10965 18680 10977 18683
rect 10744 18652 10977 18680
rect 10744 18640 10750 18652
rect 10965 18649 10977 18652
rect 11011 18680 11023 18683
rect 12805 18683 12863 18689
rect 11011 18652 12434 18680
rect 11011 18649 11023 18652
rect 10965 18643 11023 18649
rect 11057 18615 11115 18621
rect 11057 18612 11069 18615
rect 10612 18584 11069 18612
rect 11057 18581 11069 18584
rect 11103 18581 11115 18615
rect 11057 18575 11115 18581
rect 11330 18572 11336 18624
rect 11388 18612 11394 18624
rect 11606 18612 11612 18624
rect 11388 18584 11612 18612
rect 11388 18572 11394 18584
rect 11606 18572 11612 18584
rect 11664 18612 11670 18624
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 11664 18584 11989 18612
rect 11664 18572 11670 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 11977 18575 12035 18581
rect 12066 18572 12072 18624
rect 12124 18572 12130 18624
rect 12406 18612 12434 18652
rect 12805 18649 12817 18683
rect 12851 18680 12863 18683
rect 13170 18680 13176 18692
rect 12851 18652 13176 18680
rect 12851 18649 12863 18652
rect 12805 18643 12863 18649
rect 13170 18640 13176 18652
rect 13228 18640 13234 18692
rect 13538 18640 13544 18692
rect 13596 18640 13602 18692
rect 15473 18683 15531 18689
rect 13648 18652 13860 18680
rect 13648 18612 13676 18652
rect 12406 18584 13676 18612
rect 13832 18612 13860 18652
rect 15473 18649 15485 18683
rect 15519 18649 15531 18683
rect 15473 18643 15531 18649
rect 14645 18615 14703 18621
rect 14645 18612 14657 18615
rect 13832 18584 14657 18612
rect 14645 18581 14657 18584
rect 14691 18581 14703 18615
rect 14645 18575 14703 18581
rect 15286 18572 15292 18624
rect 15344 18612 15350 18624
rect 15488 18612 15516 18643
rect 16022 18640 16028 18692
rect 16080 18640 16086 18692
rect 20070 18680 20076 18692
rect 16776 18652 20076 18680
rect 16390 18612 16396 18624
rect 15344 18584 16396 18612
rect 15344 18572 15350 18584
rect 16390 18572 16396 18584
rect 16448 18612 16454 18624
rect 16776 18612 16804 18652
rect 20070 18640 20076 18652
rect 20128 18640 20134 18692
rect 16448 18584 16804 18612
rect 16448 18572 16454 18584
rect 16942 18572 16948 18624
rect 17000 18572 17006 18624
rect 17586 18572 17592 18624
rect 17644 18612 17650 18624
rect 18509 18615 18567 18621
rect 18509 18612 18521 18615
rect 17644 18584 18521 18612
rect 17644 18572 17650 18584
rect 18509 18581 18521 18584
rect 18555 18612 18567 18615
rect 18598 18612 18604 18624
rect 18555 18584 18604 18612
rect 18555 18581 18567 18584
rect 18509 18575 18567 18581
rect 18598 18572 18604 18584
rect 18656 18572 18662 18624
rect 19337 18615 19395 18621
rect 19337 18581 19349 18615
rect 19383 18612 19395 18615
rect 19518 18612 19524 18624
rect 19383 18584 19524 18612
rect 19383 18581 19395 18584
rect 19337 18575 19395 18581
rect 19518 18572 19524 18584
rect 19576 18612 19582 18624
rect 19794 18612 19800 18624
rect 19576 18584 19800 18612
rect 19576 18572 19582 18584
rect 19794 18572 19800 18584
rect 19852 18572 19858 18624
rect 20806 18572 20812 18624
rect 20864 18572 20870 18624
rect 20916 18612 20944 18720
rect 22554 18708 22560 18760
rect 22612 18708 22618 18760
rect 23492 18680 23520 18788
rect 23658 18776 23664 18828
rect 23716 18816 23722 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 23716 18788 24593 18816
rect 23716 18776 23722 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 25409 18819 25467 18825
rect 25409 18785 25421 18819
rect 25455 18816 25467 18819
rect 25774 18816 25780 18828
rect 25455 18788 25780 18816
rect 25455 18785 25467 18788
rect 25409 18779 25467 18785
rect 25774 18776 25780 18788
rect 25832 18776 25838 18828
rect 26234 18776 26240 18828
rect 26292 18816 26298 18828
rect 27617 18819 27675 18825
rect 27617 18816 27629 18819
rect 26292 18788 27629 18816
rect 26292 18776 26298 18788
rect 27617 18785 27629 18788
rect 27663 18785 27675 18819
rect 27617 18779 27675 18785
rect 30190 18776 30196 18828
rect 30248 18776 30254 18828
rect 30285 18819 30343 18825
rect 30285 18785 30297 18819
rect 30331 18785 30343 18819
rect 30285 18779 30343 18785
rect 23566 18708 23572 18760
rect 23624 18708 23630 18760
rect 23750 18708 23756 18760
rect 23808 18748 23814 18760
rect 24029 18751 24087 18757
rect 24029 18748 24041 18751
rect 23808 18720 24041 18748
rect 23808 18708 23814 18720
rect 24029 18717 24041 18720
rect 24075 18748 24087 18751
rect 25130 18748 25136 18760
rect 24075 18720 25136 18748
rect 24075 18717 24087 18720
rect 24029 18711 24087 18717
rect 25130 18708 25136 18720
rect 25188 18708 25194 18760
rect 27706 18708 27712 18760
rect 27764 18748 27770 18760
rect 27893 18751 27951 18757
rect 27893 18748 27905 18751
rect 27764 18720 27905 18748
rect 27764 18708 27770 18720
rect 27893 18717 27905 18720
rect 27939 18717 27951 18751
rect 27893 18711 27951 18717
rect 29822 18708 29828 18760
rect 29880 18748 29886 18760
rect 30300 18748 30328 18779
rect 30834 18776 30840 18828
rect 30892 18776 30898 18828
rect 31726 18816 31754 18856
rect 46934 18816 46940 18828
rect 31726 18788 46940 18816
rect 46934 18776 46940 18788
rect 46992 18776 46998 18828
rect 29880 18720 30328 18748
rect 29880 18708 29886 18720
rect 25685 18683 25743 18689
rect 23492 18652 25636 18680
rect 22094 18612 22100 18624
rect 20916 18584 22100 18612
rect 22094 18572 22100 18584
rect 22152 18572 22158 18624
rect 23382 18572 23388 18624
rect 23440 18572 23446 18624
rect 23474 18572 23480 18624
rect 23532 18612 23538 18624
rect 23842 18612 23848 18624
rect 23532 18584 23848 18612
rect 23532 18572 23538 18584
rect 23842 18572 23848 18584
rect 23900 18612 23906 18624
rect 24121 18615 24179 18621
rect 24121 18612 24133 18615
rect 23900 18584 24133 18612
rect 23900 18572 23906 18584
rect 24121 18581 24133 18584
rect 24167 18581 24179 18615
rect 25608 18612 25636 18652
rect 25685 18649 25697 18683
rect 25731 18680 25743 18683
rect 25958 18680 25964 18692
rect 25731 18652 25964 18680
rect 25731 18649 25743 18652
rect 25685 18643 25743 18649
rect 25958 18640 25964 18652
rect 26016 18640 26022 18692
rect 26970 18680 26976 18692
rect 26910 18652 26976 18680
rect 26970 18640 26976 18652
rect 27028 18640 27034 18692
rect 30650 18680 30656 18692
rect 27080 18652 30656 18680
rect 27080 18612 27108 18652
rect 30650 18640 30656 18652
rect 30708 18640 30714 18692
rect 25608 18584 27108 18612
rect 24121 18575 24179 18581
rect 29730 18572 29736 18624
rect 29788 18572 29794 18624
rect 30098 18572 30104 18624
rect 30156 18572 30162 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 5626 18408 5632 18420
rect 2746 18380 5632 18408
rect 2746 18340 2774 18380
rect 5626 18368 5632 18380
rect 5684 18368 5690 18420
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 8938 18408 8944 18420
rect 6972 18380 8944 18408
rect 6972 18368 6978 18380
rect 8938 18368 8944 18380
rect 8996 18368 9002 18420
rect 9769 18411 9827 18417
rect 9769 18377 9781 18411
rect 9815 18408 9827 18411
rect 10226 18408 10232 18420
rect 9815 18380 10232 18408
rect 9815 18377 9827 18380
rect 9769 18371 9827 18377
rect 10226 18368 10232 18380
rect 10284 18368 10290 18420
rect 10413 18411 10471 18417
rect 10413 18377 10425 18411
rect 10459 18408 10471 18411
rect 11882 18408 11888 18420
rect 10459 18380 11888 18408
rect 10459 18377 10471 18380
rect 10413 18371 10471 18377
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 12345 18411 12403 18417
rect 12345 18408 12357 18411
rect 12084 18380 12357 18408
rect 5902 18340 5908 18352
rect 1780 18312 2774 18340
rect 3620 18312 5908 18340
rect 1780 18281 1808 18312
rect 3620 18281 3648 18312
rect 5902 18300 5908 18312
rect 5960 18300 5966 18352
rect 7466 18300 7472 18352
rect 7524 18340 7530 18352
rect 9582 18340 9588 18352
rect 7524 18312 9588 18340
rect 7524 18300 7530 18312
rect 9582 18300 9588 18312
rect 9640 18300 9646 18352
rect 9953 18343 10011 18349
rect 9953 18309 9965 18343
rect 9999 18340 10011 18343
rect 10502 18340 10508 18352
rect 9999 18312 10508 18340
rect 9999 18309 10011 18312
rect 9953 18303 10011 18309
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18241 1823 18275
rect 1765 18235 1823 18241
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 5626 18232 5632 18284
rect 5684 18232 5690 18284
rect 5721 18275 5779 18281
rect 5721 18241 5733 18275
rect 5767 18272 5779 18275
rect 6086 18272 6092 18284
rect 5767 18244 6092 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 6086 18232 6092 18244
rect 6144 18272 6150 18284
rect 6638 18272 6644 18284
rect 6144 18244 6644 18272
rect 6144 18232 6150 18244
rect 6638 18232 6644 18244
rect 6696 18232 6702 18284
rect 6730 18232 6736 18284
rect 6788 18232 6794 18284
rect 7006 18232 7012 18284
rect 7064 18272 7070 18284
rect 7926 18272 7932 18284
rect 7064 18244 7932 18272
rect 7064 18232 7070 18244
rect 7926 18232 7932 18244
rect 7984 18232 7990 18284
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 8481 18275 8539 18281
rect 8481 18272 8493 18275
rect 8444 18244 8493 18272
rect 8444 18232 8450 18244
rect 8481 18241 8493 18244
rect 8527 18272 8539 18275
rect 9968 18272 9996 18303
rect 10502 18300 10508 18312
rect 10560 18300 10566 18352
rect 8527 18244 9996 18272
rect 8527 18241 8539 18244
rect 8481 18235 8539 18241
rect 10226 18232 10232 18284
rect 10284 18272 10290 18284
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 10284 18244 10793 18272
rect 10284 18232 10290 18244
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 11330 18232 11336 18284
rect 11388 18272 11394 18284
rect 12084 18272 12112 18380
rect 12345 18377 12357 18380
rect 12391 18377 12403 18411
rect 12345 18371 12403 18377
rect 12452 18380 12756 18408
rect 12452 18340 12480 18380
rect 11388 18244 12112 18272
rect 12268 18312 12480 18340
rect 12728 18340 12756 18380
rect 13722 18368 13728 18420
rect 13780 18408 13786 18420
rect 15381 18411 15439 18417
rect 15381 18408 15393 18411
rect 13780 18380 15393 18408
rect 13780 18368 13786 18380
rect 15381 18377 15393 18380
rect 15427 18377 15439 18411
rect 15381 18371 15439 18377
rect 17313 18411 17371 18417
rect 17313 18377 17325 18411
rect 17359 18408 17371 18411
rect 19334 18408 19340 18420
rect 17359 18380 19340 18408
rect 17359 18377 17371 18380
rect 17313 18371 17371 18377
rect 19334 18368 19340 18380
rect 19392 18368 19398 18420
rect 19889 18411 19947 18417
rect 19889 18408 19901 18411
rect 19812 18380 19901 18408
rect 19812 18352 19840 18380
rect 19889 18377 19901 18380
rect 19935 18377 19947 18411
rect 19889 18371 19947 18377
rect 20714 18368 20720 18420
rect 20772 18368 20778 18420
rect 20990 18368 20996 18420
rect 21048 18408 21054 18420
rect 24857 18411 24915 18417
rect 24857 18408 24869 18411
rect 21048 18380 24869 18408
rect 21048 18368 21054 18380
rect 24857 18377 24869 18380
rect 24903 18377 24915 18411
rect 24857 18371 24915 18377
rect 26789 18411 26847 18417
rect 26789 18377 26801 18411
rect 26835 18408 26847 18411
rect 26970 18408 26976 18420
rect 26835 18380 26976 18408
rect 26835 18377 26847 18380
rect 26789 18371 26847 18377
rect 26970 18368 26976 18380
rect 27028 18368 27034 18420
rect 27157 18411 27215 18417
rect 27157 18377 27169 18411
rect 27203 18408 27215 18411
rect 30098 18408 30104 18420
rect 27203 18380 30104 18408
rect 27203 18377 27215 18380
rect 27157 18371 27215 18377
rect 30098 18368 30104 18380
rect 30156 18368 30162 18420
rect 30650 18368 30656 18420
rect 30708 18408 30714 18420
rect 30745 18411 30803 18417
rect 30745 18408 30757 18411
rect 30708 18380 30757 18408
rect 30708 18368 30714 18380
rect 30745 18377 30757 18380
rect 30791 18408 30803 18411
rect 31481 18411 31539 18417
rect 31481 18408 31493 18411
rect 30791 18380 31493 18408
rect 30791 18377 30803 18380
rect 30745 18371 30803 18377
rect 31481 18377 31493 18380
rect 31527 18408 31539 18411
rect 38562 18408 38568 18420
rect 31527 18380 38568 18408
rect 31527 18377 31539 18380
rect 31481 18371 31539 18377
rect 38562 18368 38568 18380
rect 38620 18368 38626 18420
rect 13998 18340 14004 18352
rect 12728 18312 14004 18340
rect 11388 18232 11394 18244
rect 2038 18164 2044 18216
rect 2096 18164 2102 18216
rect 3786 18164 3792 18216
rect 3844 18204 3850 18216
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 3844 18176 3893 18204
rect 3844 18164 3850 18176
rect 3881 18173 3893 18176
rect 3927 18173 3939 18207
rect 3881 18167 3939 18173
rect 5902 18164 5908 18216
rect 5960 18164 5966 18216
rect 7282 18164 7288 18216
rect 7340 18164 7346 18216
rect 8570 18164 8576 18216
rect 8628 18204 8634 18216
rect 9217 18207 9275 18213
rect 9217 18204 9229 18207
rect 8628 18176 9229 18204
rect 8628 18164 8634 18176
rect 9217 18173 9229 18176
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 9490 18164 9496 18216
rect 9548 18204 9554 18216
rect 10873 18207 10931 18213
rect 10873 18204 10885 18207
rect 9548 18176 10885 18204
rect 9548 18164 9554 18176
rect 10873 18173 10885 18176
rect 10919 18173 10931 18207
rect 10873 18167 10931 18173
rect 11057 18207 11115 18213
rect 11057 18173 11069 18207
rect 11103 18204 11115 18207
rect 12268 18204 12296 18312
rect 13998 18300 14004 18312
rect 14056 18300 14062 18352
rect 14461 18343 14519 18349
rect 14461 18309 14473 18343
rect 14507 18340 14519 18343
rect 14550 18340 14556 18352
rect 14507 18312 14556 18340
rect 14507 18309 14519 18312
rect 14461 18303 14519 18309
rect 14550 18300 14556 18312
rect 14608 18300 14614 18352
rect 16022 18300 16028 18352
rect 16080 18340 16086 18352
rect 16209 18343 16267 18349
rect 16209 18340 16221 18343
rect 16080 18312 16221 18340
rect 16080 18300 16086 18312
rect 16209 18309 16221 18312
rect 16255 18309 16267 18343
rect 18141 18343 18199 18349
rect 16209 18303 16267 18309
rect 16408 18312 17356 18340
rect 12437 18275 12495 18281
rect 12437 18272 12449 18275
rect 11103 18176 12296 18204
rect 12360 18244 12449 18272
rect 11103 18173 11115 18176
rect 11057 18167 11115 18173
rect 6270 18096 6276 18148
rect 6328 18136 6334 18148
rect 7006 18136 7012 18148
rect 6328 18108 7012 18136
rect 6328 18096 6334 18108
rect 7006 18096 7012 18108
rect 7064 18096 7070 18148
rect 7926 18096 7932 18148
rect 7984 18136 7990 18148
rect 10686 18136 10692 18148
rect 7984 18108 10692 18136
rect 7984 18096 7990 18108
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 11882 18096 11888 18148
rect 11940 18136 11946 18148
rect 11977 18139 12035 18145
rect 11977 18136 11989 18139
rect 11940 18108 11989 18136
rect 11940 18096 11946 18108
rect 11977 18105 11989 18108
rect 12023 18105 12035 18139
rect 11977 18099 12035 18105
rect 1118 18068 1124 18080
rect 1044 18040 1124 18068
rect 1044 17728 1072 18040
rect 1118 18028 1124 18040
rect 1176 18028 1182 18080
rect 5261 18071 5319 18077
rect 5261 18037 5273 18071
rect 5307 18068 5319 18071
rect 6730 18068 6736 18080
rect 5307 18040 6736 18068
rect 5307 18037 5319 18040
rect 5261 18031 5319 18037
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 10045 18071 10103 18077
rect 10045 18068 10057 18071
rect 9916 18040 10057 18068
rect 9916 18028 9922 18040
rect 10045 18037 10057 18040
rect 10091 18068 10103 18071
rect 10134 18068 10140 18080
rect 10091 18040 10140 18068
rect 10091 18037 10103 18040
rect 10045 18031 10103 18037
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 11701 18071 11759 18077
rect 11701 18037 11713 18071
rect 11747 18068 11759 18071
rect 12066 18068 12072 18080
rect 11747 18040 12072 18068
rect 11747 18037 11759 18040
rect 11701 18031 11759 18037
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 12360 18068 12388 18244
rect 12437 18241 12449 18244
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 13633 18275 13691 18281
rect 13633 18241 13645 18275
rect 13679 18272 13691 18275
rect 13679 18244 13713 18272
rect 13679 18241 13691 18244
rect 13633 18235 13691 18241
rect 12621 18207 12679 18213
rect 12621 18173 12633 18207
rect 12667 18204 12679 18207
rect 12667 18176 12848 18204
rect 12667 18173 12679 18176
rect 12621 18167 12679 18173
rect 12820 18148 12848 18176
rect 13170 18164 13176 18216
rect 13228 18204 13234 18216
rect 13648 18204 13676 18235
rect 15194 18232 15200 18284
rect 15252 18272 15258 18284
rect 16408 18272 16436 18312
rect 15252 18244 16436 18272
rect 15252 18232 15258 18244
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 16632 18244 17233 18272
rect 16632 18232 16638 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17328 18272 17356 18312
rect 18141 18309 18153 18343
rect 18187 18340 18199 18343
rect 19702 18340 19708 18352
rect 18187 18312 19708 18340
rect 18187 18309 18199 18312
rect 18141 18303 18199 18309
rect 19702 18300 19708 18312
rect 19760 18300 19766 18352
rect 19794 18300 19800 18352
rect 19852 18300 19858 18352
rect 21082 18300 21088 18352
rect 21140 18300 21146 18352
rect 23474 18340 23480 18352
rect 21928 18312 23480 18340
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 17328 18244 18337 18272
rect 17221 18235 17279 18241
rect 18325 18241 18337 18244
rect 18371 18241 18383 18275
rect 19981 18275 20039 18281
rect 18325 18235 18383 18241
rect 18432 18244 19748 18272
rect 15102 18204 15108 18216
rect 13228 18176 15108 18204
rect 13228 18164 13234 18176
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 15473 18207 15531 18213
rect 15473 18173 15485 18207
rect 15519 18173 15531 18207
rect 15473 18167 15531 18173
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 16942 18204 16948 18216
rect 15703 18176 16948 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 12802 18096 12808 18148
rect 12860 18096 12866 18148
rect 15010 18096 15016 18148
rect 15068 18096 15074 18148
rect 15488 18136 15516 18167
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 17494 18164 17500 18216
rect 17552 18164 17558 18216
rect 17586 18164 17592 18216
rect 17644 18204 17650 18216
rect 18432 18204 18460 18244
rect 17644 18176 18460 18204
rect 18877 18207 18935 18213
rect 17644 18164 17650 18176
rect 18877 18173 18889 18207
rect 18923 18204 18935 18207
rect 19334 18204 19340 18216
rect 18923 18176 19340 18204
rect 18923 18173 18935 18176
rect 18877 18167 18935 18173
rect 19334 18164 19340 18176
rect 19392 18164 19398 18216
rect 19521 18139 19579 18145
rect 19521 18136 19533 18139
rect 15488 18108 19533 18136
rect 19521 18105 19533 18108
rect 19567 18105 19579 18139
rect 19720 18136 19748 18244
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 21928 18272 21956 18312
rect 23474 18300 23480 18312
rect 23532 18300 23538 18352
rect 25130 18340 25136 18352
rect 24610 18312 25136 18340
rect 25130 18300 25136 18312
rect 25188 18300 25194 18352
rect 25314 18300 25320 18352
rect 25372 18300 25378 18352
rect 26050 18300 26056 18352
rect 26108 18300 26114 18352
rect 28353 18343 28411 18349
rect 28353 18309 28365 18343
rect 28399 18340 28411 18343
rect 28626 18340 28632 18352
rect 28399 18312 28632 18340
rect 28399 18309 28411 18312
rect 28353 18303 28411 18309
rect 28626 18300 28632 18312
rect 28684 18300 28690 18352
rect 29638 18340 29644 18352
rect 29578 18312 29644 18340
rect 29638 18300 29644 18312
rect 29696 18300 29702 18352
rect 20027 18244 21956 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 19996 18136 20024 18235
rect 22002 18232 22008 18284
rect 22060 18232 22066 18284
rect 25332 18272 25360 18300
rect 26513 18275 26571 18281
rect 26513 18272 26525 18275
rect 25332 18244 26525 18272
rect 26513 18241 26525 18244
rect 26559 18241 26571 18275
rect 26513 18235 26571 18241
rect 27798 18232 27804 18284
rect 27856 18272 27862 18284
rect 28077 18275 28135 18281
rect 28077 18272 28089 18275
rect 27856 18244 28089 18272
rect 27856 18232 27862 18244
rect 28077 18241 28089 18244
rect 28123 18241 28135 18275
rect 28077 18235 28135 18241
rect 30650 18232 30656 18284
rect 30708 18272 30714 18284
rect 31018 18272 31024 18284
rect 30708 18244 31024 18272
rect 30708 18232 30714 18244
rect 31018 18232 31024 18244
rect 31076 18272 31082 18284
rect 31297 18275 31355 18281
rect 31297 18272 31309 18275
rect 31076 18244 31309 18272
rect 31076 18232 31082 18244
rect 31297 18241 31309 18244
rect 31343 18241 31355 18275
rect 31297 18235 31355 18241
rect 20070 18164 20076 18216
rect 20128 18164 20134 18216
rect 20806 18164 20812 18216
rect 20864 18204 20870 18216
rect 21177 18207 21235 18213
rect 21177 18204 21189 18207
rect 20864 18176 21189 18204
rect 20864 18164 20870 18176
rect 21177 18173 21189 18176
rect 21223 18173 21235 18207
rect 21177 18167 21235 18173
rect 21269 18207 21327 18213
rect 21269 18173 21281 18207
rect 21315 18173 21327 18207
rect 21269 18167 21327 18173
rect 19720 18108 20024 18136
rect 19521 18099 19579 18105
rect 20714 18096 20720 18148
rect 20772 18136 20778 18148
rect 21284 18136 21312 18167
rect 22462 18164 22468 18216
rect 22520 18204 22526 18216
rect 22557 18207 22615 18213
rect 22557 18204 22569 18207
rect 22520 18176 22569 18204
rect 22520 18164 22526 18176
rect 22557 18173 22569 18176
rect 22603 18204 22615 18207
rect 22833 18207 22891 18213
rect 22833 18204 22845 18207
rect 22603 18176 22845 18204
rect 22603 18173 22615 18176
rect 22557 18167 22615 18173
rect 22833 18173 22845 18176
rect 22879 18204 22891 18207
rect 22922 18204 22928 18216
rect 22879 18176 22928 18204
rect 22879 18173 22891 18176
rect 22833 18167 22891 18173
rect 22922 18164 22928 18176
rect 22980 18164 22986 18216
rect 23109 18207 23167 18213
rect 23109 18173 23121 18207
rect 23155 18173 23167 18207
rect 23109 18167 23167 18173
rect 23385 18207 23443 18213
rect 23385 18173 23397 18207
rect 23431 18204 23443 18207
rect 25222 18204 25228 18216
rect 23431 18176 25228 18204
rect 23431 18173 23443 18176
rect 23385 18167 23443 18173
rect 20772 18108 21312 18136
rect 20772 18096 20778 18108
rect 12618 18068 12624 18080
rect 12360 18040 12624 18068
rect 12618 18028 12624 18040
rect 12676 18028 12682 18080
rect 13357 18071 13415 18077
rect 13357 18037 13369 18071
rect 13403 18068 13415 18071
rect 13538 18068 13544 18080
rect 13403 18040 13544 18068
rect 13403 18037 13415 18040
rect 13357 18031 13415 18037
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 15746 18028 15752 18080
rect 15804 18068 15810 18080
rect 16025 18071 16083 18077
rect 16025 18068 16037 18071
rect 15804 18040 16037 18068
rect 15804 18028 15810 18040
rect 16025 18037 16037 18040
rect 16071 18037 16083 18071
rect 16025 18031 16083 18037
rect 16390 18028 16396 18080
rect 16448 18028 16454 18080
rect 16853 18071 16911 18077
rect 16853 18037 16865 18071
rect 16899 18068 16911 18071
rect 17678 18068 17684 18080
rect 16899 18040 17684 18068
rect 16899 18037 16911 18040
rect 16853 18031 16911 18037
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 19702 18028 19708 18080
rect 19760 18068 19766 18080
rect 22830 18068 22836 18080
rect 19760 18040 22836 18068
rect 19760 18028 19766 18040
rect 22830 18028 22836 18040
rect 22888 18028 22894 18080
rect 23124 18068 23152 18167
rect 25222 18164 25228 18176
rect 25280 18164 25286 18216
rect 27062 18164 27068 18216
rect 27120 18204 27126 18216
rect 30837 18207 30895 18213
rect 27120 18176 30328 18204
rect 27120 18164 27126 18176
rect 24486 18096 24492 18148
rect 24544 18136 24550 18148
rect 26786 18136 26792 18148
rect 24544 18108 26792 18136
rect 24544 18096 24550 18108
rect 26786 18096 26792 18108
rect 26844 18096 26850 18148
rect 30300 18145 30328 18176
rect 30837 18173 30849 18207
rect 30883 18204 30895 18207
rect 37734 18204 37740 18216
rect 30883 18176 37740 18204
rect 30883 18173 30895 18176
rect 30837 18167 30895 18173
rect 30285 18139 30343 18145
rect 30285 18105 30297 18139
rect 30331 18105 30343 18139
rect 30285 18099 30343 18105
rect 30374 18096 30380 18148
rect 30432 18136 30438 18148
rect 30852 18136 30880 18167
rect 37734 18164 37740 18176
rect 37792 18164 37798 18216
rect 30432 18108 30880 18136
rect 30432 18096 30438 18108
rect 24670 18068 24676 18080
rect 23124 18040 24676 18068
rect 24670 18028 24676 18040
rect 24728 18028 24734 18080
rect 27338 18028 27344 18080
rect 27396 18068 27402 18080
rect 29822 18068 29828 18080
rect 27396 18040 29828 18068
rect 27396 18028 27402 18040
rect 29822 18028 29828 18040
rect 29880 18028 29886 18080
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 3605 17867 3663 17873
rect 3605 17833 3617 17867
rect 3651 17864 3663 17867
rect 8386 17864 8392 17876
rect 3651 17836 8392 17864
rect 3651 17833 3663 17836
rect 3605 17827 3663 17833
rect 8386 17824 8392 17836
rect 8444 17864 8450 17876
rect 8938 17864 8944 17876
rect 8444 17836 8944 17864
rect 8444 17824 8450 17836
rect 8938 17824 8944 17836
rect 8996 17824 9002 17876
rect 10134 17864 10140 17876
rect 9646 17836 10140 17864
rect 1854 17756 1860 17808
rect 1912 17796 1918 17808
rect 4433 17799 4491 17805
rect 4433 17796 4445 17799
rect 1912 17768 4445 17796
rect 1912 17756 1918 17768
rect 4433 17765 4445 17768
rect 4479 17765 4491 17799
rect 4433 17759 4491 17765
rect 6178 17756 6184 17808
rect 6236 17796 6242 17808
rect 6641 17799 6699 17805
rect 6641 17796 6653 17799
rect 6236 17768 6653 17796
rect 6236 17756 6242 17768
rect 6641 17765 6653 17768
rect 6687 17765 6699 17799
rect 6641 17759 6699 17765
rect 7190 17756 7196 17808
rect 7248 17796 7254 17808
rect 7558 17796 7564 17808
rect 7248 17768 7564 17796
rect 7248 17756 7254 17768
rect 7558 17756 7564 17768
rect 7616 17756 7622 17808
rect 7834 17756 7840 17808
rect 7892 17756 7898 17808
rect 9646 17796 9674 17836
rect 10134 17824 10140 17836
rect 10192 17824 10198 17876
rect 10318 17824 10324 17876
rect 10376 17864 10382 17876
rect 10597 17867 10655 17873
rect 10597 17864 10609 17867
rect 10376 17836 10609 17864
rect 10376 17824 10382 17836
rect 10597 17833 10609 17836
rect 10643 17833 10655 17867
rect 10597 17827 10655 17833
rect 12342 17824 12348 17876
rect 12400 17864 12406 17876
rect 13725 17867 13783 17873
rect 13725 17864 13737 17867
rect 12400 17836 13737 17864
rect 12400 17824 12406 17836
rect 13725 17833 13737 17836
rect 13771 17833 13783 17867
rect 13725 17827 13783 17833
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 16390 17864 16396 17876
rect 15252 17836 16396 17864
rect 15252 17824 15258 17836
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 16666 17824 16672 17876
rect 16724 17864 16730 17876
rect 21174 17864 21180 17876
rect 16724 17836 21180 17864
rect 16724 17824 16730 17836
rect 21174 17824 21180 17836
rect 21232 17824 21238 17876
rect 21266 17824 21272 17876
rect 21324 17864 21330 17876
rect 21726 17864 21732 17876
rect 21324 17836 21732 17864
rect 21324 17824 21330 17836
rect 21726 17824 21732 17836
rect 21784 17864 21790 17876
rect 21913 17867 21971 17873
rect 21913 17864 21925 17867
rect 21784 17836 21925 17864
rect 21784 17824 21790 17836
rect 21913 17833 21925 17836
rect 21959 17864 21971 17867
rect 23750 17864 23756 17876
rect 21959 17836 23756 17864
rect 21959 17833 21971 17836
rect 21913 17827 21971 17833
rect 23750 17824 23756 17836
rect 23808 17824 23814 17876
rect 30929 17867 30987 17873
rect 30929 17864 30941 17867
rect 23860 17836 30941 17864
rect 8404 17768 9674 17796
rect 1118 17728 1124 17740
rect 1044 17700 1124 17728
rect 1118 17688 1124 17700
rect 1176 17688 1182 17740
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 1780 17700 7389 17728
rect 1780 17669 1808 17700
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7576 17728 7604 17756
rect 8404 17737 8432 17768
rect 9766 17756 9772 17808
rect 9824 17796 9830 17808
rect 11882 17796 11888 17808
rect 9824 17768 11888 17796
rect 9824 17756 9830 17768
rect 11882 17756 11888 17768
rect 11940 17756 11946 17808
rect 13262 17756 13268 17808
rect 13320 17796 13326 17808
rect 16206 17796 16212 17808
rect 13320 17768 16212 17796
rect 13320 17756 13326 17768
rect 16206 17756 16212 17768
rect 16264 17756 16270 17808
rect 17586 17756 17592 17808
rect 17644 17796 17650 17808
rect 20717 17799 20775 17805
rect 20717 17796 20729 17799
rect 17644 17768 20729 17796
rect 17644 17756 17650 17768
rect 20717 17765 20729 17768
rect 20763 17765 20775 17799
rect 20717 17759 20775 17765
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7576 17700 8401 17728
rect 7377 17691 7435 17697
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 9732 17700 9873 17728
rect 9732 17688 9738 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 10042 17688 10048 17740
rect 10100 17728 10106 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10100 17700 11161 17728
rect 10100 17688 10106 17700
rect 11149 17697 11161 17700
rect 11195 17697 11207 17731
rect 11149 17691 11207 17697
rect 12253 17731 12311 17737
rect 12253 17697 12265 17731
rect 12299 17728 12311 17731
rect 12894 17728 12900 17740
rect 12299 17700 12900 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 12894 17688 12900 17700
rect 12952 17728 12958 17740
rect 13630 17728 13636 17740
rect 12952 17700 13636 17728
rect 12952 17688 12958 17700
rect 13630 17688 13636 17700
rect 13688 17688 13694 17740
rect 16298 17688 16304 17740
rect 16356 17688 16362 17740
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 16942 17728 16948 17740
rect 16623 17700 16948 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 16942 17688 16948 17700
rect 17000 17688 17006 17740
rect 18966 17688 18972 17740
rect 19024 17728 19030 17740
rect 19429 17731 19487 17737
rect 19429 17728 19441 17731
rect 19024 17700 19441 17728
rect 19024 17688 19030 17700
rect 19429 17697 19441 17700
rect 19475 17697 19487 17731
rect 19429 17691 19487 17697
rect 19610 17688 19616 17740
rect 19668 17728 19674 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 19668 17700 19717 17728
rect 19668 17688 19674 17700
rect 19705 17697 19717 17700
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 20346 17688 20352 17740
rect 20404 17728 20410 17740
rect 21269 17731 21327 17737
rect 21269 17728 21281 17731
rect 20404 17700 21281 17728
rect 20404 17688 20410 17700
rect 21269 17697 21281 17700
rect 21315 17728 21327 17731
rect 23750 17728 23756 17740
rect 21315 17700 23756 17728
rect 21315 17697 21327 17700
rect 21269 17691 21327 17697
rect 23750 17688 23756 17700
rect 23808 17688 23814 17740
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17629 1823 17663
rect 1765 17623 1823 17629
rect 3786 17620 3792 17672
rect 3844 17620 3850 17672
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4614 17660 4620 17672
rect 4212 17632 4620 17660
rect 4212 17620 4218 17632
rect 4614 17620 4620 17632
rect 4672 17660 4678 17672
rect 4893 17663 4951 17669
rect 4893 17660 4905 17663
rect 4672 17632 4905 17660
rect 4672 17620 4678 17632
rect 4893 17629 4905 17632
rect 4939 17629 4951 17663
rect 4893 17623 4951 17629
rect 7098 17620 7104 17672
rect 7156 17660 7162 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7156 17632 8217 17660
rect 7156 17620 7162 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8205 17623 8263 17629
rect 8938 17620 8944 17672
rect 8996 17660 9002 17672
rect 9122 17660 9128 17672
rect 8996 17632 9128 17660
rect 8996 17620 9002 17632
rect 9122 17620 9128 17632
rect 9180 17620 9186 17672
rect 9490 17620 9496 17672
rect 9548 17660 9554 17672
rect 11057 17663 11115 17669
rect 11057 17660 11069 17663
rect 9548 17632 11069 17660
rect 9548 17620 9554 17632
rect 11057 17629 11069 17632
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 11698 17620 11704 17672
rect 11756 17620 11762 17672
rect 11974 17620 11980 17672
rect 12032 17620 12038 17672
rect 19334 17620 19340 17672
rect 19392 17660 19398 17672
rect 21085 17663 21143 17669
rect 21085 17660 21097 17663
rect 19392 17632 21097 17660
rect 19392 17620 19398 17632
rect 21085 17629 21097 17632
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 22002 17620 22008 17672
rect 22060 17660 22066 17672
rect 22281 17663 22339 17669
rect 22281 17660 22293 17663
rect 22060 17632 22293 17660
rect 22060 17620 22066 17632
rect 22281 17629 22293 17632
rect 22327 17629 22339 17663
rect 22281 17623 22339 17629
rect 23658 17620 23664 17672
rect 23716 17620 23722 17672
rect 1210 17552 1216 17604
rect 1268 17592 1274 17604
rect 2501 17595 2559 17601
rect 2501 17592 2513 17595
rect 1268 17564 2513 17592
rect 1268 17552 1274 17564
rect 2501 17561 2513 17564
rect 2547 17561 2559 17595
rect 2501 17555 2559 17561
rect 3421 17595 3479 17601
rect 3421 17561 3433 17595
rect 3467 17592 3479 17595
rect 4062 17592 4068 17604
rect 3467 17564 4068 17592
rect 3467 17561 3479 17564
rect 3421 17555 3479 17561
rect 4062 17552 4068 17564
rect 4120 17552 4126 17604
rect 4249 17595 4307 17601
rect 4249 17561 4261 17595
rect 4295 17592 4307 17595
rect 4798 17592 4804 17604
rect 4295 17564 4804 17592
rect 4295 17561 4307 17564
rect 4249 17555 4307 17561
rect 4798 17552 4804 17564
rect 4856 17552 4862 17604
rect 5169 17595 5227 17601
rect 5169 17561 5181 17595
rect 5215 17561 5227 17595
rect 5169 17555 5227 17561
rect 5184 17524 5212 17555
rect 5442 17552 5448 17604
rect 5500 17592 5506 17604
rect 5500 17564 5658 17592
rect 5500 17552 5506 17564
rect 7190 17552 7196 17604
rect 7248 17552 7254 17604
rect 8297 17595 8355 17601
rect 8297 17561 8309 17595
rect 8343 17592 8355 17595
rect 9398 17592 9404 17604
rect 8343 17564 9404 17592
rect 8343 17561 8355 17564
rect 8297 17555 8355 17561
rect 9398 17552 9404 17564
rect 9456 17552 9462 17604
rect 10965 17595 11023 17601
rect 10965 17561 10977 17595
rect 11011 17592 11023 17595
rect 12250 17592 12256 17604
rect 11011 17564 12256 17592
rect 11011 17561 11023 17564
rect 10965 17555 11023 17561
rect 12250 17552 12256 17564
rect 12308 17552 12314 17604
rect 13538 17592 13544 17604
rect 13478 17564 13544 17592
rect 13538 17552 13544 17564
rect 13596 17592 13602 17604
rect 13998 17592 14004 17604
rect 13596 17564 14004 17592
rect 13596 17552 13602 17564
rect 13998 17552 14004 17564
rect 14056 17552 14062 17604
rect 14369 17595 14427 17601
rect 14369 17561 14381 17595
rect 14415 17592 14427 17595
rect 18325 17595 18383 17601
rect 18325 17592 18337 17595
rect 14415 17564 14964 17592
rect 14415 17561 14427 17564
rect 14369 17555 14427 17561
rect 7374 17524 7380 17536
rect 5184 17496 7380 17524
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 8018 17484 8024 17536
rect 8076 17524 8082 17536
rect 14274 17524 14280 17536
rect 8076 17496 14280 17524
rect 8076 17484 8082 17496
rect 14274 17484 14280 17496
rect 14332 17484 14338 17536
rect 14458 17484 14464 17536
rect 14516 17484 14522 17536
rect 14936 17533 14964 17564
rect 16408 17564 17066 17592
rect 17880 17564 18337 17592
rect 16408 17536 16436 17564
rect 14921 17527 14979 17533
rect 14921 17493 14933 17527
rect 14967 17524 14979 17527
rect 15010 17524 15016 17536
rect 14967 17496 15016 17524
rect 14967 17493 14979 17496
rect 14921 17487 14979 17493
rect 15010 17484 15016 17496
rect 15068 17484 15074 17536
rect 15102 17484 15108 17536
rect 15160 17484 15166 17536
rect 15378 17484 15384 17536
rect 15436 17484 15442 17536
rect 16022 17484 16028 17536
rect 16080 17524 16086 17536
rect 16390 17524 16396 17536
rect 16080 17496 16396 17524
rect 16080 17484 16086 17496
rect 16390 17484 16396 17496
rect 16448 17484 16454 17536
rect 16960 17524 16988 17564
rect 17880 17524 17908 17564
rect 18325 17561 18337 17564
rect 18371 17561 18383 17595
rect 20714 17592 20720 17604
rect 18325 17555 18383 17561
rect 18524 17564 20720 17592
rect 18524 17536 18552 17564
rect 20714 17552 20720 17564
rect 20772 17552 20778 17604
rect 21177 17595 21235 17601
rect 21177 17561 21189 17595
rect 21223 17592 21235 17595
rect 21223 17564 22094 17592
rect 21223 17561 21235 17564
rect 21177 17555 21235 17561
rect 16960 17496 17908 17524
rect 18049 17527 18107 17533
rect 18049 17493 18061 17527
rect 18095 17524 18107 17527
rect 18506 17524 18512 17536
rect 18095 17496 18512 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 18506 17484 18512 17496
rect 18564 17484 18570 17536
rect 18693 17527 18751 17533
rect 18693 17493 18705 17527
rect 18739 17524 18751 17527
rect 20438 17524 20444 17536
rect 18739 17496 20444 17524
rect 18739 17493 18751 17496
rect 18693 17487 18751 17493
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 20990 17484 20996 17536
rect 21048 17524 21054 17536
rect 21729 17527 21787 17533
rect 21729 17524 21741 17527
rect 21048 17496 21741 17524
rect 21048 17484 21054 17496
rect 21729 17493 21741 17496
rect 21775 17524 21787 17527
rect 21818 17524 21824 17536
rect 21775 17496 21824 17524
rect 21775 17493 21787 17496
rect 21729 17487 21787 17493
rect 21818 17484 21824 17496
rect 21876 17484 21882 17536
rect 22066 17524 22094 17564
rect 22554 17552 22560 17604
rect 22612 17552 22618 17604
rect 23860 17524 23888 17836
rect 30929 17833 30941 17836
rect 30975 17833 30987 17867
rect 30929 17827 30987 17833
rect 26602 17756 26608 17808
rect 26660 17756 26666 17808
rect 28442 17756 28448 17808
rect 28500 17796 28506 17808
rect 29733 17799 29791 17805
rect 29733 17796 29745 17799
rect 28500 17768 29745 17796
rect 28500 17756 28506 17768
rect 29733 17765 29745 17768
rect 29779 17765 29791 17799
rect 29733 17759 29791 17765
rect 24670 17688 24676 17740
rect 24728 17728 24734 17740
rect 24857 17731 24915 17737
rect 24857 17728 24869 17731
rect 24728 17700 24869 17728
rect 24728 17688 24734 17700
rect 24857 17697 24869 17700
rect 24903 17728 24915 17731
rect 25774 17728 25780 17740
rect 24903 17700 25780 17728
rect 24903 17697 24915 17700
rect 24857 17691 24915 17697
rect 25774 17688 25780 17700
rect 25832 17728 25838 17740
rect 27065 17731 27123 17737
rect 27065 17728 27077 17731
rect 25832 17700 27077 17728
rect 25832 17688 25838 17700
rect 27065 17697 27077 17700
rect 27111 17728 27123 17731
rect 27798 17728 27804 17740
rect 27111 17700 27804 17728
rect 27111 17697 27123 17700
rect 27065 17691 27123 17697
rect 27798 17688 27804 17700
rect 27856 17688 27862 17740
rect 28813 17731 28871 17737
rect 28813 17697 28825 17731
rect 28859 17697 28871 17731
rect 28813 17691 28871 17697
rect 29181 17731 29239 17737
rect 29181 17697 29193 17731
rect 29227 17728 29239 17731
rect 29638 17728 29644 17740
rect 29227 17700 29644 17728
rect 29227 17697 29239 17700
rect 29181 17691 29239 17697
rect 28828 17660 28856 17691
rect 29638 17688 29644 17700
rect 29696 17688 29702 17740
rect 30282 17688 30288 17740
rect 30340 17688 30346 17740
rect 31481 17731 31539 17737
rect 31481 17728 31493 17731
rect 30392 17700 31493 17728
rect 29086 17660 29092 17672
rect 28828 17632 29092 17660
rect 29086 17620 29092 17632
rect 29144 17660 29150 17672
rect 30392 17660 30420 17700
rect 31481 17697 31493 17700
rect 31527 17697 31539 17731
rect 31481 17691 31539 17697
rect 29144 17632 30420 17660
rect 29144 17620 29150 17632
rect 30834 17620 30840 17672
rect 30892 17660 30898 17672
rect 31294 17660 31300 17672
rect 30892 17632 31300 17660
rect 30892 17620 30898 17632
rect 31294 17620 31300 17632
rect 31352 17620 31358 17672
rect 31389 17663 31447 17669
rect 31389 17629 31401 17663
rect 31435 17660 31447 17663
rect 37366 17660 37372 17672
rect 31435 17632 37372 17660
rect 31435 17629 31447 17632
rect 31389 17623 31447 17629
rect 37366 17620 37372 17632
rect 37424 17620 37430 17672
rect 25130 17592 25136 17604
rect 24044 17564 25136 17592
rect 24044 17533 24072 17564
rect 25130 17552 25136 17564
rect 25188 17552 25194 17604
rect 26970 17592 26976 17604
rect 26358 17564 26976 17592
rect 26970 17552 26976 17564
rect 27028 17552 27034 17604
rect 27338 17552 27344 17604
rect 27396 17552 27402 17604
rect 29638 17592 29644 17604
rect 28566 17564 29644 17592
rect 29638 17552 29644 17564
rect 29696 17552 29702 17604
rect 30101 17595 30159 17601
rect 30101 17561 30113 17595
rect 30147 17592 30159 17595
rect 30926 17592 30932 17604
rect 30147 17564 30932 17592
rect 30147 17561 30159 17564
rect 30101 17555 30159 17561
rect 22066 17496 23888 17524
rect 24029 17527 24087 17533
rect 24029 17493 24041 17527
rect 24075 17493 24087 17527
rect 24029 17487 24087 17493
rect 24394 17484 24400 17536
rect 24452 17524 24458 17536
rect 30116 17524 30144 17555
rect 30926 17552 30932 17564
rect 30984 17552 30990 17604
rect 24452 17496 30144 17524
rect 24452 17484 24458 17496
rect 30190 17484 30196 17536
rect 30248 17484 30254 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 3970 17280 3976 17332
rect 4028 17320 4034 17332
rect 4890 17320 4896 17332
rect 4028 17292 4896 17320
rect 4028 17280 4034 17292
rect 4890 17280 4896 17292
rect 4948 17320 4954 17332
rect 5077 17323 5135 17329
rect 5077 17320 5089 17323
rect 4948 17292 5089 17320
rect 4948 17280 4954 17292
rect 5077 17289 5089 17292
rect 5123 17320 5135 17323
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 5123 17292 5641 17320
rect 5123 17289 5135 17292
rect 5077 17283 5135 17289
rect 5629 17289 5641 17292
rect 5675 17289 5687 17323
rect 5629 17283 5687 17289
rect 6822 17280 6828 17332
rect 6880 17280 6886 17332
rect 7742 17280 7748 17332
rect 7800 17320 7806 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7800 17292 8033 17320
rect 7800 17280 7806 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 11885 17323 11943 17329
rect 11885 17320 11897 17323
rect 8021 17283 8079 17289
rect 8128 17292 11897 17320
rect 4338 17212 4344 17264
rect 4396 17212 4402 17264
rect 7193 17255 7251 17261
rect 7193 17221 7205 17255
rect 7239 17252 7251 17255
rect 7282 17252 7288 17264
rect 7239 17224 7288 17252
rect 7239 17221 7251 17224
rect 7193 17215 7251 17221
rect 7282 17212 7288 17224
rect 7340 17212 7346 17264
rect 1762 17144 1768 17196
rect 1820 17144 1826 17196
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 8128 17184 8156 17292
rect 11885 17289 11897 17292
rect 11931 17289 11943 17323
rect 11885 17283 11943 17289
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12529 17323 12587 17329
rect 12529 17320 12541 17323
rect 12492 17292 12541 17320
rect 12492 17280 12498 17292
rect 12529 17289 12541 17292
rect 12575 17289 12587 17323
rect 13354 17320 13360 17332
rect 12529 17283 12587 17289
rect 12728 17292 13360 17320
rect 9582 17212 9588 17264
rect 9640 17252 9646 17264
rect 9953 17255 10011 17261
rect 9953 17252 9965 17255
rect 9640 17224 9965 17252
rect 9640 17212 9646 17224
rect 9953 17221 9965 17224
rect 9999 17221 10011 17255
rect 9953 17215 10011 17221
rect 10781 17255 10839 17261
rect 10781 17221 10793 17255
rect 10827 17252 10839 17255
rect 12728 17252 12756 17292
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 13722 17280 13728 17332
rect 13780 17280 13786 17332
rect 14274 17280 14280 17332
rect 14332 17320 14338 17332
rect 16117 17323 16175 17329
rect 16117 17320 16129 17323
rect 14332 17292 16129 17320
rect 14332 17280 14338 17292
rect 16117 17289 16129 17292
rect 16163 17289 16175 17323
rect 16117 17283 16175 17289
rect 16206 17280 16212 17332
rect 16264 17320 16270 17332
rect 17126 17320 17132 17332
rect 16264 17292 17132 17320
rect 16264 17280 16270 17292
rect 17126 17280 17132 17292
rect 17184 17280 17190 17332
rect 17862 17280 17868 17332
rect 17920 17320 17926 17332
rect 22005 17323 22063 17329
rect 22005 17320 22017 17323
rect 17920 17292 22017 17320
rect 17920 17280 17926 17292
rect 22005 17289 22017 17292
rect 22051 17289 22063 17323
rect 22005 17283 22063 17289
rect 22373 17323 22431 17329
rect 22373 17289 22385 17323
rect 22419 17320 22431 17323
rect 22462 17320 22468 17332
rect 22419 17292 22468 17320
rect 22419 17289 22431 17292
rect 22373 17283 22431 17289
rect 22462 17280 22468 17292
rect 22520 17280 22526 17332
rect 24394 17320 24400 17332
rect 23676 17292 24400 17320
rect 10827 17224 12756 17252
rect 10827 17221 10839 17224
rect 10781 17215 10839 17221
rect 3651 17156 8156 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 8386 17144 8392 17196
rect 8444 17144 8450 17196
rect 8754 17184 8760 17196
rect 8680 17156 8760 17184
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1360 17088 2053 17116
rect 1360 17076 1366 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 3510 17076 3516 17128
rect 3568 17116 3574 17128
rect 4614 17116 4620 17128
rect 3568 17088 4620 17116
rect 3568 17076 3574 17088
rect 4614 17076 4620 17088
rect 4672 17116 4678 17128
rect 5721 17119 5779 17125
rect 5721 17116 5733 17119
rect 4672 17088 5733 17116
rect 4672 17076 4678 17088
rect 5721 17085 5733 17088
rect 5767 17085 5779 17119
rect 5721 17079 5779 17085
rect 5902 17076 5908 17128
rect 5960 17116 5966 17128
rect 6362 17116 6368 17128
rect 5960 17088 6368 17116
rect 5960 17076 5966 17088
rect 6362 17076 6368 17088
rect 6420 17076 6426 17128
rect 6454 17076 6460 17128
rect 6512 17076 6518 17128
rect 7285 17119 7343 17125
rect 7285 17085 7297 17119
rect 7331 17085 7343 17119
rect 7285 17079 7343 17085
rect 7469 17119 7527 17125
rect 7469 17085 7481 17119
rect 7515 17116 7527 17119
rect 7558 17116 7564 17128
rect 7515 17088 7564 17116
rect 7515 17085 7527 17088
rect 7469 17079 7527 17085
rect 5261 17051 5319 17057
rect 5261 17017 5273 17051
rect 5307 17048 5319 17051
rect 7300 17048 7328 17079
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 8481 17119 8539 17125
rect 8481 17085 8493 17119
rect 8527 17116 8539 17119
rect 8570 17116 8576 17128
rect 8527 17088 8576 17116
rect 8527 17085 8539 17088
rect 8481 17079 8539 17085
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 8680 17125 8708 17156
rect 8754 17144 8760 17156
rect 8812 17144 8818 17196
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 9364 17156 9674 17184
rect 9364 17144 9370 17156
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17085 8723 17119
rect 9646 17116 9674 17156
rect 9858 17144 9864 17196
rect 9916 17144 9922 17196
rect 9968 17184 9996 17215
rect 12802 17212 12808 17264
rect 12860 17252 12866 17264
rect 14185 17255 14243 17261
rect 14185 17252 14197 17255
rect 12860 17224 14197 17252
rect 12860 17212 12866 17224
rect 14185 17221 14197 17224
rect 14231 17252 14243 17255
rect 14737 17255 14795 17261
rect 14737 17252 14749 17255
rect 14231 17224 14749 17252
rect 14231 17221 14243 17224
rect 14185 17215 14243 17221
rect 14737 17221 14749 17224
rect 14783 17221 14795 17255
rect 17770 17252 17776 17264
rect 14737 17215 14795 17221
rect 14936 17224 17776 17252
rect 9968 17156 11744 17184
rect 10045 17119 10103 17125
rect 10045 17116 10057 17119
rect 9646 17088 10057 17116
rect 8665 17079 8723 17085
rect 10045 17085 10057 17088
rect 10091 17116 10103 17119
rect 10318 17116 10324 17128
rect 10091 17088 10324 17116
rect 10091 17085 10103 17088
rect 10045 17079 10103 17085
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 11716 17116 11744 17156
rect 11790 17144 11796 17196
rect 11848 17144 11854 17196
rect 12897 17187 12955 17193
rect 12897 17184 12909 17187
rect 12406 17156 12909 17184
rect 12250 17116 12256 17128
rect 11716 17088 12256 17116
rect 12250 17076 12256 17088
rect 12308 17116 12314 17128
rect 12406 17116 12434 17156
rect 12897 17153 12909 17156
rect 12943 17153 12955 17187
rect 12897 17147 12955 17153
rect 12989 17187 13047 17193
rect 12989 17153 13001 17187
rect 13035 17184 13047 17187
rect 13035 17156 13860 17184
rect 13035 17153 13047 17156
rect 12989 17147 13047 17153
rect 12308 17088 12434 17116
rect 13081 17119 13139 17125
rect 12308 17076 12314 17088
rect 13081 17085 13093 17119
rect 13127 17085 13139 17119
rect 13832 17116 13860 17156
rect 13906 17144 13912 17196
rect 13964 17184 13970 17196
rect 14936 17193 14964 17224
rect 17770 17212 17776 17224
rect 17828 17212 17834 17264
rect 18138 17212 18144 17264
rect 18196 17252 18202 17264
rect 18417 17255 18475 17261
rect 18417 17252 18429 17255
rect 18196 17224 18429 17252
rect 18196 17212 18202 17224
rect 18417 17221 18429 17224
rect 18463 17252 18475 17255
rect 18506 17252 18512 17264
rect 18463 17224 18512 17252
rect 18463 17221 18475 17224
rect 18417 17215 18475 17221
rect 18506 17212 18512 17224
rect 18564 17212 18570 17264
rect 22554 17252 22560 17264
rect 20180 17224 22560 17252
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 13964 17156 14105 17184
rect 13964 17144 13970 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 14921 17187 14979 17193
rect 14921 17184 14933 17187
rect 14093 17147 14151 17153
rect 14292 17156 14933 17184
rect 14292 17116 14320 17156
rect 14921 17153 14933 17156
rect 14967 17153 14979 17187
rect 14921 17147 14979 17153
rect 15654 17144 15660 17196
rect 15712 17144 15718 17196
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17184 16359 17187
rect 16666 17184 16672 17196
rect 16347 17156 16672 17184
rect 16347 17153 16359 17156
rect 16301 17147 16359 17153
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 17218 17144 17224 17196
rect 17276 17144 17282 17196
rect 19794 17184 19800 17196
rect 19550 17156 19800 17184
rect 19794 17144 19800 17156
rect 19852 17144 19858 17196
rect 13832 17088 14320 17116
rect 14369 17119 14427 17125
rect 13081 17079 13139 17085
rect 14369 17085 14381 17119
rect 14415 17116 14427 17119
rect 15286 17116 15292 17128
rect 14415 17088 15292 17116
rect 14415 17085 14427 17088
rect 14369 17079 14427 17085
rect 5307 17020 7328 17048
rect 5307 17017 5319 17020
rect 5261 17011 5319 17017
rect 8754 17008 8760 17060
rect 8812 17048 8818 17060
rect 9493 17051 9551 17057
rect 9493 17048 9505 17051
rect 8812 17020 9505 17048
rect 8812 17008 8818 17020
rect 9493 17017 9505 17020
rect 9539 17017 9551 17051
rect 9493 17011 9551 17017
rect 12342 17008 12348 17060
rect 12400 17048 12406 17060
rect 13096 17048 13124 17079
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 15838 17076 15844 17128
rect 15896 17116 15902 17128
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 15896 17088 17325 17116
rect 15896 17076 15902 17088
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17402 17076 17408 17128
rect 17460 17076 17466 17128
rect 18141 17119 18199 17125
rect 18141 17085 18153 17119
rect 18187 17085 18199 17119
rect 20180 17116 20208 17224
rect 22554 17212 22560 17224
rect 22612 17212 22618 17264
rect 20622 17144 20628 17196
rect 20680 17184 20686 17196
rect 21082 17184 21088 17196
rect 20680 17156 21088 17184
rect 20680 17144 20686 17156
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 21266 17144 21272 17196
rect 21324 17184 21330 17196
rect 23676 17193 23704 17292
rect 24394 17280 24400 17292
rect 24452 17280 24458 17332
rect 29086 17320 29092 17332
rect 24964 17292 29092 17320
rect 23750 17212 23756 17264
rect 23808 17212 23814 17264
rect 24964 17261 24992 17292
rect 29086 17280 29092 17292
rect 29144 17280 29150 17332
rect 29638 17280 29644 17332
rect 29696 17320 29702 17332
rect 29825 17323 29883 17329
rect 29825 17320 29837 17323
rect 29696 17292 29837 17320
rect 29696 17280 29702 17292
rect 29825 17289 29837 17292
rect 29871 17289 29883 17323
rect 29825 17283 29883 17289
rect 30190 17280 30196 17332
rect 30248 17320 30254 17332
rect 30561 17323 30619 17329
rect 30561 17320 30573 17323
rect 30248 17292 30573 17320
rect 30248 17280 30254 17292
rect 30561 17289 30573 17292
rect 30607 17289 30619 17323
rect 30561 17283 30619 17289
rect 30834 17280 30840 17332
rect 30892 17280 30898 17332
rect 30926 17280 30932 17332
rect 30984 17280 30990 17332
rect 24949 17255 25007 17261
rect 24949 17221 24961 17255
rect 24995 17221 25007 17255
rect 26789 17255 26847 17261
rect 26789 17252 26801 17255
rect 26174 17224 26801 17252
rect 24949 17215 25007 17221
rect 26789 17221 26801 17224
rect 26835 17252 26847 17255
rect 26970 17252 26976 17264
rect 26835 17224 26976 17252
rect 26835 17221 26847 17224
rect 26789 17215 26847 17221
rect 26970 17212 26976 17224
rect 27028 17212 27034 17264
rect 29656 17252 29684 17280
rect 29302 17224 31708 17252
rect 23661 17187 23719 17193
rect 23661 17184 23673 17187
rect 21324 17156 23673 17184
rect 21324 17144 21330 17156
rect 23661 17153 23673 17156
rect 23707 17153 23719 17187
rect 23768 17184 23796 17212
rect 24397 17187 24455 17193
rect 23768 17156 24256 17184
rect 23661 17147 23719 17153
rect 18141 17079 18199 17085
rect 19904 17088 20208 17116
rect 21177 17119 21235 17125
rect 12400 17020 13124 17048
rect 12400 17008 12406 17020
rect 13446 17008 13452 17060
rect 13504 17048 13510 17060
rect 15473 17051 15531 17057
rect 15473 17048 15485 17051
rect 13504 17020 15485 17048
rect 13504 17008 13510 17020
rect 15473 17017 15485 17020
rect 15519 17017 15531 17051
rect 15473 17011 15531 17017
rect 17034 17008 17040 17060
rect 17092 17048 17098 17060
rect 18156 17048 18184 17079
rect 17092 17020 18184 17048
rect 17092 17008 17098 17020
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 9125 16983 9183 16989
rect 9125 16980 9137 16983
rect 3384 16952 9137 16980
rect 3384 16940 3390 16952
rect 9125 16949 9137 16952
rect 9171 16980 9183 16983
rect 9766 16980 9772 16992
rect 9171 16952 9772 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 9766 16940 9772 16952
rect 9824 16980 9830 16992
rect 10502 16980 10508 16992
rect 9824 16952 10508 16980
rect 9824 16940 9830 16952
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 10870 16940 10876 16992
rect 10928 16940 10934 16992
rect 11333 16983 11391 16989
rect 11333 16949 11345 16983
rect 11379 16980 11391 16983
rect 11606 16980 11612 16992
rect 11379 16952 11612 16980
rect 11379 16949 11391 16952
rect 11333 16943 11391 16949
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 12066 16940 12072 16992
rect 12124 16980 12130 16992
rect 13722 16980 13728 16992
rect 12124 16952 13728 16980
rect 12124 16940 12130 16952
rect 13722 16940 13728 16952
rect 13780 16940 13786 16992
rect 15197 16983 15255 16989
rect 15197 16949 15209 16983
rect 15243 16980 15255 16983
rect 15286 16980 15292 16992
rect 15243 16952 15292 16980
rect 15243 16949 15255 16952
rect 15197 16943 15255 16949
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 16850 16940 16856 16992
rect 16908 16940 16914 16992
rect 17494 16940 17500 16992
rect 17552 16980 17558 16992
rect 19904 16989 19932 17088
rect 21177 17085 21189 17119
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 21361 17119 21419 17125
rect 21361 17085 21373 17119
rect 21407 17085 21419 17119
rect 21361 17079 21419 17085
rect 20070 17008 20076 17060
rect 20128 17048 20134 17060
rect 20349 17051 20407 17057
rect 20349 17048 20361 17051
rect 20128 17020 20361 17048
rect 20128 17008 20134 17020
rect 20349 17017 20361 17020
rect 20395 17048 20407 17051
rect 21192 17048 21220 17079
rect 20395 17020 21220 17048
rect 21376 17048 21404 17079
rect 21726 17076 21732 17128
rect 21784 17116 21790 17128
rect 22465 17119 22523 17125
rect 22465 17116 22477 17119
rect 21784 17088 22477 17116
rect 21784 17076 21790 17088
rect 22465 17085 22477 17088
rect 22511 17085 22523 17119
rect 22465 17079 22523 17085
rect 22554 17076 22560 17128
rect 22612 17076 22618 17128
rect 23750 17076 23756 17128
rect 23808 17076 23814 17128
rect 23845 17119 23903 17125
rect 23845 17085 23857 17119
rect 23891 17085 23903 17119
rect 24228 17116 24256 17156
rect 24397 17153 24409 17187
rect 24443 17184 24455 17187
rect 24486 17184 24492 17196
rect 24443 17156 24492 17184
rect 24443 17153 24455 17156
rect 24397 17147 24455 17153
rect 24486 17144 24492 17156
rect 24544 17144 24550 17196
rect 24670 17144 24676 17196
rect 24728 17144 24734 17196
rect 27798 17144 27804 17196
rect 27856 17144 27862 17196
rect 31680 17184 31708 17224
rect 37274 17212 37280 17264
rect 37332 17252 37338 17264
rect 48498 17252 48504 17264
rect 37332 17224 48504 17252
rect 37332 17212 37338 17224
rect 48498 17212 48504 17224
rect 48556 17212 48562 17264
rect 31754 17184 31760 17196
rect 31680 17156 31760 17184
rect 31754 17144 31760 17156
rect 31812 17144 31818 17196
rect 26421 17119 26479 17125
rect 26421 17116 26433 17119
rect 24228 17088 26433 17116
rect 23845 17079 23903 17085
rect 26421 17085 26433 17088
rect 26467 17085 26479 17119
rect 26421 17079 26479 17085
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17116 27215 17119
rect 27614 17116 27620 17128
rect 27203 17088 27620 17116
rect 27203 17085 27215 17088
rect 27157 17079 27215 17085
rect 22186 17048 22192 17060
rect 21376 17020 22192 17048
rect 20395 17017 20407 17020
rect 20349 17011 20407 17017
rect 19889 16983 19947 16989
rect 19889 16980 19901 16983
rect 17552 16952 19901 16980
rect 17552 16940 17558 16952
rect 19889 16949 19901 16952
rect 19935 16949 19947 16983
rect 19889 16943 19947 16949
rect 20162 16940 20168 16992
rect 20220 16980 20226 16992
rect 20622 16980 20628 16992
rect 20220 16952 20628 16980
rect 20220 16940 20226 16952
rect 20622 16940 20628 16952
rect 20680 16940 20686 16992
rect 20714 16940 20720 16992
rect 20772 16940 20778 16992
rect 21192 16980 21220 17020
rect 22186 17008 22192 17020
rect 22244 17048 22250 17060
rect 23860 17048 23888 17079
rect 27614 17076 27620 17088
rect 27672 17076 27678 17128
rect 28077 17119 28135 17125
rect 28077 17085 28089 17119
rect 28123 17116 28135 17119
rect 30282 17116 30288 17128
rect 28123 17088 30288 17116
rect 28123 17085 28135 17088
rect 28077 17079 28135 17085
rect 30282 17076 30288 17088
rect 30340 17076 30346 17128
rect 22244 17020 23888 17048
rect 22244 17008 22250 17020
rect 30190 17008 30196 17060
rect 30248 17048 30254 17060
rect 30248 17020 30880 17048
rect 30248 17008 30254 17020
rect 21542 16980 21548 16992
rect 21192 16952 21548 16980
rect 21542 16940 21548 16952
rect 21600 16940 21606 16992
rect 21726 16940 21732 16992
rect 21784 16980 21790 16992
rect 22554 16980 22560 16992
rect 21784 16952 22560 16980
rect 21784 16940 21790 16952
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 23290 16940 23296 16992
rect 23348 16940 23354 16992
rect 25314 16940 25320 16992
rect 25372 16980 25378 16992
rect 25958 16980 25964 16992
rect 25372 16952 25964 16980
rect 25372 16940 25378 16952
rect 25958 16940 25964 16952
rect 26016 16940 26022 16992
rect 27154 16940 27160 16992
rect 27212 16980 27218 16992
rect 29549 16983 29607 16989
rect 29549 16980 29561 16983
rect 27212 16952 29561 16980
rect 27212 16940 27218 16952
rect 29549 16949 29561 16952
rect 29595 16949 29607 16983
rect 30852 16980 30880 17020
rect 30926 17008 30932 17060
rect 30984 17048 30990 17060
rect 47394 17048 47400 17060
rect 30984 17020 47400 17048
rect 30984 17008 30990 17020
rect 47394 17008 47400 17020
rect 47452 17008 47458 17060
rect 47118 16980 47124 16992
rect 30852 16952 47124 16980
rect 29549 16943 29607 16949
rect 47118 16940 47124 16952
rect 47176 16940 47182 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 1762 16736 1768 16788
rect 1820 16776 1826 16788
rect 10870 16776 10876 16788
rect 1820 16748 10876 16776
rect 1820 16736 1826 16748
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 11698 16736 11704 16788
rect 11756 16776 11762 16788
rect 16850 16776 16856 16788
rect 11756 16748 16856 16776
rect 11756 16736 11762 16748
rect 16850 16736 16856 16748
rect 16908 16736 16914 16788
rect 17126 16736 17132 16788
rect 17184 16776 17190 16788
rect 19702 16776 19708 16788
rect 17184 16748 19708 16776
rect 17184 16736 17190 16748
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 19794 16736 19800 16788
rect 19852 16776 19858 16788
rect 20990 16776 20996 16788
rect 19852 16748 20996 16776
rect 19852 16736 19858 16748
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 23750 16736 23756 16788
rect 23808 16776 23814 16788
rect 30190 16776 30196 16788
rect 23808 16748 30196 16776
rect 23808 16736 23814 16748
rect 30190 16736 30196 16748
rect 30248 16736 30254 16788
rect 2130 16668 2136 16720
rect 2188 16708 2194 16720
rect 3421 16711 3479 16717
rect 3421 16708 3433 16711
rect 2188 16680 3433 16708
rect 2188 16668 2194 16680
rect 3421 16677 3433 16680
rect 3467 16708 3479 16711
rect 3510 16708 3516 16720
rect 3467 16680 3516 16708
rect 3467 16677 3479 16680
rect 3421 16671 3479 16677
rect 3510 16668 3516 16680
rect 3568 16668 3574 16720
rect 3605 16711 3663 16717
rect 3605 16677 3617 16711
rect 3651 16708 3663 16711
rect 4062 16708 4068 16720
rect 3651 16680 4068 16708
rect 3651 16677 3663 16680
rect 3605 16671 3663 16677
rect 4062 16668 4068 16680
rect 4120 16668 4126 16720
rect 5534 16668 5540 16720
rect 5592 16708 5598 16720
rect 6089 16711 6147 16717
rect 6089 16708 6101 16711
rect 5592 16680 6101 16708
rect 5592 16668 5598 16680
rect 6089 16677 6101 16680
rect 6135 16677 6147 16711
rect 9401 16711 9459 16717
rect 9401 16708 9413 16711
rect 6089 16671 6147 16677
rect 7208 16680 9413 16708
rect 2314 16600 2320 16652
rect 2372 16640 2378 16652
rect 3326 16640 3332 16652
rect 2372 16612 3332 16640
rect 2372 16600 2378 16612
rect 3326 16600 3332 16612
rect 3384 16600 3390 16652
rect 4522 16600 4528 16652
rect 4580 16600 4586 16652
rect 5718 16600 5724 16652
rect 5776 16640 5782 16652
rect 6270 16640 6276 16652
rect 5776 16612 6276 16640
rect 5776 16600 5782 16612
rect 6270 16600 6276 16612
rect 6328 16640 6334 16652
rect 7101 16643 7159 16649
rect 7101 16640 7113 16643
rect 6328 16612 7113 16640
rect 6328 16600 6334 16612
rect 7101 16609 7113 16612
rect 7147 16609 7159 16643
rect 7101 16603 7159 16609
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 1811 16544 2774 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 2746 16504 2774 16544
rect 3970 16532 3976 16584
rect 4028 16532 4034 16584
rect 7208 16572 7236 16680
rect 9401 16677 9413 16680
rect 9447 16677 9459 16711
rect 9401 16671 9459 16677
rect 9769 16711 9827 16717
rect 9769 16677 9781 16711
rect 9815 16708 9827 16711
rect 10410 16708 10416 16720
rect 9815 16680 10416 16708
rect 9815 16677 9827 16680
rect 9769 16671 9827 16677
rect 10410 16668 10416 16680
rect 10468 16668 10474 16720
rect 10704 16680 11928 16708
rect 10704 16649 10732 16680
rect 7285 16643 7343 16649
rect 7285 16609 7297 16643
rect 7331 16640 7343 16643
rect 8481 16643 8539 16649
rect 8481 16640 8493 16643
rect 7331 16612 8493 16640
rect 7331 16609 7343 16612
rect 7285 16603 7343 16609
rect 8481 16609 8493 16612
rect 8527 16640 8539 16643
rect 10689 16643 10747 16649
rect 10689 16640 10701 16643
rect 8527 16612 10701 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 10689 16609 10701 16612
rect 10735 16609 10747 16643
rect 10689 16603 10747 16609
rect 11606 16600 11612 16652
rect 11664 16640 11670 16652
rect 11900 16649 11928 16680
rect 12250 16668 12256 16720
rect 12308 16708 12314 16720
rect 12437 16711 12495 16717
rect 12437 16708 12449 16711
rect 12308 16680 12449 16708
rect 12308 16668 12314 16680
rect 12437 16677 12449 16680
rect 12483 16677 12495 16711
rect 12437 16671 12495 16677
rect 12986 16668 12992 16720
rect 13044 16668 13050 16720
rect 13262 16668 13268 16720
rect 13320 16708 13326 16720
rect 13538 16708 13544 16720
rect 13320 16680 13544 16708
rect 13320 16668 13326 16680
rect 13538 16668 13544 16680
rect 13596 16668 13602 16720
rect 18138 16708 18144 16720
rect 13648 16680 18144 16708
rect 11701 16643 11759 16649
rect 11701 16640 11713 16643
rect 11664 16612 11713 16640
rect 11664 16600 11670 16612
rect 11701 16609 11713 16612
rect 11747 16609 11759 16643
rect 11701 16603 11759 16609
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16640 11943 16643
rect 12342 16640 12348 16652
rect 11931 16612 12348 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 13648 16649 13676 16680
rect 18138 16668 18144 16680
rect 18196 16668 18202 16720
rect 21082 16668 21088 16720
rect 21140 16708 21146 16720
rect 21450 16708 21456 16720
rect 21140 16680 21456 16708
rect 21140 16668 21146 16680
rect 21450 16668 21456 16680
rect 21508 16668 21514 16720
rect 25130 16668 25136 16720
rect 25188 16708 25194 16720
rect 25188 16680 28488 16708
rect 25188 16668 25194 16680
rect 12713 16643 12771 16649
rect 12713 16640 12725 16643
rect 12584 16612 12725 16640
rect 12584 16600 12590 16612
rect 12713 16609 12725 16612
rect 12759 16640 12771 16643
rect 13449 16643 13507 16649
rect 13449 16640 13461 16643
rect 12759 16612 13461 16640
rect 12759 16609 12771 16612
rect 12713 16603 12771 16609
rect 13449 16609 13461 16612
rect 13495 16609 13507 16643
rect 13449 16603 13507 16609
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16609 13691 16643
rect 13633 16603 13691 16609
rect 14458 16600 14464 16652
rect 14516 16640 14522 16652
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 14516 16612 15485 16640
rect 14516 16600 14522 16612
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16640 15715 16643
rect 16298 16640 16304 16652
rect 15703 16612 16304 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 16761 16643 16819 16649
rect 16761 16609 16773 16643
rect 16807 16640 16819 16643
rect 17218 16640 17224 16652
rect 16807 16612 17224 16640
rect 16807 16609 16819 16612
rect 16761 16603 16819 16609
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 18506 16640 18512 16652
rect 18248 16612 18512 16640
rect 4080 16544 7236 16572
rect 4080 16504 4108 16544
rect 7742 16532 7748 16584
rect 7800 16572 7806 16584
rect 7800 16544 9076 16572
rect 7800 16532 7806 16544
rect 2746 16476 4108 16504
rect 2501 16467 2559 16473
rect 5902 16464 5908 16516
rect 5960 16464 5966 16516
rect 7009 16507 7067 16513
rect 7009 16473 7021 16507
rect 7055 16504 7067 16507
rect 7926 16504 7932 16516
rect 7055 16476 7932 16504
rect 7055 16473 7067 16476
rect 7009 16467 7067 16473
rect 7926 16464 7932 16476
rect 7984 16464 7990 16516
rect 8202 16464 8208 16516
rect 8260 16504 8266 16516
rect 8938 16504 8944 16516
rect 8260 16476 8944 16504
rect 8260 16464 8266 16476
rect 8938 16464 8944 16476
rect 8996 16464 9002 16516
rect 6641 16439 6699 16445
rect 6641 16405 6653 16439
rect 6687 16436 6699 16439
rect 6822 16436 6828 16448
rect 6687 16408 6828 16436
rect 6687 16405 6699 16408
rect 6641 16399 6699 16405
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 7834 16396 7840 16448
rect 7892 16396 7898 16448
rect 8110 16396 8116 16448
rect 8168 16436 8174 16448
rect 8297 16439 8355 16445
rect 8297 16436 8309 16439
rect 8168 16408 8309 16436
rect 8168 16396 8174 16408
rect 8297 16405 8309 16408
rect 8343 16405 8355 16439
rect 9048 16436 9076 16544
rect 10410 16532 10416 16584
rect 10468 16532 10474 16584
rect 10502 16532 10508 16584
rect 10560 16532 10566 16584
rect 14553 16575 14611 16581
rect 12728 16544 13492 16572
rect 9217 16507 9275 16513
rect 9217 16473 9229 16507
rect 9263 16504 9275 16507
rect 12728 16504 12756 16544
rect 9263 16476 12756 16504
rect 9263 16473 9275 16476
rect 9217 16467 9275 16473
rect 12802 16464 12808 16516
rect 12860 16504 12866 16516
rect 13357 16507 13415 16513
rect 13357 16504 13369 16507
rect 12860 16476 13369 16504
rect 12860 16464 12866 16476
rect 13357 16473 13369 16476
rect 13403 16473 13415 16507
rect 13464 16504 13492 16544
rect 14553 16541 14565 16575
rect 14599 16572 14611 16575
rect 14642 16572 14648 16584
rect 14599 16544 14648 16572
rect 14599 16541 14611 16544
rect 14553 16535 14611 16541
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 15378 16532 15384 16584
rect 15436 16532 15442 16584
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 15620 16544 15884 16572
rect 15620 16532 15626 16544
rect 13538 16504 13544 16516
rect 13464 16476 13544 16504
rect 13357 16467 13415 16473
rect 13538 16464 13544 16476
rect 13596 16464 13602 16516
rect 10045 16439 10103 16445
rect 10045 16436 10057 16439
rect 9048 16408 10057 16436
rect 8297 16399 8355 16405
rect 10045 16405 10057 16408
rect 10091 16405 10103 16439
rect 10045 16399 10103 16405
rect 11238 16396 11244 16448
rect 11296 16396 11302 16448
rect 11609 16439 11667 16445
rect 11609 16405 11621 16439
rect 11655 16436 11667 16439
rect 11882 16436 11888 16448
rect 11655 16408 11888 16436
rect 11655 16405 11667 16408
rect 11609 16399 11667 16405
rect 11882 16396 11888 16408
rect 11940 16436 11946 16448
rect 12253 16439 12311 16445
rect 12253 16436 12265 16439
rect 11940 16408 12265 16436
rect 11940 16396 11946 16408
rect 12253 16405 12265 16408
rect 12299 16405 12311 16439
rect 12253 16399 12311 16405
rect 14366 16396 14372 16448
rect 14424 16396 14430 16448
rect 15013 16439 15071 16445
rect 15013 16405 15025 16439
rect 15059 16436 15071 16439
rect 15562 16436 15568 16448
rect 15059 16408 15568 16436
rect 15059 16405 15071 16408
rect 15013 16399 15071 16405
rect 15562 16396 15568 16408
rect 15620 16396 15626 16448
rect 15856 16436 15884 16544
rect 15930 16532 15936 16584
rect 15988 16572 15994 16584
rect 18248 16581 18276 16612
rect 18506 16600 18512 16612
rect 18564 16600 18570 16652
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 20346 16640 20352 16652
rect 19751 16612 20352 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 20346 16600 20352 16612
rect 20404 16600 20410 16652
rect 20714 16600 20720 16652
rect 20772 16640 20778 16652
rect 22465 16643 22523 16649
rect 22465 16640 22477 16643
rect 20772 16612 22477 16640
rect 20772 16600 20778 16612
rect 22465 16609 22477 16612
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 22554 16600 22560 16652
rect 22612 16600 22618 16652
rect 23750 16600 23756 16652
rect 23808 16600 23814 16652
rect 24578 16600 24584 16652
rect 24636 16640 24642 16652
rect 25222 16640 25228 16652
rect 24636 16612 25228 16640
rect 24636 16600 24642 16612
rect 25222 16600 25228 16612
rect 25280 16600 25286 16652
rect 25317 16643 25375 16649
rect 25317 16609 25329 16643
rect 25363 16640 25375 16643
rect 25774 16640 25780 16652
rect 25363 16612 25780 16640
rect 25363 16609 25375 16612
rect 25317 16603 25375 16609
rect 25774 16600 25780 16612
rect 25832 16600 25838 16652
rect 25958 16600 25964 16652
rect 26016 16600 26022 16652
rect 27062 16600 27068 16652
rect 27120 16600 27126 16652
rect 27154 16600 27160 16652
rect 27212 16600 27218 16652
rect 28460 16649 28488 16680
rect 28445 16643 28503 16649
rect 28445 16609 28457 16643
rect 28491 16640 28503 16643
rect 28718 16640 28724 16652
rect 28491 16612 28724 16640
rect 28491 16609 28503 16612
rect 28445 16603 28503 16609
rect 28718 16600 28724 16612
rect 28776 16600 28782 16652
rect 30834 16640 30840 16652
rect 28920 16612 30840 16640
rect 16209 16575 16267 16581
rect 16209 16572 16221 16575
rect 15988 16544 16221 16572
rect 15988 16532 15994 16544
rect 16209 16541 16221 16544
rect 16255 16541 16267 16575
rect 16209 16535 16267 16541
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 18233 16575 18291 16581
rect 18233 16541 18245 16575
rect 18279 16541 18291 16575
rect 18233 16535 18291 16541
rect 17604 16504 17632 16535
rect 18322 16532 18328 16584
rect 18380 16572 18386 16584
rect 19150 16572 19156 16584
rect 18380 16544 19156 16572
rect 18380 16532 18386 16544
rect 19150 16532 19156 16544
rect 19208 16532 19214 16584
rect 19426 16532 19432 16584
rect 19484 16532 19490 16584
rect 22373 16575 22431 16581
rect 22373 16541 22385 16575
rect 22419 16572 22431 16575
rect 23290 16572 23296 16584
rect 22419 16544 23296 16572
rect 22419 16541 22431 16544
rect 22373 16535 22431 16541
rect 23290 16532 23296 16544
rect 23348 16532 23354 16584
rect 23569 16575 23627 16581
rect 23569 16541 23581 16575
rect 23615 16572 23627 16575
rect 23658 16572 23664 16584
rect 23615 16544 23664 16572
rect 23615 16541 23627 16544
rect 23569 16535 23627 16541
rect 23658 16532 23664 16544
rect 23716 16572 23722 16584
rect 24486 16572 24492 16584
rect 23716 16544 24492 16572
rect 23716 16532 23722 16544
rect 24486 16532 24492 16544
rect 24544 16532 24550 16584
rect 25038 16532 25044 16584
rect 25096 16572 25102 16584
rect 25096 16544 26740 16572
rect 25096 16532 25102 16544
rect 20990 16504 20996 16516
rect 17604 16476 20024 16504
rect 20930 16476 20996 16504
rect 16025 16439 16083 16445
rect 16025 16436 16037 16439
rect 15856 16408 16037 16436
rect 16025 16405 16037 16408
rect 16071 16405 16083 16439
rect 16025 16399 16083 16405
rect 16390 16396 16396 16448
rect 16448 16396 16454 16448
rect 16850 16396 16856 16448
rect 16908 16436 16914 16448
rect 17405 16439 17463 16445
rect 17405 16436 17417 16439
rect 16908 16408 17417 16436
rect 16908 16396 16914 16408
rect 17405 16405 17417 16408
rect 17451 16405 17463 16439
rect 17405 16399 17463 16405
rect 18049 16439 18107 16445
rect 18049 16405 18061 16439
rect 18095 16436 18107 16439
rect 18322 16436 18328 16448
rect 18095 16408 18328 16436
rect 18095 16405 18107 16408
rect 18049 16399 18107 16405
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 18598 16396 18604 16448
rect 18656 16436 18662 16448
rect 18693 16439 18751 16445
rect 18693 16436 18705 16439
rect 18656 16408 18705 16436
rect 18656 16396 18662 16408
rect 18693 16405 18705 16408
rect 18739 16405 18751 16439
rect 19996 16436 20024 16476
rect 20990 16464 20996 16476
rect 21048 16464 21054 16516
rect 21174 16464 21180 16516
rect 21232 16504 21238 16516
rect 21453 16507 21511 16513
rect 21453 16504 21465 16507
rect 21232 16476 21465 16504
rect 21232 16464 21238 16476
rect 21453 16473 21465 16476
rect 21499 16473 21511 16507
rect 25314 16504 25320 16516
rect 21453 16467 21511 16473
rect 25056 16476 25320 16504
rect 20070 16436 20076 16448
rect 19996 16408 20076 16436
rect 18693 16399 18751 16405
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20714 16396 20720 16448
rect 20772 16436 20778 16448
rect 22005 16439 22063 16445
rect 22005 16436 22017 16439
rect 20772 16408 22017 16436
rect 20772 16396 20778 16408
rect 22005 16405 22017 16408
rect 22051 16405 22063 16439
rect 22005 16399 22063 16405
rect 22370 16396 22376 16448
rect 22428 16436 22434 16448
rect 23201 16439 23259 16445
rect 23201 16436 23213 16439
rect 22428 16408 23213 16436
rect 22428 16396 22434 16408
rect 23201 16405 23213 16408
rect 23247 16405 23259 16439
rect 23201 16399 23259 16405
rect 23661 16439 23719 16445
rect 23661 16405 23673 16439
rect 23707 16436 23719 16439
rect 23842 16436 23848 16448
rect 23707 16408 23848 16436
rect 23707 16405 23719 16408
rect 23661 16399 23719 16405
rect 23842 16396 23848 16408
rect 23900 16436 23906 16448
rect 24578 16436 24584 16448
rect 23900 16408 24584 16436
rect 23900 16396 23906 16408
rect 24578 16396 24584 16408
rect 24636 16396 24642 16448
rect 24670 16396 24676 16448
rect 24728 16396 24734 16448
rect 25056 16445 25084 16476
rect 25314 16464 25320 16476
rect 25372 16464 25378 16516
rect 25498 16464 25504 16516
rect 25556 16504 25562 16516
rect 25556 16476 26648 16504
rect 25556 16464 25562 16476
rect 25041 16439 25099 16445
rect 25041 16405 25053 16439
rect 25087 16405 25099 16439
rect 25041 16399 25099 16405
rect 25130 16396 25136 16448
rect 25188 16436 25194 16448
rect 25682 16436 25688 16448
rect 25188 16408 25688 16436
rect 25188 16396 25194 16408
rect 25682 16396 25688 16408
rect 25740 16396 25746 16448
rect 26620 16445 26648 16476
rect 26605 16439 26663 16445
rect 26605 16405 26617 16439
rect 26651 16405 26663 16439
rect 26712 16436 26740 16544
rect 27614 16532 27620 16584
rect 27672 16572 27678 16584
rect 28169 16575 28227 16581
rect 28169 16572 28181 16575
rect 27672 16544 28181 16572
rect 27672 16532 27678 16544
rect 28169 16541 28181 16544
rect 28215 16541 28227 16575
rect 28169 16535 28227 16541
rect 28261 16575 28319 16581
rect 28261 16541 28273 16575
rect 28307 16572 28319 16575
rect 28350 16572 28356 16584
rect 28307 16544 28356 16572
rect 28307 16541 28319 16544
rect 28261 16535 28319 16541
rect 28350 16532 28356 16544
rect 28408 16572 28414 16584
rect 28920 16572 28948 16612
rect 30834 16600 30840 16612
rect 30892 16600 30898 16652
rect 28408 16544 28948 16572
rect 28408 16532 28414 16544
rect 26973 16507 27031 16513
rect 26973 16473 26985 16507
rect 27019 16504 27031 16507
rect 28442 16504 28448 16516
rect 27019 16476 28448 16504
rect 27019 16473 27031 16476
rect 26973 16467 27031 16473
rect 28442 16464 28448 16476
rect 28500 16464 28506 16516
rect 27801 16439 27859 16445
rect 27801 16436 27813 16439
rect 26712 16408 27813 16436
rect 26605 16399 26663 16405
rect 27801 16405 27813 16408
rect 27847 16405 27859 16439
rect 27801 16399 27859 16405
rect 28258 16396 28264 16448
rect 28316 16436 28322 16448
rect 28534 16436 28540 16448
rect 28316 16408 28540 16436
rect 28316 16396 28322 16408
rect 28534 16396 28540 16408
rect 28592 16396 28598 16448
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 3970 16192 3976 16244
rect 4028 16232 4034 16244
rect 6914 16232 6920 16244
rect 4028 16204 6920 16232
rect 4028 16192 4034 16204
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 7006 16192 7012 16244
rect 7064 16232 7070 16244
rect 7285 16235 7343 16241
rect 7285 16232 7297 16235
rect 7064 16204 7297 16232
rect 7064 16192 7070 16204
rect 7285 16201 7297 16204
rect 7331 16201 7343 16235
rect 10229 16235 10287 16241
rect 7285 16195 7343 16201
rect 7392 16204 10088 16232
rect 4246 16124 4252 16176
rect 4304 16164 4310 16176
rect 4341 16167 4399 16173
rect 4341 16164 4353 16167
rect 4304 16136 4353 16164
rect 4304 16124 4310 16136
rect 4341 16133 4353 16136
rect 4387 16133 4399 16167
rect 4341 16127 4399 16133
rect 5718 16124 5724 16176
rect 5776 16124 5782 16176
rect 5810 16124 5816 16176
rect 5868 16164 5874 16176
rect 7392 16164 7420 16204
rect 5868 16136 7420 16164
rect 5868 16124 5874 16136
rect 9766 16124 9772 16176
rect 9824 16124 9830 16176
rect 10060 16164 10088 16204
rect 10229 16201 10241 16235
rect 10275 16232 10287 16235
rect 10502 16232 10508 16244
rect 10275 16204 10508 16232
rect 10275 16201 10287 16204
rect 10229 16195 10287 16201
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 10594 16192 10600 16244
rect 10652 16192 10658 16244
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 11514 16232 11520 16244
rect 11204 16204 11520 16232
rect 11204 16192 11210 16204
rect 11514 16192 11520 16204
rect 11572 16232 11578 16244
rect 11609 16235 11667 16241
rect 11609 16232 11621 16235
rect 11572 16204 11621 16232
rect 11572 16192 11578 16204
rect 11609 16201 11621 16204
rect 11655 16201 11667 16235
rect 11609 16195 11667 16201
rect 13630 16192 13636 16244
rect 13688 16232 13694 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 13688 16204 13737 16232
rect 13688 16192 13694 16204
rect 13725 16201 13737 16204
rect 13771 16201 13783 16235
rect 13725 16195 13783 16201
rect 14568 16204 16620 16232
rect 12526 16164 12532 16176
rect 10060 16136 12532 16164
rect 12526 16124 12532 16136
rect 12584 16124 12590 16176
rect 13998 16164 14004 16176
rect 13478 16136 14004 16164
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 1811 16068 2774 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2746 16028 2774 16068
rect 3510 16056 3516 16108
rect 3568 16056 3574 16108
rect 3694 16056 3700 16108
rect 3752 16096 3758 16108
rect 5629 16099 5687 16105
rect 5629 16096 5641 16099
rect 3752 16068 5641 16096
rect 3752 16056 3758 16068
rect 5629 16065 5641 16068
rect 5675 16065 5687 16099
rect 5629 16059 5687 16065
rect 7282 16056 7288 16108
rect 7340 16096 7346 16108
rect 7653 16099 7711 16105
rect 7653 16096 7665 16099
rect 7340 16068 7665 16096
rect 7340 16056 7346 16068
rect 7653 16065 7665 16068
rect 7699 16065 7711 16099
rect 7653 16059 7711 16065
rect 8478 16056 8484 16108
rect 8536 16056 8542 16108
rect 11149 16099 11207 16105
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11195 16068 11928 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 4706 16028 4712 16040
rect 2746 16000 4712 16028
rect 2041 15991 2099 15997
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 16028 5963 16031
rect 5994 16028 6000 16040
rect 5951 16000 6000 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 5994 15988 6000 16000
rect 6052 16028 6058 16040
rect 6546 16028 6552 16040
rect 6052 16000 6552 16028
rect 6052 15988 6058 16000
rect 6546 15988 6552 16000
rect 6604 15988 6610 16040
rect 6638 15988 6644 16040
rect 6696 15988 6702 16040
rect 7374 15988 7380 16040
rect 7432 16028 7438 16040
rect 7745 16031 7803 16037
rect 7745 16028 7757 16031
rect 7432 16000 7757 16028
rect 7432 15988 7438 16000
rect 7745 15997 7757 16000
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 7926 15988 7932 16040
rect 7984 15988 7990 16040
rect 8757 16031 8815 16037
rect 8757 16028 8769 16031
rect 8588 16000 8769 16028
rect 6362 15920 6368 15972
rect 6420 15960 6426 15972
rect 8478 15960 8484 15972
rect 6420 15932 8484 15960
rect 6420 15920 6426 15932
rect 8478 15920 8484 15932
rect 8536 15960 8542 15972
rect 8588 15960 8616 16000
rect 8757 15997 8769 16000
rect 8803 16028 8815 16031
rect 9950 16028 9956 16040
rect 8803 16000 9956 16028
rect 8803 15997 8815 16000
rect 8757 15991 8815 15997
rect 9950 15988 9956 16000
rect 10008 16028 10014 16040
rect 10134 16028 10140 16040
rect 10008 16000 10140 16028
rect 10008 15988 10014 16000
rect 10134 15988 10140 16000
rect 10192 16028 10198 16040
rect 10870 16028 10876 16040
rect 10192 16000 10876 16028
rect 10192 15988 10198 16000
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 8536 15932 8616 15960
rect 8536 15920 8542 15932
rect 10962 15920 10968 15972
rect 11020 15920 11026 15972
rect 5258 15852 5264 15904
rect 5316 15852 5322 15904
rect 7006 15852 7012 15904
rect 7064 15892 7070 15904
rect 11790 15892 11796 15904
rect 7064 15864 11796 15892
rect 7064 15852 7070 15864
rect 11790 15852 11796 15864
rect 11848 15852 11854 15904
rect 11900 15892 11928 16068
rect 11974 16056 11980 16108
rect 12032 16056 12038 16108
rect 12250 15988 12256 16040
rect 12308 15988 12314 16040
rect 12342 15988 12348 16040
rect 12400 16028 12406 16040
rect 14568 16028 14596 16204
rect 14645 16167 14703 16173
rect 14645 16133 14657 16167
rect 14691 16164 14703 16167
rect 16482 16164 16488 16176
rect 14691 16136 16488 16164
rect 14691 16133 14703 16136
rect 14645 16127 14703 16133
rect 16482 16124 16488 16136
rect 16540 16124 16546 16176
rect 16592 16164 16620 16204
rect 16666 16192 16672 16244
rect 16724 16232 16730 16244
rect 16942 16232 16948 16244
rect 16724 16204 16948 16232
rect 16724 16192 16730 16204
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 17126 16192 17132 16244
rect 17184 16192 17190 16244
rect 17405 16235 17463 16241
rect 17405 16201 17417 16235
rect 17451 16232 17463 16235
rect 17494 16232 17500 16244
rect 17451 16204 17500 16232
rect 17451 16201 17463 16204
rect 17405 16195 17463 16201
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 17862 16192 17868 16244
rect 17920 16192 17926 16244
rect 19702 16192 19708 16244
rect 19760 16232 19766 16244
rect 20533 16235 20591 16241
rect 20533 16232 20545 16235
rect 19760 16204 20545 16232
rect 19760 16192 19766 16204
rect 20533 16201 20545 16204
rect 20579 16201 20591 16235
rect 21174 16232 21180 16244
rect 20533 16195 20591 16201
rect 20640 16204 21180 16232
rect 20640 16164 20668 16204
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 24946 16192 24952 16244
rect 25004 16232 25010 16244
rect 26605 16235 26663 16241
rect 26605 16232 26617 16235
rect 25004 16204 26617 16232
rect 25004 16192 25010 16204
rect 26605 16201 26617 16204
rect 26651 16201 26663 16235
rect 26605 16195 26663 16201
rect 26970 16192 26976 16244
rect 27028 16192 27034 16244
rect 27614 16192 27620 16244
rect 27672 16232 27678 16244
rect 27709 16235 27767 16241
rect 27709 16232 27721 16235
rect 27672 16204 27721 16232
rect 27672 16192 27678 16204
rect 27709 16201 27721 16204
rect 27755 16232 27767 16235
rect 28350 16232 28356 16244
rect 27755 16204 28356 16232
rect 27755 16201 27767 16204
rect 27709 16195 27767 16201
rect 28350 16192 28356 16204
rect 28408 16192 28414 16244
rect 24397 16167 24455 16173
rect 16592 16136 20668 16164
rect 21560 16136 24348 16164
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16096 14795 16099
rect 15010 16096 15016 16108
rect 14783 16068 15016 16096
rect 14783 16065 14795 16068
rect 14737 16059 14795 16065
rect 15010 16056 15016 16068
rect 15068 16096 15074 16108
rect 16301 16099 16359 16105
rect 15068 16068 15608 16096
rect 15068 16056 15074 16068
rect 12400 16000 14596 16028
rect 14829 16031 14887 16037
rect 12400 15988 12406 16000
rect 14829 15997 14841 16031
rect 14875 15997 14887 16031
rect 14829 15991 14887 15997
rect 13630 15920 13636 15972
rect 13688 15960 13694 15972
rect 14844 15960 14872 15991
rect 14918 15988 14924 16040
rect 14976 15988 14982 16040
rect 15470 15988 15476 16040
rect 15528 15988 15534 16040
rect 15580 16028 15608 16068
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 17586 16096 17592 16108
rect 16347 16068 17592 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 17586 16056 17592 16068
rect 17644 16056 17650 16108
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16065 17831 16099
rect 17773 16059 17831 16065
rect 16574 16028 16580 16040
rect 15580 16000 16580 16028
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 16666 15988 16672 16040
rect 16724 16028 16730 16040
rect 17788 16028 17816 16059
rect 17862 16056 17868 16108
rect 17920 16096 17926 16108
rect 18601 16099 18659 16105
rect 17920 16068 18552 16096
rect 17920 16056 17926 16068
rect 17957 16031 18015 16037
rect 17957 16028 17969 16031
rect 16724 16000 17816 16028
rect 17880 16000 17969 16028
rect 16724 15988 16730 16000
rect 13688 15932 14872 15960
rect 14936 15960 14964 15988
rect 14936 15932 17540 15960
rect 13688 15920 13694 15932
rect 12434 15892 12440 15904
rect 11900 15864 12440 15892
rect 12434 15852 12440 15864
rect 12492 15852 12498 15904
rect 13722 15852 13728 15904
rect 13780 15892 13786 15904
rect 14277 15895 14335 15901
rect 14277 15892 14289 15895
rect 13780 15864 14289 15892
rect 13780 15852 13786 15864
rect 14277 15861 14289 15864
rect 14323 15861 14335 15895
rect 14277 15855 14335 15861
rect 14918 15852 14924 15904
rect 14976 15892 14982 15904
rect 16117 15895 16175 15901
rect 16117 15892 16129 15895
rect 14976 15864 16129 15892
rect 14976 15852 14982 15864
rect 16117 15861 16129 15864
rect 16163 15861 16175 15895
rect 16117 15855 16175 15861
rect 16390 15852 16396 15904
rect 16448 15892 16454 15904
rect 16574 15892 16580 15904
rect 16448 15864 16580 15892
rect 16448 15852 16454 15864
rect 16574 15852 16580 15864
rect 16632 15892 16638 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 16632 15864 16681 15892
rect 16632 15852 16638 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 17512 15892 17540 15932
rect 17586 15920 17592 15972
rect 17644 15960 17650 15972
rect 17880 15960 17908 16000
rect 17957 15997 17969 16000
rect 18003 15997 18015 16031
rect 17957 15991 18015 15997
rect 17644 15932 17908 15960
rect 18524 15960 18552 16068
rect 18601 16065 18613 16099
rect 18647 16096 18659 16099
rect 18690 16096 18696 16108
rect 18647 16068 18696 16096
rect 18647 16065 18659 16068
rect 18601 16059 18659 16065
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 18874 16056 18880 16108
rect 18932 16056 18938 16108
rect 20438 16056 20444 16108
rect 20496 16056 20502 16108
rect 21450 16056 21456 16108
rect 21508 16056 21514 16108
rect 20717 16031 20775 16037
rect 20717 15997 20729 16031
rect 20763 16028 20775 16031
rect 21560 16028 21588 16136
rect 23658 16056 23664 16108
rect 23716 16056 23722 16108
rect 23753 16099 23811 16105
rect 23753 16065 23765 16099
rect 23799 16096 23811 16099
rect 23842 16096 23848 16108
rect 23799 16068 23848 16096
rect 23799 16065 23811 16068
rect 23753 16059 23811 16065
rect 23842 16056 23848 16068
rect 23900 16056 23906 16108
rect 20763 16000 21588 16028
rect 20763 15997 20775 16000
rect 20717 15991 20775 15997
rect 21634 15988 21640 16040
rect 21692 16028 21698 16040
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 21692 16000 22017 16028
rect 21692 15988 21698 16000
rect 22005 15997 22017 16000
rect 22051 15997 22063 16031
rect 22005 15991 22063 15997
rect 22278 15988 22284 16040
rect 22336 15988 22342 16040
rect 23937 16031 23995 16037
rect 23937 15997 23949 16031
rect 23983 16028 23995 16031
rect 24026 16028 24032 16040
rect 23983 16000 24032 16028
rect 23983 15997 23995 16000
rect 23937 15991 23995 15997
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 24320 16028 24348 16136
rect 24397 16133 24409 16167
rect 24443 16164 24455 16167
rect 24486 16164 24492 16176
rect 24443 16136 24492 16164
rect 24443 16133 24455 16136
rect 24397 16127 24455 16133
rect 24486 16124 24492 16136
rect 24544 16124 24550 16176
rect 24578 16124 24584 16176
rect 24636 16124 24642 16176
rect 26988 16164 27016 16192
rect 26358 16136 27016 16164
rect 24854 16056 24860 16108
rect 24912 16056 24918 16108
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24320 16000 25145 16028
rect 25133 15997 25145 16000
rect 25179 16028 25191 16031
rect 27154 16028 27160 16040
rect 25179 16000 27160 16028
rect 25179 15997 25191 16000
rect 25133 15991 25191 15997
rect 27154 15988 27160 16000
rect 27212 15988 27218 16040
rect 20073 15963 20131 15969
rect 18524 15932 19334 15960
rect 17644 15920 17650 15932
rect 18598 15892 18604 15904
rect 17512 15864 18604 15892
rect 16669 15855 16727 15861
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 19306 15892 19334 15932
rect 20073 15929 20085 15963
rect 20119 15960 20131 15963
rect 23382 15960 23388 15972
rect 20119 15932 23388 15960
rect 20119 15929 20131 15932
rect 20073 15923 20131 15929
rect 23382 15920 23388 15932
rect 23440 15920 23446 15972
rect 21269 15895 21327 15901
rect 21269 15892 21281 15895
rect 19306 15864 21281 15892
rect 21269 15861 21281 15864
rect 21315 15861 21327 15895
rect 21269 15855 21327 15861
rect 22462 15852 22468 15904
rect 22520 15892 22526 15904
rect 23293 15895 23351 15901
rect 23293 15892 23305 15895
rect 22520 15864 23305 15892
rect 22520 15852 22526 15864
rect 23293 15861 23305 15864
rect 23339 15861 23351 15895
rect 23293 15855 23351 15861
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 5810 15688 5816 15700
rect 4540 15660 5816 15688
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 1360 15524 2053 15552
rect 1360 15512 1366 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 3878 15512 3884 15564
rect 3936 15552 3942 15564
rect 4433 15555 4491 15561
rect 4433 15552 4445 15555
rect 3936 15524 4445 15552
rect 3936 15512 3942 15524
rect 4433 15521 4445 15524
rect 4479 15552 4491 15555
rect 4540 15552 4568 15660
rect 5810 15648 5816 15660
rect 5868 15648 5874 15700
rect 7190 15648 7196 15700
rect 7248 15688 7254 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7248 15660 7849 15688
rect 7248 15648 7254 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 7926 15648 7932 15700
rect 7984 15688 7990 15700
rect 8570 15688 8576 15700
rect 7984 15660 8576 15688
rect 7984 15648 7990 15660
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 8662 15648 8668 15700
rect 8720 15688 8726 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 8720 15660 9321 15688
rect 8720 15648 8726 15660
rect 9309 15657 9321 15660
rect 9355 15657 9367 15691
rect 12802 15688 12808 15700
rect 9309 15651 9367 15657
rect 10244 15660 12808 15688
rect 5994 15620 6000 15632
rect 4632 15592 6000 15620
rect 4632 15561 4660 15592
rect 5994 15580 6000 15592
rect 6052 15580 6058 15632
rect 7006 15620 7012 15632
rect 6656 15592 7012 15620
rect 4479 15524 4568 15552
rect 4617 15555 4675 15561
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 4617 15521 4629 15555
rect 4663 15521 4675 15555
rect 4617 15515 4675 15521
rect 5166 15512 5172 15564
rect 5224 15552 5230 15564
rect 5629 15555 5687 15561
rect 5629 15552 5641 15555
rect 5224 15524 5641 15552
rect 5224 15512 5230 15524
rect 5629 15521 5641 15524
rect 5675 15521 5687 15555
rect 5629 15515 5687 15521
rect 5813 15555 5871 15561
rect 5813 15521 5825 15555
rect 5859 15552 5871 15555
rect 6656 15552 6684 15592
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 7469 15623 7527 15629
rect 7469 15589 7481 15623
rect 7515 15620 7527 15623
rect 8294 15620 8300 15632
rect 7515 15592 8300 15620
rect 7515 15589 7527 15592
rect 7469 15583 7527 15589
rect 8294 15580 8300 15592
rect 8352 15620 8358 15632
rect 9214 15620 9220 15632
rect 8352 15592 9220 15620
rect 8352 15580 8358 15592
rect 9214 15580 9220 15592
rect 9272 15580 9278 15632
rect 5859 15524 6684 15552
rect 5859 15521 5871 15524
rect 5813 15515 5871 15521
rect 6730 15512 6736 15564
rect 6788 15552 6794 15564
rect 6825 15555 6883 15561
rect 6825 15552 6837 15555
rect 6788 15524 6837 15552
rect 6788 15512 6794 15524
rect 6825 15521 6837 15524
rect 6871 15521 6883 15555
rect 6825 15515 6883 15521
rect 6914 15512 6920 15564
rect 6972 15512 6978 15564
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 7156 15524 8156 15552
rect 7156 15512 7162 15524
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 3418 15484 3424 15496
rect 1811 15456 3424 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 3896 15456 6500 15484
rect 2774 15376 2780 15428
rect 2832 15416 2838 15428
rect 3329 15419 3387 15425
rect 3329 15416 3341 15419
rect 2832 15388 3341 15416
rect 2832 15376 2838 15388
rect 3329 15385 3341 15388
rect 3375 15416 3387 15419
rect 3896 15416 3924 15456
rect 5537 15419 5595 15425
rect 5537 15416 5549 15419
rect 3375 15388 3924 15416
rect 3988 15388 5549 15416
rect 3375 15385 3387 15388
rect 3329 15379 3387 15385
rect 3605 15351 3663 15357
rect 3605 15317 3617 15351
rect 3651 15348 3663 15351
rect 3786 15348 3792 15360
rect 3651 15320 3792 15348
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 3786 15308 3792 15320
rect 3844 15308 3850 15360
rect 3988 15357 4016 15388
rect 5537 15385 5549 15388
rect 5583 15385 5595 15419
rect 5537 15379 5595 15385
rect 3973 15351 4031 15357
rect 3973 15317 3985 15351
rect 4019 15317 4031 15351
rect 3973 15311 4031 15317
rect 4338 15308 4344 15360
rect 4396 15308 4402 15360
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 5718 15348 5724 15360
rect 5215 15320 5724 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 6362 15308 6368 15360
rect 6420 15308 6426 15360
rect 6472 15348 6500 15456
rect 6638 15444 6644 15496
rect 6696 15484 6702 15496
rect 8018 15484 8024 15496
rect 6696 15456 8024 15484
rect 6696 15444 6702 15456
rect 8018 15444 8024 15456
rect 8076 15444 8082 15496
rect 6733 15419 6791 15425
rect 6733 15385 6745 15419
rect 6779 15416 6791 15419
rect 7926 15416 7932 15428
rect 6779 15388 7932 15416
rect 6779 15385 6791 15388
rect 6733 15379 6791 15385
rect 7926 15376 7932 15388
rect 7984 15376 7990 15428
rect 8128 15416 8156 15524
rect 8202 15512 8208 15564
rect 8260 15552 8266 15564
rect 8260 15524 8432 15552
rect 8260 15512 8266 15524
rect 8404 15484 8432 15524
rect 8478 15512 8484 15564
rect 8536 15512 8542 15564
rect 10244 15561 10272 15660
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 13538 15648 13544 15700
rect 13596 15648 13602 15700
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 15470 15688 15476 15700
rect 14884 15660 15476 15688
rect 14884 15648 14890 15660
rect 15470 15648 15476 15660
rect 15528 15648 15534 15700
rect 15838 15648 15844 15700
rect 15896 15648 15902 15700
rect 19889 15691 19947 15697
rect 19889 15688 19901 15691
rect 16132 15660 19901 15688
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 16132 15620 16160 15660
rect 19889 15657 19901 15660
rect 19935 15657 19947 15691
rect 19889 15651 19947 15657
rect 20070 15648 20076 15700
rect 20128 15688 20134 15700
rect 20128 15660 21588 15688
rect 20128 15648 20134 15660
rect 19610 15620 19616 15632
rect 10744 15592 16160 15620
rect 16316 15592 16601 15620
rect 10744 15580 10750 15592
rect 10229 15555 10287 15561
rect 10229 15521 10241 15555
rect 10275 15521 10287 15555
rect 10229 15515 10287 15521
rect 10870 15512 10876 15564
rect 10928 15552 10934 15564
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 10928 15524 11437 15552
rect 10928 15512 10934 15524
rect 11425 15521 11437 15524
rect 11471 15521 11483 15555
rect 11425 15515 11483 15521
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 13354 15552 13360 15564
rect 12759 15524 13360 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 13354 15512 13360 15524
rect 13412 15512 13418 15564
rect 14550 15512 14556 15564
rect 14608 15552 14614 15564
rect 14921 15555 14979 15561
rect 14921 15552 14933 15555
rect 14608 15524 14933 15552
rect 14608 15512 14614 15524
rect 14921 15521 14933 15524
rect 14967 15521 14979 15555
rect 14921 15515 14979 15521
rect 15105 15555 15163 15561
rect 15105 15521 15117 15555
rect 15151 15521 15163 15555
rect 15105 15515 15163 15521
rect 8404 15456 9536 15484
rect 8205 15419 8263 15425
rect 8205 15416 8217 15419
rect 8128 15388 8217 15416
rect 8205 15385 8217 15388
rect 8251 15385 8263 15419
rect 8205 15379 8263 15385
rect 9214 15376 9220 15428
rect 9272 15376 9278 15428
rect 9508 15416 9536 15456
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 9916 15456 11345 15484
rect 9916 15444 9922 15456
rect 11333 15453 11345 15456
rect 11379 15484 11391 15487
rect 11514 15484 11520 15496
rect 11379 15456 11520 15484
rect 11379 15453 11391 15456
rect 11333 15447 11391 15453
rect 11514 15444 11520 15456
rect 11572 15444 11578 15496
rect 11790 15444 11796 15496
rect 11848 15484 11854 15496
rect 13630 15484 13636 15496
rect 11848 15456 13636 15484
rect 11848 15444 11854 15456
rect 13630 15444 13636 15456
rect 13688 15444 13694 15496
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 12437 15419 12495 15425
rect 12437 15416 12449 15419
rect 9508 15388 12449 15416
rect 12437 15385 12449 15388
rect 12483 15385 12495 15419
rect 12437 15379 12495 15385
rect 13265 15419 13323 15425
rect 13265 15385 13277 15419
rect 13311 15416 13323 15419
rect 13740 15416 13768 15447
rect 14826 15444 14832 15496
rect 14884 15444 14890 15496
rect 13311 15388 14964 15416
rect 13311 15385 13323 15388
rect 13265 15379 13323 15385
rect 8297 15351 8355 15357
rect 8297 15348 8309 15351
rect 6472 15320 8309 15348
rect 8297 15317 8309 15320
rect 8343 15317 8355 15351
rect 8297 15311 8355 15317
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 9306 15348 9312 15360
rect 8996 15320 9312 15348
rect 8996 15308 9002 15320
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 9766 15308 9772 15360
rect 9824 15308 9830 15360
rect 9858 15308 9864 15360
rect 9916 15308 9922 15360
rect 10318 15308 10324 15360
rect 10376 15348 10382 15360
rect 10686 15348 10692 15360
rect 10376 15320 10692 15348
rect 10376 15308 10382 15320
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 10870 15308 10876 15360
rect 10928 15308 10934 15360
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 11241 15351 11299 15357
rect 11241 15348 11253 15351
rect 11204 15320 11253 15348
rect 11204 15308 11210 15320
rect 11241 15317 11253 15320
rect 11287 15317 11299 15351
rect 11241 15311 11299 15317
rect 12066 15308 12072 15360
rect 12124 15308 12130 15360
rect 12526 15308 12532 15360
rect 12584 15308 12590 15360
rect 13998 15308 14004 15360
rect 14056 15348 14062 15360
rect 14093 15351 14151 15357
rect 14093 15348 14105 15351
rect 14056 15320 14105 15348
rect 14056 15308 14062 15320
rect 14093 15317 14105 15320
rect 14139 15317 14151 15351
rect 14093 15311 14151 15317
rect 14366 15308 14372 15360
rect 14424 15348 14430 15360
rect 14461 15351 14519 15357
rect 14461 15348 14473 15351
rect 14424 15320 14473 15348
rect 14424 15308 14430 15320
rect 14461 15317 14473 15320
rect 14507 15317 14519 15351
rect 14936 15348 14964 15388
rect 15010 15376 15016 15428
rect 15068 15416 15074 15428
rect 15120 15416 15148 15515
rect 16316 15484 16344 15592
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15521 16543 15555
rect 16573 15552 16601 15592
rect 18340 15592 19616 15620
rect 18340 15552 18368 15592
rect 19610 15580 19616 15592
rect 19668 15580 19674 15632
rect 21560 15620 21588 15660
rect 21634 15648 21640 15700
rect 21692 15688 21698 15700
rect 22465 15691 22523 15697
rect 22465 15688 22477 15691
rect 21692 15660 22477 15688
rect 21692 15648 21698 15660
rect 22465 15657 22477 15660
rect 22511 15657 22523 15691
rect 22465 15651 22523 15657
rect 22756 15660 23060 15688
rect 22756 15620 22784 15660
rect 21560 15592 22784 15620
rect 22833 15623 22891 15629
rect 22833 15589 22845 15623
rect 22879 15620 22891 15623
rect 22922 15620 22928 15632
rect 22879 15592 22928 15620
rect 22879 15589 22891 15592
rect 22833 15583 22891 15589
rect 22922 15580 22928 15592
rect 22980 15580 22986 15632
rect 23032 15620 23060 15660
rect 23658 15648 23664 15700
rect 23716 15688 23722 15700
rect 24489 15691 24547 15697
rect 24489 15688 24501 15691
rect 23716 15660 24501 15688
rect 23716 15648 23722 15660
rect 24489 15657 24501 15660
rect 24535 15688 24547 15691
rect 24578 15688 24584 15700
rect 24535 15660 24584 15688
rect 24535 15657 24547 15660
rect 24489 15651 24547 15657
rect 24578 15648 24584 15660
rect 24636 15648 24642 15700
rect 29730 15620 29736 15632
rect 23032 15592 29736 15620
rect 29730 15580 29736 15592
rect 29788 15580 29794 15632
rect 16573 15524 18368 15552
rect 16485 15515 16543 15521
rect 15068 15388 15148 15416
rect 15212 15456 16344 15484
rect 15068 15376 15074 15388
rect 15212 15348 15240 15456
rect 16209 15419 16267 15425
rect 16209 15416 16221 15419
rect 15488 15388 16221 15416
rect 15488 15360 15516 15388
rect 16209 15385 16221 15388
rect 16255 15385 16267 15419
rect 16500 15416 16528 15515
rect 19426 15512 19432 15564
rect 19484 15552 19490 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 19484 15524 20269 15552
rect 19484 15512 19490 15524
rect 20257 15521 20269 15524
rect 20303 15552 20315 15555
rect 20622 15552 20628 15564
rect 20303 15524 20628 15552
rect 20303 15521 20315 15524
rect 20257 15515 20315 15521
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 20990 15512 20996 15564
rect 21048 15552 21054 15564
rect 21048 15524 22692 15552
rect 21048 15512 21054 15524
rect 17034 15444 17040 15496
rect 17092 15444 17098 15496
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15484 19671 15487
rect 20162 15484 20168 15496
rect 19659 15456 20168 15484
rect 19659 15453 19671 15456
rect 19613 15447 19671 15453
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 21652 15470 21680 15524
rect 22554 15484 22560 15496
rect 21836 15456 22560 15484
rect 17310 15416 17316 15428
rect 16500 15388 17316 15416
rect 16209 15379 16267 15385
rect 17310 15376 17316 15388
rect 17368 15376 17374 15428
rect 17770 15376 17776 15428
rect 17828 15376 17834 15428
rect 19150 15376 19156 15428
rect 19208 15416 19214 15428
rect 20533 15419 20591 15425
rect 20533 15416 20545 15419
rect 19208 15388 20545 15416
rect 19208 15376 19214 15388
rect 20533 15385 20545 15388
rect 20579 15385 20591 15419
rect 20533 15379 20591 15385
rect 14936 15320 15240 15348
rect 14461 15311 14519 15317
rect 15470 15308 15476 15360
rect 15528 15308 15534 15360
rect 16114 15308 16120 15360
rect 16172 15348 16178 15360
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 16172 15320 16313 15348
rect 16172 15308 16178 15320
rect 16301 15317 16313 15320
rect 16347 15348 16359 15351
rect 16390 15348 16396 15360
rect 16347 15320 16396 15348
rect 16347 15317 16359 15320
rect 16301 15311 16359 15317
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 17402 15308 17408 15360
rect 17460 15348 17466 15360
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 17460 15320 18797 15348
rect 17460 15308 17466 15320
rect 18785 15317 18797 15320
rect 18831 15317 18843 15351
rect 18785 15311 18843 15317
rect 19334 15308 19340 15360
rect 19392 15348 19398 15360
rect 19429 15351 19487 15357
rect 19429 15348 19441 15351
rect 19392 15320 19441 15348
rect 19392 15308 19398 15320
rect 19429 15317 19441 15320
rect 19475 15317 19487 15351
rect 20548 15348 20576 15379
rect 21836 15348 21864 15456
rect 22554 15444 22560 15456
rect 22612 15444 22618 15496
rect 20548 15320 21864 15348
rect 19429 15311 19487 15317
rect 21910 15308 21916 15360
rect 21968 15348 21974 15360
rect 22005 15351 22063 15357
rect 22005 15348 22017 15351
rect 21968 15320 22017 15348
rect 21968 15308 21974 15320
rect 22005 15317 22017 15320
rect 22051 15317 22063 15351
rect 22005 15311 22063 15317
rect 22373 15351 22431 15357
rect 22373 15317 22385 15351
rect 22419 15348 22431 15351
rect 22664 15348 22692 15524
rect 22940 15484 22968 15580
rect 25774 15512 25780 15564
rect 25832 15512 25838 15564
rect 23109 15487 23167 15493
rect 23109 15484 23121 15487
rect 22940 15456 23121 15484
rect 23109 15453 23121 15456
rect 23155 15484 23167 15487
rect 23290 15484 23296 15496
rect 23155 15456 23296 15484
rect 23155 15453 23167 15456
rect 23109 15447 23167 15453
rect 23290 15444 23296 15456
rect 23348 15444 23354 15496
rect 26142 15444 26148 15496
rect 26200 15484 26206 15496
rect 37274 15484 37280 15496
rect 26200 15456 37280 15484
rect 26200 15444 26206 15456
rect 37274 15444 37280 15456
rect 37332 15444 37338 15496
rect 23934 15376 23940 15428
rect 23992 15376 23998 15428
rect 25685 15419 25743 15425
rect 25685 15385 25697 15419
rect 25731 15416 25743 15419
rect 25731 15388 26556 15416
rect 25731 15385 25743 15388
rect 25685 15379 25743 15385
rect 23382 15348 23388 15360
rect 22419 15320 23388 15348
rect 22419 15317 22431 15320
rect 22373 15311 22431 15317
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 25222 15308 25228 15360
rect 25280 15308 25286 15360
rect 25590 15308 25596 15360
rect 25648 15348 25654 15360
rect 26142 15348 26148 15360
rect 25648 15320 26148 15348
rect 25648 15308 25654 15320
rect 26142 15308 26148 15320
rect 26200 15348 26206 15360
rect 26528 15357 26556 15388
rect 26237 15351 26295 15357
rect 26237 15348 26249 15351
rect 26200 15320 26249 15348
rect 26200 15308 26206 15320
rect 26237 15317 26249 15320
rect 26283 15317 26295 15351
rect 26237 15311 26295 15317
rect 26513 15351 26571 15357
rect 26513 15317 26525 15351
rect 26559 15348 26571 15351
rect 26878 15348 26884 15360
rect 26559 15320 26884 15348
rect 26559 15317 26571 15320
rect 26513 15311 26571 15317
rect 26878 15308 26884 15320
rect 26936 15348 26942 15360
rect 44818 15348 44824 15360
rect 26936 15320 44824 15348
rect 26936 15308 26942 15320
rect 44818 15308 44824 15320
rect 44876 15308 44882 15360
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 3510 15104 3516 15156
rect 3568 15104 3574 15156
rect 3786 15104 3792 15156
rect 3844 15144 3850 15156
rect 4614 15144 4620 15156
rect 3844 15116 4620 15144
rect 3844 15104 3850 15116
rect 4614 15104 4620 15116
rect 4672 15104 4678 15156
rect 4706 15104 4712 15156
rect 4764 15144 4770 15156
rect 6733 15147 6791 15153
rect 6733 15144 6745 15147
rect 4764 15116 6745 15144
rect 4764 15104 4770 15116
rect 6733 15113 6745 15116
rect 6779 15113 6791 15147
rect 6733 15107 6791 15113
rect 7653 15147 7711 15153
rect 7653 15113 7665 15147
rect 7699 15144 7711 15147
rect 7926 15144 7932 15156
rect 7699 15116 7932 15144
rect 7699 15113 7711 15116
rect 7653 15107 7711 15113
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 9585 15147 9643 15153
rect 9585 15113 9597 15147
rect 9631 15144 9643 15147
rect 11238 15144 11244 15156
rect 9631 15116 11244 15144
rect 9631 15113 9643 15116
rect 9585 15107 9643 15113
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 15470 15144 15476 15156
rect 12406 15116 15476 15144
rect 4430 15076 4436 15088
rect 1780 15048 4436 15076
rect 1780 15017 1808 15048
rect 4430 15036 4436 15048
rect 4488 15036 4494 15088
rect 5810 15036 5816 15088
rect 5868 15076 5874 15088
rect 7745 15079 7803 15085
rect 7745 15076 7757 15079
rect 5868 15048 7757 15076
rect 5868 15036 5874 15048
rect 7745 15045 7757 15048
rect 7791 15045 7803 15079
rect 7745 15039 7803 15045
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 14977 1823 15011
rect 1765 14971 1823 14977
rect 2866 14968 2872 15020
rect 2924 15008 2930 15020
rect 3510 15008 3516 15020
rect 2924 14980 3516 15008
rect 2924 14968 2930 14980
rect 3510 14968 3516 14980
rect 3568 15008 3574 15020
rect 3697 15011 3755 15017
rect 3697 15008 3709 15011
rect 3568 14980 3709 15008
rect 3568 14968 3574 14980
rect 3697 14977 3709 14980
rect 3743 14977 3755 15011
rect 3697 14971 3755 14977
rect 4154 14968 4160 15020
rect 4212 14968 4218 15020
rect 5534 14968 5540 15020
rect 5592 14968 5598 15020
rect 6454 14968 6460 15020
rect 6512 15008 6518 15020
rect 6641 15011 6699 15017
rect 6641 15008 6653 15011
rect 6512 14980 6653 15008
rect 6512 14968 6518 14980
rect 6641 14977 6653 14980
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 7760 15008 7788 15039
rect 8846 15036 8852 15088
rect 8904 15076 8910 15088
rect 9677 15079 9735 15085
rect 9677 15076 9689 15079
rect 8904 15048 9689 15076
rect 8904 15036 8910 15048
rect 9677 15045 9689 15048
rect 9723 15045 9735 15079
rect 9677 15039 9735 15045
rect 10042 15036 10048 15088
rect 10100 15076 10106 15088
rect 10502 15076 10508 15088
rect 10100 15048 10508 15076
rect 10100 15036 10106 15048
rect 10502 15036 10508 15048
rect 10560 15036 10566 15088
rect 10594 15036 10600 15088
rect 10652 15076 10658 15088
rect 10781 15079 10839 15085
rect 10781 15076 10793 15079
rect 10652 15048 10793 15076
rect 10652 15036 10658 15048
rect 10781 15045 10793 15048
rect 10827 15045 10839 15079
rect 12406 15076 12434 15116
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 22094 15144 22100 15156
rect 18472 15116 22100 15144
rect 18472 15104 18478 15116
rect 22094 15104 22100 15116
rect 22152 15104 22158 15156
rect 22554 15104 22560 15156
rect 22612 15144 22618 15156
rect 23753 15147 23811 15153
rect 23753 15144 23765 15147
rect 22612 15116 23765 15144
rect 22612 15104 22618 15116
rect 23753 15113 23765 15116
rect 23799 15113 23811 15147
rect 23753 15107 23811 15113
rect 24946 15104 24952 15156
rect 25004 15104 25010 15156
rect 27062 15104 27068 15156
rect 27120 15104 27126 15156
rect 14918 15076 14924 15088
rect 10781 15039 10839 15045
rect 10888 15048 12434 15076
rect 12544 15048 14924 15076
rect 8573 15011 8631 15017
rect 6788 14980 7696 15008
rect 7760 14980 8524 15008
rect 6788 14968 6794 14980
rect 1302 14900 1308 14952
rect 1360 14940 1366 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 1360 14912 2053 14940
rect 1360 14900 1366 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 4433 14943 4491 14949
rect 4433 14909 4445 14943
rect 4479 14940 4491 14943
rect 4798 14940 4804 14952
rect 4479 14912 4804 14940
rect 4479 14909 4491 14912
rect 4433 14903 4491 14909
rect 4798 14900 4804 14912
rect 4856 14900 4862 14952
rect 4890 14900 4896 14952
rect 4948 14940 4954 14952
rect 4948 14912 5580 14940
rect 4948 14900 4954 14912
rect 5552 14872 5580 14912
rect 5902 14900 5908 14952
rect 5960 14940 5966 14952
rect 7668 14940 7696 14980
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 5960 14912 7512 14940
rect 7668 14912 7849 14940
rect 5960 14900 5966 14912
rect 7484 14872 7512 14912
rect 7837 14909 7849 14912
rect 7883 14909 7895 14943
rect 8496 14940 8524 14980
rect 8573 14977 8585 15011
rect 8619 15008 8631 15011
rect 8662 15008 8668 15020
rect 8619 14980 8668 15008
rect 8619 14977 8631 14980
rect 8573 14971 8631 14977
rect 8662 14968 8668 14980
rect 8720 14968 8726 15020
rect 9306 14968 9312 15020
rect 9364 15008 9370 15020
rect 10888 15017 10916 15048
rect 10873 15011 10931 15017
rect 10873 15008 10885 15011
rect 9364 14980 10885 15008
rect 9364 14968 9370 14980
rect 10873 14977 10885 14980
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 11698 14968 11704 15020
rect 11756 14968 11762 15020
rect 11974 14968 11980 15020
rect 12032 14968 12038 15020
rect 9582 14940 9588 14952
rect 8496 14912 9588 14940
rect 7837 14903 7895 14909
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 9674 14900 9680 14952
rect 9732 14940 9738 14952
rect 9861 14943 9919 14949
rect 9861 14940 9873 14943
rect 9732 14912 9873 14940
rect 9732 14900 9738 14912
rect 9861 14909 9873 14912
rect 9907 14940 9919 14943
rect 10778 14940 10784 14952
rect 9907 14912 10784 14940
rect 9907 14909 9919 14912
rect 9861 14903 9919 14909
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 10965 14943 11023 14949
rect 10965 14940 10977 14943
rect 10888 14912 10977 14940
rect 7926 14872 7932 14884
rect 5552 14844 7420 14872
rect 7484 14844 7932 14872
rect 4430 14764 4436 14816
rect 4488 14804 4494 14816
rect 5905 14807 5963 14813
rect 5905 14804 5917 14807
rect 4488 14776 5917 14804
rect 4488 14764 4494 14776
rect 5905 14773 5917 14776
rect 5951 14804 5963 14807
rect 6914 14804 6920 14816
rect 5951 14776 6920 14804
rect 5951 14773 5963 14776
rect 5905 14767 5963 14773
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 7282 14764 7288 14816
rect 7340 14764 7346 14816
rect 7392 14804 7420 14844
rect 7926 14832 7932 14844
rect 7984 14872 7990 14884
rect 10318 14872 10324 14884
rect 7984 14844 10324 14872
rect 7984 14832 7990 14844
rect 10318 14832 10324 14844
rect 10376 14832 10382 14884
rect 10413 14875 10471 14881
rect 10413 14841 10425 14875
rect 10459 14872 10471 14875
rect 10594 14872 10600 14884
rect 10459 14844 10600 14872
rect 10459 14841 10471 14844
rect 10413 14835 10471 14841
rect 10594 14832 10600 14844
rect 10652 14832 10658 14884
rect 8202 14804 8208 14816
rect 7392 14776 8208 14804
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 8478 14764 8484 14816
rect 8536 14804 8542 14816
rect 8665 14807 8723 14813
rect 8665 14804 8677 14807
rect 8536 14776 8677 14804
rect 8536 14764 8542 14776
rect 8665 14773 8677 14776
rect 8711 14773 8723 14807
rect 8665 14767 8723 14773
rect 8846 14764 8852 14816
rect 8904 14804 8910 14816
rect 9217 14807 9275 14813
rect 9217 14804 9229 14807
rect 8904 14776 9229 14804
rect 8904 14764 8910 14776
rect 9217 14773 9229 14776
rect 9263 14773 9275 14807
rect 9217 14767 9275 14773
rect 9398 14764 9404 14816
rect 9456 14804 9462 14816
rect 10888 14804 10916 14912
rect 10965 14909 10977 14912
rect 11011 14909 11023 14943
rect 10965 14903 11023 14909
rect 11790 14900 11796 14952
rect 11848 14940 11854 14952
rect 12544 14940 12572 15048
rect 14918 15036 14924 15048
rect 14976 15036 14982 15088
rect 15378 15036 15384 15088
rect 15436 15036 15442 15088
rect 16390 15036 16396 15088
rect 16448 15076 16454 15088
rect 16761 15079 16819 15085
rect 16761 15076 16773 15079
rect 16448 15048 16773 15076
rect 16448 15036 16454 15048
rect 16761 15045 16773 15048
rect 16807 15076 16819 15079
rect 16807 15048 20208 15076
rect 16807 15045 16819 15048
rect 16761 15039 16819 15045
rect 13354 14968 13360 15020
rect 13412 14968 13418 15020
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 15008 13507 15011
rect 14001 15011 14059 15017
rect 14001 15008 14013 15011
rect 13495 14980 14013 15008
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 14001 14977 14013 14980
rect 14047 15008 14059 15011
rect 14047 14980 14228 15008
rect 14047 14977 14059 14980
rect 14001 14971 14059 14977
rect 11848 14912 12572 14940
rect 11848 14900 11854 14912
rect 13262 14900 13268 14952
rect 13320 14940 13326 14952
rect 13541 14943 13599 14949
rect 13541 14940 13553 14943
rect 13320 14912 13553 14940
rect 13320 14900 13326 14912
rect 13541 14909 13553 14912
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 12618 14832 12624 14884
rect 12676 14872 12682 14884
rect 12989 14875 13047 14881
rect 12989 14872 13001 14875
rect 12676 14844 13001 14872
rect 12676 14832 12682 14844
rect 12989 14841 13001 14844
rect 13035 14841 13047 14875
rect 13556 14872 13584 14903
rect 13722 14872 13728 14884
rect 13556 14844 13728 14872
rect 12989 14835 13047 14841
rect 13722 14832 13728 14844
rect 13780 14832 13786 14884
rect 14200 14872 14228 14980
rect 17126 14968 17132 15020
rect 17184 14968 17190 15020
rect 17770 14968 17776 15020
rect 17828 15008 17834 15020
rect 19153 15011 19211 15017
rect 19153 15008 19165 15011
rect 17828 14980 19165 15008
rect 17828 14968 17834 14980
rect 19153 14977 19165 14980
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 19484 14980 20085 15008
rect 19484 14968 19490 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20180 15008 20208 15048
rect 20254 15036 20260 15088
rect 20312 15076 20318 15088
rect 20714 15076 20720 15088
rect 20312 15048 20720 15076
rect 20312 15036 20318 15048
rect 20714 15036 20720 15048
rect 20772 15036 20778 15088
rect 20901 15079 20959 15085
rect 20901 15045 20913 15079
rect 20947 15076 20959 15079
rect 20990 15076 20996 15088
rect 20947 15048 20996 15076
rect 20947 15045 20959 15048
rect 20901 15039 20959 15045
rect 20990 15036 20996 15048
rect 21048 15036 21054 15088
rect 22186 15036 22192 15088
rect 22244 15076 22250 15088
rect 22281 15079 22339 15085
rect 22281 15076 22293 15079
rect 22244 15048 22293 15076
rect 22244 15036 22250 15048
rect 22281 15045 22293 15048
rect 22327 15045 22339 15079
rect 24964 15076 24992 15104
rect 25133 15079 25191 15085
rect 25133 15076 25145 15079
rect 24964 15048 25145 15076
rect 22281 15039 22339 15045
rect 25133 15045 25145 15048
rect 25179 15045 25191 15079
rect 27080 15076 27108 15104
rect 26358 15048 27108 15076
rect 25133 15039 25191 15045
rect 20180 14980 20484 15008
rect 20073 14971 20131 14977
rect 14274 14900 14280 14952
rect 14332 14940 14338 14952
rect 14553 14943 14611 14949
rect 14553 14940 14565 14943
rect 14332 14912 14565 14940
rect 14332 14900 14338 14912
rect 14553 14909 14565 14912
rect 14599 14909 14611 14943
rect 14553 14903 14611 14909
rect 14829 14943 14887 14949
rect 14829 14909 14841 14943
rect 14875 14940 14887 14943
rect 14918 14940 14924 14952
rect 14875 14912 14924 14940
rect 14875 14909 14887 14912
rect 14829 14903 14887 14909
rect 14918 14900 14924 14912
rect 14976 14900 14982 14952
rect 15562 14900 15568 14952
rect 15620 14940 15626 14952
rect 19610 14940 19616 14952
rect 15620 14912 19616 14940
rect 15620 14900 15626 14912
rect 19610 14900 19616 14912
rect 19668 14900 19674 14952
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14940 20223 14943
rect 20254 14940 20260 14952
rect 20211 14912 20260 14940
rect 20211 14909 20223 14912
rect 20165 14903 20223 14909
rect 20254 14900 20260 14912
rect 20312 14900 20318 14952
rect 20349 14943 20407 14949
rect 20349 14909 20361 14943
rect 20395 14909 20407 14943
rect 20456 14940 20484 14980
rect 20622 14968 20628 15020
rect 20680 15008 20686 15020
rect 22002 15008 22008 15020
rect 20680 14980 22008 15008
rect 20680 14968 20686 14980
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 23382 14968 23388 15020
rect 23440 14968 23446 15020
rect 23934 14968 23940 15020
rect 23992 15008 23998 15020
rect 24857 15011 24915 15017
rect 24857 15008 24869 15011
rect 23992 14980 24869 15008
rect 23992 14968 23998 14980
rect 24857 14977 24869 14980
rect 24903 14977 24915 15011
rect 24857 14971 24915 14977
rect 20456 14912 24992 14940
rect 20349 14903 20407 14909
rect 16942 14872 16948 14884
rect 14200 14844 14688 14872
rect 9456 14776 10916 14804
rect 9456 14764 9462 14776
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 13814 14804 13820 14816
rect 11204 14776 13820 14804
rect 11204 14764 11210 14776
rect 13814 14764 13820 14776
rect 13872 14804 13878 14816
rect 14185 14807 14243 14813
rect 14185 14804 14197 14807
rect 13872 14776 14197 14804
rect 13872 14764 13878 14776
rect 14185 14773 14197 14776
rect 14231 14773 14243 14807
rect 14660 14804 14688 14844
rect 16224 14844 16948 14872
rect 16224 14804 16252 14844
rect 16942 14832 16948 14844
rect 17000 14832 17006 14884
rect 17494 14832 17500 14884
rect 17552 14872 17558 14884
rect 19705 14875 19763 14881
rect 17552 14844 19472 14872
rect 17552 14832 17558 14844
rect 14660 14776 16252 14804
rect 14185 14767 14243 14773
rect 16298 14764 16304 14816
rect 16356 14764 16362 14816
rect 16960 14804 16988 14832
rect 19242 14804 19248 14816
rect 16960 14776 19248 14804
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 19334 14764 19340 14816
rect 19392 14764 19398 14816
rect 19444 14804 19472 14844
rect 19705 14841 19717 14875
rect 19751 14872 19763 14875
rect 19978 14872 19984 14884
rect 19751 14844 19984 14872
rect 19751 14841 19763 14844
rect 19705 14835 19763 14841
rect 19978 14832 19984 14844
rect 20036 14832 20042 14884
rect 20364 14872 20392 14903
rect 21910 14872 21916 14884
rect 20364 14844 21916 14872
rect 21910 14832 21916 14844
rect 21968 14832 21974 14884
rect 23382 14832 23388 14884
rect 23440 14872 23446 14884
rect 23440 14844 23888 14872
rect 23440 14832 23446 14844
rect 23860 14816 23888 14844
rect 20717 14807 20775 14813
rect 20717 14804 20729 14807
rect 19444 14776 20729 14804
rect 20717 14773 20729 14776
rect 20763 14804 20775 14807
rect 20990 14804 20996 14816
rect 20763 14776 20996 14804
rect 20763 14773 20775 14776
rect 20717 14767 20775 14773
rect 20990 14764 20996 14776
rect 21048 14764 21054 14816
rect 23842 14764 23848 14816
rect 23900 14804 23906 14816
rect 24029 14807 24087 14813
rect 24029 14804 24041 14807
rect 23900 14776 24041 14804
rect 23900 14764 23906 14776
rect 24029 14773 24041 14776
rect 24075 14804 24087 14807
rect 24213 14807 24271 14813
rect 24213 14804 24225 14807
rect 24075 14776 24225 14804
rect 24075 14773 24087 14776
rect 24029 14767 24087 14773
rect 24213 14773 24225 14776
rect 24259 14773 24271 14807
rect 24964 14804 24992 14912
rect 25314 14804 25320 14816
rect 24964 14776 25320 14804
rect 24213 14767 24271 14773
rect 25314 14764 25320 14776
rect 25372 14764 25378 14816
rect 26602 14764 26608 14816
rect 26660 14764 26666 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 3973 14603 4031 14609
rect 3973 14569 3985 14603
rect 4019 14600 4031 14603
rect 4019 14572 5580 14600
rect 4019 14569 4031 14572
rect 3973 14563 4031 14569
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 5350 14532 5356 14544
rect 4212 14504 5356 14532
rect 4212 14492 4218 14504
rect 5350 14492 5356 14504
rect 5408 14492 5414 14544
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1360 14436 2053 14464
rect 1360 14424 1366 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 4430 14424 4436 14476
rect 4488 14464 4494 14476
rect 4801 14467 4859 14473
rect 4801 14464 4813 14467
rect 4488 14436 4813 14464
rect 4488 14424 4494 14436
rect 4801 14433 4813 14436
rect 4847 14433 4859 14467
rect 5552 14464 5580 14572
rect 5718 14560 5724 14612
rect 5776 14600 5782 14612
rect 9401 14603 9459 14609
rect 5776 14572 8524 14600
rect 5776 14560 5782 14572
rect 6822 14492 6828 14544
rect 6880 14532 6886 14544
rect 8202 14532 8208 14544
rect 6880 14504 8208 14532
rect 6880 14492 6886 14504
rect 8202 14492 8208 14504
rect 8260 14492 8266 14544
rect 8496 14532 8524 14572
rect 9401 14569 9413 14603
rect 9447 14600 9459 14603
rect 9490 14600 9496 14612
rect 9447 14572 9496 14600
rect 9447 14569 9459 14572
rect 9401 14563 9459 14569
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 9640 14572 11621 14600
rect 9640 14560 9646 14572
rect 11609 14569 11621 14572
rect 11655 14600 11667 14603
rect 13354 14600 13360 14612
rect 11655 14572 13360 14600
rect 11655 14569 11667 14572
rect 11609 14563 11667 14569
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 13722 14560 13728 14612
rect 13780 14560 13786 14612
rect 14369 14603 14427 14609
rect 14369 14569 14381 14603
rect 14415 14600 14427 14603
rect 14734 14600 14740 14612
rect 14415 14572 14740 14600
rect 14415 14569 14427 14572
rect 14369 14563 14427 14569
rect 14734 14560 14740 14572
rect 14792 14560 14798 14612
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 18601 14603 18659 14609
rect 18601 14600 18613 14603
rect 14976 14572 18613 14600
rect 14976 14560 14982 14572
rect 18601 14569 18613 14572
rect 18647 14569 18659 14603
rect 18601 14563 18659 14569
rect 19429 14603 19487 14609
rect 19429 14569 19441 14603
rect 19475 14600 19487 14603
rect 35066 14600 35072 14612
rect 19475 14572 35072 14600
rect 19475 14569 19487 14572
rect 19429 14563 19487 14569
rect 35066 14560 35072 14572
rect 35124 14560 35130 14612
rect 11790 14532 11796 14544
rect 8496 14504 11796 14532
rect 11790 14492 11796 14504
rect 11848 14492 11854 14544
rect 13814 14492 13820 14544
rect 13872 14532 13878 14544
rect 14182 14532 14188 14544
rect 13872 14504 14188 14532
rect 13872 14492 13878 14504
rect 14182 14492 14188 14504
rect 14240 14492 14246 14544
rect 14274 14492 14280 14544
rect 14332 14532 14338 14544
rect 14332 14504 14688 14532
rect 14332 14492 14338 14504
rect 6454 14464 6460 14476
rect 5552 14436 6460 14464
rect 4801 14427 4859 14433
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 6730 14424 6736 14476
rect 6788 14464 6794 14476
rect 6914 14464 6920 14476
rect 6788 14436 6920 14464
rect 6788 14424 6794 14436
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 7006 14424 7012 14476
rect 7064 14464 7070 14476
rect 7193 14467 7251 14473
rect 7193 14464 7205 14467
rect 7064 14436 7205 14464
rect 7064 14424 7070 14436
rect 7193 14433 7205 14436
rect 7239 14433 7251 14467
rect 7193 14427 7251 14433
rect 7742 14424 7748 14476
rect 7800 14464 7806 14476
rect 8297 14467 8355 14473
rect 8297 14464 8309 14467
rect 7800 14436 8309 14464
rect 7800 14424 7806 14436
rect 8297 14433 8309 14436
rect 8343 14433 8355 14467
rect 8297 14427 8355 14433
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14464 8539 14467
rect 9674 14464 9680 14476
rect 8527 14436 9680 14464
rect 8527 14433 8539 14436
rect 8481 14427 8539 14433
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 10042 14424 10048 14476
rect 10100 14424 10106 14476
rect 10410 14424 10416 14476
rect 10468 14464 10474 14476
rect 10594 14464 10600 14476
rect 10468 14436 10600 14464
rect 10468 14424 10474 14436
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 10962 14464 10968 14476
rect 10744 14436 10968 14464
rect 10744 14424 10750 14436
rect 10962 14424 10968 14436
rect 11020 14464 11026 14476
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 11020 14436 11161 14464
rect 11020 14424 11026 14436
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 11149 14427 11207 14433
rect 12253 14467 12311 14473
rect 12253 14433 12265 14467
rect 12299 14464 12311 14467
rect 13446 14464 13452 14476
rect 12299 14436 13452 14464
rect 12299 14433 12311 14436
rect 12253 14427 12311 14433
rect 13446 14424 13452 14436
rect 13504 14464 13510 14476
rect 13722 14464 13728 14476
rect 13504 14436 13728 14464
rect 13504 14424 13510 14436
rect 13722 14424 13728 14436
rect 13780 14424 13786 14476
rect 14660 14473 14688 14504
rect 21542 14492 21548 14544
rect 21600 14532 21606 14544
rect 21729 14535 21787 14541
rect 21729 14532 21741 14535
rect 21600 14504 21741 14532
rect 21600 14492 21606 14504
rect 21729 14501 21741 14504
rect 21775 14501 21787 14535
rect 21729 14495 21787 14501
rect 23566 14492 23572 14544
rect 23624 14532 23630 14544
rect 24029 14535 24087 14541
rect 24029 14532 24041 14535
rect 23624 14504 24041 14532
rect 23624 14492 23630 14504
rect 24029 14501 24041 14504
rect 24075 14532 24087 14535
rect 25774 14532 25780 14544
rect 24075 14504 25780 14532
rect 24075 14501 24087 14504
rect 24029 14495 24087 14501
rect 25774 14492 25780 14504
rect 25832 14492 25838 14544
rect 26878 14532 26884 14544
rect 26252 14504 26884 14532
rect 14645 14467 14703 14473
rect 14645 14433 14657 14467
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 16298 14464 16304 14476
rect 14967 14436 16304 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 16853 14467 16911 14473
rect 16853 14433 16865 14467
rect 16899 14464 16911 14467
rect 17126 14464 17132 14476
rect 16899 14436 17132 14464
rect 16899 14433 16911 14436
rect 16853 14427 16911 14433
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 17218 14424 17224 14476
rect 17276 14464 17282 14476
rect 20070 14464 20076 14476
rect 17276 14436 20076 14464
rect 17276 14424 17282 14436
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 20162 14424 20168 14476
rect 20220 14464 20226 14476
rect 21085 14467 21143 14473
rect 21085 14464 21097 14467
rect 20220 14436 21097 14464
rect 20220 14424 20226 14436
rect 21085 14433 21097 14436
rect 21131 14433 21143 14467
rect 21085 14427 21143 14433
rect 22002 14424 22008 14476
rect 22060 14464 22066 14476
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 22060 14436 22293 14464
rect 22060 14424 22066 14436
rect 22281 14433 22293 14436
rect 22327 14464 22339 14467
rect 23934 14464 23940 14476
rect 22327 14436 23940 14464
rect 22327 14433 22339 14436
rect 22281 14427 22339 14433
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 25133 14467 25191 14473
rect 25133 14433 25145 14467
rect 25179 14433 25191 14467
rect 25133 14427 25191 14433
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 1811 14368 5120 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 2590 14288 2596 14340
rect 2648 14328 2654 14340
rect 4617 14331 4675 14337
rect 4617 14328 4629 14331
rect 2648 14300 4629 14328
rect 2648 14288 2654 14300
rect 4617 14297 4629 14300
rect 4663 14297 4675 14331
rect 4617 14291 4675 14297
rect 2866 14220 2872 14272
rect 2924 14260 2930 14272
rect 3329 14263 3387 14269
rect 3329 14260 3341 14263
rect 2924 14232 3341 14260
rect 2924 14220 2930 14232
rect 3329 14229 3341 14232
rect 3375 14260 3387 14263
rect 3513 14263 3571 14269
rect 3513 14260 3525 14263
rect 3375 14232 3525 14260
rect 3375 14229 3387 14232
rect 3329 14223 3387 14229
rect 3513 14229 3525 14232
rect 3559 14229 3571 14263
rect 3513 14223 3571 14229
rect 4249 14263 4307 14269
rect 4249 14229 4261 14263
rect 4295 14260 4307 14263
rect 4522 14260 4528 14272
rect 4295 14232 4528 14260
rect 4295 14229 4307 14232
rect 4249 14223 4307 14229
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 4706 14220 4712 14272
rect 4764 14220 4770 14272
rect 5092 14260 5120 14368
rect 5166 14356 5172 14408
rect 5224 14396 5230 14408
rect 5445 14399 5503 14405
rect 5445 14396 5457 14399
rect 5224 14368 5457 14396
rect 5224 14356 5230 14368
rect 5445 14365 5457 14368
rect 5491 14365 5503 14399
rect 5445 14359 5503 14365
rect 6822 14356 6828 14408
rect 6880 14356 6886 14408
rect 6932 14396 6960 14424
rect 9398 14396 9404 14408
rect 6932 14368 9404 14396
rect 9398 14356 9404 14368
rect 9456 14356 9462 14408
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14396 9919 14399
rect 10870 14396 10876 14408
rect 9907 14368 10876 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 11974 14356 11980 14408
rect 12032 14356 12038 14408
rect 18138 14356 18144 14408
rect 18196 14396 18202 14408
rect 18877 14399 18935 14405
rect 18877 14396 18889 14399
rect 18196 14368 18889 14396
rect 18196 14356 18202 14368
rect 18877 14365 18889 14368
rect 18923 14365 18935 14399
rect 18877 14359 18935 14365
rect 19610 14356 19616 14408
rect 19668 14356 19674 14408
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20772 14368 20913 14396
rect 20772 14356 20778 14368
rect 20901 14365 20913 14368
rect 20947 14396 20959 14399
rect 21545 14399 21603 14405
rect 21545 14396 21557 14399
rect 20947 14368 21557 14396
rect 20947 14365 20959 14368
rect 20901 14359 20959 14365
rect 21545 14365 21557 14368
rect 21591 14396 21603 14399
rect 21818 14396 21824 14408
rect 21591 14368 21824 14396
rect 21591 14365 21603 14368
rect 21545 14359 21603 14365
rect 21818 14356 21824 14368
rect 21876 14356 21882 14408
rect 25148 14396 25176 14427
rect 25590 14424 25596 14476
rect 25648 14464 25654 14476
rect 26252 14473 26280 14504
rect 26878 14492 26884 14504
rect 26936 14492 26942 14544
rect 26237 14467 26295 14473
rect 26237 14464 26249 14467
rect 25648 14436 26249 14464
rect 25648 14424 25654 14436
rect 26237 14433 26249 14436
rect 26283 14433 26295 14467
rect 26237 14427 26295 14433
rect 26329 14467 26387 14473
rect 26329 14433 26341 14467
rect 26375 14464 26387 14467
rect 26602 14464 26608 14476
rect 26375 14436 26608 14464
rect 26375 14433 26387 14436
rect 26329 14427 26387 14433
rect 26344 14396 26372 14427
rect 26602 14424 26608 14436
rect 26660 14424 26666 14476
rect 23952 14368 26372 14396
rect 5721 14331 5779 14337
rect 5721 14297 5733 14331
rect 5767 14328 5779 14331
rect 5994 14328 6000 14340
rect 5767 14300 6000 14328
rect 5767 14297 5779 14300
rect 5721 14291 5779 14297
rect 5994 14288 6000 14300
rect 6052 14288 6058 14340
rect 8478 14288 8484 14340
rect 8536 14328 8542 14340
rect 10965 14331 11023 14337
rect 8536 14300 10732 14328
rect 8536 14288 8542 14300
rect 6730 14260 6736 14272
rect 5092 14232 6736 14260
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 7834 14220 7840 14272
rect 7892 14220 7898 14272
rect 8202 14220 8208 14272
rect 8260 14220 8266 14272
rect 8662 14220 8668 14272
rect 8720 14260 8726 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8720 14232 9045 14260
rect 8720 14220 8726 14232
rect 9033 14229 9045 14232
rect 9079 14260 9091 14263
rect 9306 14260 9312 14272
rect 9079 14232 9312 14260
rect 9079 14229 9091 14232
rect 9033 14223 9091 14229
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 9674 14220 9680 14272
rect 9732 14260 9738 14272
rect 9769 14263 9827 14269
rect 9769 14260 9781 14263
rect 9732 14232 9781 14260
rect 9732 14220 9738 14232
rect 9769 14229 9781 14232
rect 9815 14229 9827 14263
rect 9769 14223 9827 14229
rect 10594 14220 10600 14272
rect 10652 14220 10658 14272
rect 10704 14260 10732 14300
rect 10965 14297 10977 14331
rect 11011 14328 11023 14331
rect 11514 14328 11520 14340
rect 11011 14300 11520 14328
rect 11011 14297 11023 14300
rect 10965 14291 11023 14297
rect 11514 14288 11520 14300
rect 11572 14328 11578 14340
rect 13998 14328 14004 14340
rect 11572 14300 12434 14328
rect 13478 14300 14004 14328
rect 11572 14288 11578 14300
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 10704 14232 11069 14260
rect 11057 14229 11069 14232
rect 11103 14260 11115 14263
rect 11146 14260 11152 14272
rect 11103 14232 11152 14260
rect 11103 14229 11115 14232
rect 11057 14223 11115 14229
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 12406 14260 12434 14300
rect 13998 14288 14004 14300
rect 14056 14328 14062 14340
rect 14093 14331 14151 14337
rect 14093 14328 14105 14331
rect 14056 14300 14105 14328
rect 14056 14288 14062 14300
rect 14093 14297 14105 14300
rect 14139 14328 14151 14331
rect 15378 14328 15384 14340
rect 14139 14300 15384 14328
rect 14139 14297 14151 14300
rect 14093 14291 14151 14297
rect 15378 14288 15384 14300
rect 15436 14288 15442 14340
rect 16850 14328 16856 14340
rect 16224 14300 16856 14328
rect 12618 14260 12624 14272
rect 12406 14232 12624 14260
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 12894 14220 12900 14272
rect 12952 14260 12958 14272
rect 16224 14260 16252 14300
rect 16850 14288 16856 14300
rect 16908 14288 16914 14340
rect 17129 14331 17187 14337
rect 17129 14297 17141 14331
rect 17175 14328 17187 14331
rect 17402 14328 17408 14340
rect 17175 14300 17408 14328
rect 17175 14297 17187 14300
rect 17129 14291 17187 14297
rect 17402 14288 17408 14300
rect 17460 14288 17466 14340
rect 17770 14288 17776 14340
rect 17828 14288 17834 14340
rect 21910 14288 21916 14340
rect 21968 14328 21974 14340
rect 22557 14331 22615 14337
rect 22557 14328 22569 14331
rect 21968 14300 22569 14328
rect 21968 14288 21974 14300
rect 22557 14297 22569 14300
rect 22603 14297 22615 14331
rect 23842 14328 23848 14340
rect 23782 14300 23848 14328
rect 22557 14291 22615 14297
rect 23842 14288 23848 14300
rect 23900 14288 23906 14340
rect 12952 14232 16252 14260
rect 12952 14220 12958 14232
rect 16390 14220 16396 14272
rect 16448 14220 16454 14272
rect 16574 14220 16580 14272
rect 16632 14260 16638 14272
rect 18506 14260 18512 14272
rect 16632 14232 18512 14260
rect 16632 14220 16638 14232
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 20530 14220 20536 14272
rect 20588 14220 20594 14272
rect 20993 14263 21051 14269
rect 20993 14229 21005 14263
rect 21039 14260 21051 14263
rect 21542 14260 21548 14272
rect 21039 14232 21548 14260
rect 21039 14229 21051 14232
rect 20993 14223 21051 14229
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 22002 14220 22008 14272
rect 22060 14260 22066 14272
rect 22830 14260 22836 14272
rect 22060 14232 22836 14260
rect 22060 14220 22066 14232
rect 22830 14220 22836 14232
rect 22888 14220 22894 14272
rect 23382 14220 23388 14272
rect 23440 14260 23446 14272
rect 23952 14260 23980 14368
rect 25041 14331 25099 14337
rect 25041 14297 25053 14331
rect 25087 14328 25099 14331
rect 25130 14328 25136 14340
rect 25087 14300 25136 14328
rect 25087 14297 25099 14300
rect 25041 14291 25099 14297
rect 25130 14288 25136 14300
rect 25188 14288 25194 14340
rect 26142 14288 26148 14340
rect 26200 14328 26206 14340
rect 26973 14331 27031 14337
rect 26973 14328 26985 14331
rect 26200 14300 26985 14328
rect 26200 14288 26206 14300
rect 26973 14297 26985 14300
rect 27019 14297 27031 14331
rect 26973 14291 27031 14297
rect 23440 14232 23980 14260
rect 23440 14220 23446 14232
rect 24578 14220 24584 14272
rect 24636 14220 24642 14272
rect 24949 14263 25007 14269
rect 24949 14229 24961 14263
rect 24995 14260 25007 14263
rect 25314 14260 25320 14272
rect 24995 14232 25320 14260
rect 24995 14229 25007 14232
rect 24949 14223 25007 14229
rect 25314 14220 25320 14232
rect 25372 14220 25378 14272
rect 25774 14220 25780 14272
rect 25832 14220 25838 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3418 14016 3424 14068
rect 3476 14016 3482 14068
rect 4065 14059 4123 14065
rect 4065 14025 4077 14059
rect 4111 14056 4123 14059
rect 4706 14056 4712 14068
rect 4111 14028 4712 14056
rect 4111 14025 4123 14028
rect 4065 14019 4123 14025
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 5629 14059 5687 14065
rect 5629 14025 5641 14059
rect 5675 14056 5687 14059
rect 6362 14056 6368 14068
rect 5675 14028 6368 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 6546 14016 6552 14068
rect 6604 14016 6610 14068
rect 6917 14059 6975 14065
rect 6917 14025 6929 14059
rect 6963 14025 6975 14059
rect 6917 14019 6975 14025
rect 2590 13948 2596 14000
rect 2648 13988 2654 14000
rect 4525 13991 4583 13997
rect 4525 13988 4537 13991
rect 2648 13960 4537 13988
rect 2648 13948 2654 13960
rect 4525 13957 4537 13960
rect 4571 13957 4583 13991
rect 4525 13951 4583 13957
rect 4614 13948 4620 14000
rect 4672 13988 4678 14000
rect 5721 13991 5779 13997
rect 5721 13988 5733 13991
rect 4672 13960 5733 13988
rect 4672 13948 4678 13960
rect 5721 13957 5733 13960
rect 5767 13957 5779 13991
rect 5721 13951 5779 13957
rect 6454 13948 6460 14000
rect 6512 13948 6518 14000
rect 6932 13988 6960 14019
rect 7282 14016 7288 14068
rect 7340 14016 7346 14068
rect 7466 14016 7472 14068
rect 7524 14056 7530 14068
rect 7742 14056 7748 14068
rect 7524 14028 7748 14056
rect 7524 14016 7530 14028
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 9214 14056 9220 14068
rect 8159 14028 9220 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9324 14028 10916 14056
rect 8481 13991 8539 13997
rect 8481 13988 8493 13991
rect 6932 13960 8493 13988
rect 8481 13957 8493 13960
rect 8527 13957 8539 13991
rect 8481 13951 8539 13957
rect 8570 13948 8576 14000
rect 8628 13948 8634 14000
rect 1762 13880 1768 13932
rect 1820 13880 1826 13932
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13920 4491 13923
rect 4890 13920 4896 13932
rect 4479 13892 4896 13920
rect 4479 13889 4491 13892
rect 4433 13883 4491 13889
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 3620 13852 3648 13883
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 5258 13880 5264 13932
rect 5316 13920 5322 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 5316 13892 7389 13920
rect 5316 13880 5322 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 9324 13920 9352 14028
rect 10318 13948 10324 14000
rect 10376 13948 10382 14000
rect 10888 13988 10916 14028
rect 11146 14016 11152 14068
rect 11204 14056 11210 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11204 14028 11989 14056
rect 11204 14016 11210 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 12250 14056 12256 14068
rect 11977 14019 12035 14025
rect 12084 14028 12256 14056
rect 11238 13988 11244 14000
rect 10888 13960 11244 13988
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 11606 13948 11612 14000
rect 11664 13948 11670 14000
rect 11790 13948 11796 14000
rect 11848 13988 11854 14000
rect 12084 13988 12112 14028
rect 12250 14016 12256 14028
rect 12308 14056 12314 14068
rect 12345 14059 12403 14065
rect 12345 14056 12357 14059
rect 12308 14028 12357 14056
rect 12308 14016 12314 14028
rect 12345 14025 12357 14028
rect 12391 14025 12403 14059
rect 12345 14019 12403 14025
rect 12618 14016 12624 14068
rect 12676 14056 12682 14068
rect 13078 14056 13084 14068
rect 12676 14028 13084 14056
rect 12676 14016 12682 14028
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 13173 14059 13231 14065
rect 13173 14025 13185 14059
rect 13219 14056 13231 14059
rect 13219 14028 14136 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 11848 13960 12112 13988
rect 11848 13948 11854 13960
rect 12158 13948 12164 14000
rect 12216 13988 12222 14000
rect 12437 13991 12495 13997
rect 12437 13988 12449 13991
rect 12216 13960 12449 13988
rect 12216 13948 12222 13960
rect 12437 13957 12449 13960
rect 12483 13957 12495 13991
rect 13633 13991 13691 13997
rect 13633 13988 13645 13991
rect 12437 13951 12495 13957
rect 12544 13960 13645 13988
rect 7377 13883 7435 13889
rect 7576 13892 9352 13920
rect 3620 13824 4660 13852
rect 2041 13815 2099 13821
rect 4632 13784 4660 13824
rect 4706 13812 4712 13864
rect 4764 13812 4770 13864
rect 5902 13812 5908 13864
rect 5960 13812 5966 13864
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 6788 13824 6960 13852
rect 6788 13812 6794 13824
rect 5718 13784 5724 13796
rect 4632 13756 5724 13784
rect 5718 13744 5724 13756
rect 5776 13744 5782 13796
rect 6086 13744 6092 13796
rect 6144 13784 6150 13796
rect 6362 13784 6368 13796
rect 6144 13756 6368 13784
rect 6144 13744 6150 13756
rect 6362 13744 6368 13756
rect 6420 13744 6426 13796
rect 6932 13784 6960 13824
rect 7006 13812 7012 13864
rect 7064 13852 7070 13864
rect 7469 13855 7527 13861
rect 7469 13852 7481 13855
rect 7064 13824 7481 13852
rect 7064 13812 7070 13824
rect 7469 13821 7481 13824
rect 7515 13821 7527 13855
rect 7469 13815 7527 13821
rect 7576 13784 7604 13892
rect 8478 13812 8484 13864
rect 8536 13852 8542 13864
rect 8665 13855 8723 13861
rect 8665 13852 8677 13855
rect 8536 13824 8677 13852
rect 8536 13812 8542 13824
rect 8665 13821 8677 13824
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 9306 13812 9312 13864
rect 9364 13812 9370 13864
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 11057 13855 11115 13861
rect 11057 13852 11069 13855
rect 10836 13824 11069 13852
rect 10836 13812 10842 13824
rect 11057 13821 11069 13824
rect 11103 13821 11115 13855
rect 11624 13852 11652 13948
rect 12544 13852 12572 13960
rect 13633 13957 13645 13960
rect 13679 13957 13691 13991
rect 14108 13988 14136 14028
rect 14182 14016 14188 14068
rect 14240 14056 14246 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 14240 14028 14749 14056
rect 14240 14016 14246 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 14737 14019 14795 14025
rect 14826 14016 14832 14068
rect 14884 14016 14890 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 16574 14056 16580 14068
rect 15611 14028 16580 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 17310 14016 17316 14068
rect 17368 14056 17374 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 17368 14028 18889 14056
rect 17368 14016 17374 14028
rect 18877 14025 18889 14028
rect 18923 14025 18935 14059
rect 18877 14019 18935 14025
rect 19429 14059 19487 14065
rect 19429 14025 19441 14059
rect 19475 14025 19487 14059
rect 19429 14019 19487 14025
rect 16666 13988 16672 14000
rect 14108 13960 16672 13988
rect 13633 13951 13691 13957
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 17862 13988 17868 14000
rect 17052 13960 17868 13988
rect 13538 13880 13544 13932
rect 13596 13880 13602 13932
rect 15746 13920 15752 13932
rect 13740 13892 15752 13920
rect 11624 13824 12572 13852
rect 12621 13855 12679 13861
rect 11057 13815 11115 13821
rect 12621 13821 12633 13855
rect 12667 13821 12679 13855
rect 12621 13815 12679 13821
rect 12342 13784 12348 13796
rect 6932 13756 7604 13784
rect 10612 13756 12348 13784
rect 5258 13676 5264 13728
rect 5316 13676 5322 13728
rect 5350 13676 5356 13728
rect 5408 13716 5414 13728
rect 9030 13716 9036 13728
rect 5408 13688 9036 13716
rect 5408 13676 5414 13688
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 9572 13719 9630 13725
rect 9572 13685 9584 13719
rect 9618 13716 9630 13719
rect 10612 13716 10640 13756
rect 12342 13744 12348 13756
rect 12400 13784 12406 13796
rect 12636 13784 12664 13815
rect 13078 13812 13084 13864
rect 13136 13852 13142 13864
rect 13740 13852 13768 13892
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 15930 13880 15936 13932
rect 15988 13880 15994 13932
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 16942 13920 16948 13932
rect 16071 13892 16948 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 13136 13824 13768 13852
rect 13136 13812 13142 13824
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 14458 13852 14464 13864
rect 14384 13824 14464 13852
rect 14384 13793 14412 13824
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 14918 13812 14924 13864
rect 14976 13812 14982 13864
rect 16206 13812 16212 13864
rect 16264 13812 16270 13864
rect 17052 13852 17080 13960
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 19444 13988 19472 14019
rect 20070 14016 20076 14068
rect 20128 14016 20134 14068
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 20990 14056 20996 14068
rect 20404 14028 20996 14056
rect 20404 14016 20410 14028
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 21174 14016 21180 14068
rect 21232 14056 21238 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 21232 14028 23397 14056
rect 21232 14016 21238 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 24949 14059 25007 14065
rect 24949 14025 24961 14059
rect 24995 14056 25007 14059
rect 25774 14056 25780 14068
rect 24995 14028 25780 14056
rect 24995 14025 25007 14028
rect 24949 14019 25007 14025
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 20898 13988 20904 14000
rect 19444 13960 20904 13988
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 21818 13948 21824 14000
rect 21876 13988 21882 14000
rect 22649 13991 22707 13997
rect 22649 13988 22661 13991
rect 21876 13960 22661 13988
rect 21876 13948 21882 13960
rect 22649 13957 22661 13960
rect 22695 13988 22707 13991
rect 22695 13960 23888 13988
rect 22695 13957 22707 13960
rect 22649 13951 22707 13957
rect 19613 13923 19671 13929
rect 19613 13920 19625 13923
rect 18616 13892 19625 13920
rect 16684 13824 17080 13852
rect 14369 13787 14427 13793
rect 12400 13756 12664 13784
rect 13096 13756 13400 13784
rect 12400 13744 12406 13756
rect 9618 13688 10640 13716
rect 9618 13685 9630 13688
rect 9572 13679 9630 13685
rect 10686 13676 10692 13728
rect 10744 13716 10750 13728
rect 13096 13716 13124 13756
rect 10744 13688 13124 13716
rect 13372 13716 13400 13756
rect 14369 13753 14381 13787
rect 14415 13753 14427 13787
rect 14369 13747 14427 13753
rect 14826 13744 14832 13796
rect 14884 13784 14890 13796
rect 15194 13784 15200 13796
rect 14884 13756 15200 13784
rect 14884 13744 14890 13756
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 16684 13728 16712 13824
rect 17126 13812 17132 13864
rect 17184 13812 17190 13864
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 18616 13852 18644 13892
rect 19613 13889 19625 13892
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 20438 13880 20444 13932
rect 20496 13880 20502 13932
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13920 20591 13923
rect 22370 13920 22376 13932
rect 20579 13892 22376 13920
rect 20579 13889 20591 13892
rect 20533 13883 20591 13889
rect 22370 13880 22376 13892
rect 22428 13880 22434 13932
rect 22554 13880 22560 13932
rect 22612 13920 22618 13932
rect 23860 13929 23888 13960
rect 24578 13948 24584 14000
rect 24636 13988 24642 14000
rect 25041 13991 25099 13997
rect 25041 13988 25053 13991
rect 24636 13960 25053 13988
rect 24636 13948 24642 13960
rect 25041 13957 25053 13960
rect 25087 13957 25099 13991
rect 25041 13951 25099 13957
rect 25130 13948 25136 14000
rect 25188 13988 25194 14000
rect 25593 13991 25651 13997
rect 25593 13988 25605 13991
rect 25188 13960 25605 13988
rect 25188 13948 25194 13960
rect 25593 13957 25605 13960
rect 25639 13957 25651 13991
rect 25593 13951 25651 13957
rect 23753 13923 23811 13929
rect 23753 13920 23765 13923
rect 22612 13892 23765 13920
rect 22612 13880 22618 13892
rect 23753 13889 23765 13892
rect 23799 13889 23811 13923
rect 23753 13883 23811 13889
rect 23845 13923 23903 13929
rect 23845 13889 23857 13923
rect 23891 13920 23903 13923
rect 24118 13920 24124 13932
rect 23891 13892 24124 13920
rect 23891 13889 23903 13892
rect 23845 13883 23903 13889
rect 17828 13824 18644 13852
rect 17828 13812 17834 13824
rect 18782 13812 18788 13864
rect 18840 13852 18846 13864
rect 20346 13852 20352 13864
rect 18840 13824 20352 13852
rect 18840 13812 18846 13824
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 20717 13855 20775 13861
rect 20717 13821 20729 13855
rect 20763 13821 20775 13855
rect 20717 13815 20775 13821
rect 19242 13744 19248 13796
rect 19300 13784 19306 13796
rect 19300 13756 20208 13784
rect 19300 13744 19306 13756
rect 14458 13716 14464 13728
rect 13372 13688 14464 13716
rect 10744 13676 10750 13688
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 16666 13676 16672 13728
rect 16724 13676 16730 13728
rect 17402 13725 17408 13728
rect 17392 13719 17408 13725
rect 17392 13685 17404 13719
rect 17392 13679 17408 13685
rect 17402 13676 17408 13679
rect 17460 13676 17466 13728
rect 20180 13716 20208 13756
rect 20622 13744 20628 13796
rect 20680 13784 20686 13796
rect 20732 13784 20760 13815
rect 20990 13812 20996 13864
rect 21048 13852 21054 13864
rect 22833 13855 22891 13861
rect 21048 13824 22232 13852
rect 21048 13812 21054 13824
rect 22204 13793 22232 13824
rect 22833 13821 22845 13855
rect 22879 13821 22891 13855
rect 23768 13852 23796 13883
rect 24118 13880 24124 13892
rect 24176 13880 24182 13932
rect 25314 13880 25320 13932
rect 25372 13920 25378 13932
rect 25777 13923 25835 13929
rect 25777 13920 25789 13923
rect 25372 13892 25789 13920
rect 25372 13880 25378 13892
rect 25777 13889 25789 13892
rect 25823 13889 25835 13923
rect 25777 13883 25835 13889
rect 23768 13824 23888 13852
rect 22833 13815 22891 13821
rect 22189 13787 22247 13793
rect 20680 13756 20760 13784
rect 20824 13756 22094 13784
rect 20680 13744 20686 13756
rect 20824 13716 20852 13756
rect 20180 13688 20852 13716
rect 22066 13716 22094 13756
rect 22189 13753 22201 13787
rect 22235 13753 22247 13787
rect 22189 13747 22247 13753
rect 22738 13744 22744 13796
rect 22796 13784 22802 13796
rect 22848 13784 22876 13815
rect 23750 13784 23756 13796
rect 22796 13756 23756 13784
rect 22796 13744 22802 13756
rect 23750 13744 23756 13756
rect 23808 13744 23814 13796
rect 23860 13784 23888 13824
rect 24026 13812 24032 13864
rect 24084 13812 24090 13864
rect 25130 13812 25136 13864
rect 25188 13852 25194 13864
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 25188 13824 25237 13852
rect 25188 13812 25194 13824
rect 25225 13821 25237 13824
rect 25271 13852 25283 13855
rect 26145 13855 26203 13861
rect 26145 13852 26157 13855
rect 25271 13824 26157 13852
rect 25271 13821 25283 13824
rect 25225 13815 25283 13821
rect 26145 13821 26157 13824
rect 26191 13821 26203 13855
rect 26145 13815 26203 13821
rect 25961 13787 26019 13793
rect 25961 13784 25973 13787
rect 23860 13756 25973 13784
rect 25961 13753 25973 13756
rect 26007 13753 26019 13787
rect 25961 13747 26019 13753
rect 22830 13716 22836 13728
rect 22066 13688 22836 13716
rect 22830 13676 22836 13688
rect 22888 13676 22894 13728
rect 24578 13676 24584 13728
rect 24636 13676 24642 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 3421 13515 3479 13521
rect 3421 13481 3433 13515
rect 3467 13512 3479 13515
rect 4246 13512 4252 13524
rect 3467 13484 4252 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 4246 13472 4252 13484
rect 4304 13512 4310 13524
rect 4614 13512 4620 13524
rect 4304 13484 4620 13512
rect 4304 13472 4310 13484
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 7432 13484 8064 13512
rect 7432 13472 7438 13484
rect 5442 13404 5448 13456
rect 5500 13444 5506 13456
rect 6365 13447 6423 13453
rect 6365 13444 6377 13447
rect 5500 13416 6377 13444
rect 5500 13404 5506 13416
rect 6365 13413 6377 13416
rect 6411 13413 6423 13447
rect 8036 13444 8064 13484
rect 9030 13472 9036 13524
rect 9088 13512 9094 13524
rect 14366 13512 14372 13524
rect 9088 13484 14372 13512
rect 9088 13472 9094 13484
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 15010 13472 15016 13524
rect 15068 13512 15074 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15068 13484 16037 13512
rect 15068 13472 15074 13484
rect 16025 13481 16037 13484
rect 16071 13481 16083 13515
rect 16025 13475 16083 13481
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 17460 13484 18889 13512
rect 17460 13472 17466 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 20346 13472 20352 13524
rect 20404 13512 20410 13524
rect 22097 13515 22155 13521
rect 20404 13484 21680 13512
rect 20404 13472 20410 13484
rect 10686 13444 10692 13456
rect 8036 13416 10692 13444
rect 6365 13407 6423 13413
rect 2038 13336 2044 13388
rect 2096 13336 2102 13388
rect 4157 13379 4215 13385
rect 4157 13345 4169 13379
rect 4203 13376 4215 13379
rect 5166 13376 5172 13388
rect 4203 13348 5172 13376
rect 4203 13345 4215 13348
rect 4157 13339 4215 13345
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 1762 13268 1768 13320
rect 1820 13268 1826 13320
rect 5534 13268 5540 13320
rect 5592 13268 5598 13320
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 6181 13311 6239 13317
rect 6181 13308 6193 13311
rect 5868 13280 6193 13308
rect 5868 13268 5874 13280
rect 6181 13277 6193 13280
rect 6227 13277 6239 13311
rect 6181 13271 6239 13277
rect 4430 13200 4436 13252
rect 4488 13200 4494 13252
rect 4522 13200 4528 13252
rect 4580 13240 4586 13252
rect 4580 13212 4922 13240
rect 4580 13200 4586 13212
rect 1854 13132 1860 13184
rect 1912 13172 1918 13184
rect 3513 13175 3571 13181
rect 3513 13172 3525 13175
rect 1912 13144 3525 13172
rect 1912 13132 1918 13144
rect 3513 13141 3525 13144
rect 3559 13172 3571 13175
rect 3786 13172 3792 13184
rect 3559 13144 3792 13172
rect 3559 13141 3571 13144
rect 3513 13135 3571 13141
rect 3786 13132 3792 13144
rect 3844 13132 3850 13184
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 4706 13172 4712 13184
rect 3927 13144 4712 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 4816 13172 4844 13212
rect 5552 13172 5580 13268
rect 5828 13212 6224 13240
rect 5828 13172 5856 13212
rect 6196 13184 6224 13212
rect 4816 13144 5856 13172
rect 5902 13132 5908 13184
rect 5960 13132 5966 13184
rect 6178 13132 6184 13184
rect 6236 13132 6242 13184
rect 6380 13172 6408 13407
rect 10686 13404 10692 13416
rect 10744 13404 10750 13456
rect 11514 13404 11520 13456
rect 11572 13404 11578 13456
rect 11701 13447 11759 13453
rect 11701 13413 11713 13447
rect 11747 13444 11759 13447
rect 11790 13444 11796 13456
rect 11747 13416 11796 13444
rect 11747 13413 11759 13416
rect 11701 13407 11759 13413
rect 6733 13379 6791 13385
rect 6733 13345 6745 13379
rect 6779 13376 6791 13379
rect 7466 13376 7472 13388
rect 6779 13348 7472 13376
rect 6779 13345 6791 13348
rect 6733 13339 6791 13345
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 8478 13336 8484 13388
rect 8536 13336 8542 13388
rect 9030 13336 9036 13388
rect 9088 13376 9094 13388
rect 9125 13379 9183 13385
rect 9125 13376 9137 13379
rect 9088 13348 9137 13376
rect 9088 13336 9094 13348
rect 9125 13345 9137 13348
rect 9171 13345 9183 13379
rect 9125 13339 9183 13345
rect 9398 13336 9404 13388
rect 9456 13336 9462 13388
rect 10870 13336 10876 13388
rect 10928 13336 10934 13388
rect 10965 13379 11023 13385
rect 10965 13345 10977 13379
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 8496 13308 8524 13336
rect 10980 13308 11008 13339
rect 11238 13336 11244 13388
rect 11296 13376 11302 13388
rect 11716 13376 11744 13407
rect 11790 13404 11796 13416
rect 11848 13404 11854 13456
rect 13722 13404 13728 13456
rect 13780 13404 13786 13456
rect 21652 13444 21680 13484
rect 22097 13481 22109 13515
rect 22143 13512 22155 13515
rect 22186 13512 22192 13524
rect 22143 13484 22192 13512
rect 22143 13481 22155 13484
rect 22097 13475 22155 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 22554 13472 22560 13524
rect 22612 13472 22618 13524
rect 23290 13472 23296 13524
rect 23348 13512 23354 13524
rect 23934 13512 23940 13524
rect 23348 13484 23940 13512
rect 23348 13472 23354 13484
rect 23934 13472 23940 13484
rect 23992 13472 23998 13524
rect 24118 13472 24124 13524
rect 24176 13472 24182 13524
rect 32490 13512 32496 13524
rect 31726 13484 32496 13512
rect 21652 13416 22784 13444
rect 11296 13348 11744 13376
rect 11296 13336 11302 13348
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 14553 13379 14611 13385
rect 12032 13348 14320 13376
rect 12032 13336 12038 13348
rect 14292 13320 14320 13348
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15194 13376 15200 13388
rect 14599 13348 15200 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 15194 13336 15200 13348
rect 15252 13376 15258 13388
rect 16390 13376 16396 13388
rect 15252 13348 16396 13376
rect 15252 13336 15258 13348
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 17126 13336 17132 13388
rect 17184 13376 17190 13388
rect 17494 13376 17500 13388
rect 17184 13348 17500 13376
rect 17184 13336 17190 13348
rect 17494 13336 17500 13348
rect 17552 13376 17558 13388
rect 20070 13376 20076 13388
rect 17552 13348 20076 13376
rect 17552 13336 17558 13348
rect 20070 13336 20076 13348
rect 20128 13336 20134 13388
rect 20349 13379 20407 13385
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 22186 13376 22192 13388
rect 20395 13348 22192 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 22186 13336 22192 13348
rect 22244 13336 22250 13388
rect 22756 13376 22784 13416
rect 22830 13404 22836 13456
rect 22888 13444 22894 13456
rect 31726 13444 31754 13484
rect 32490 13472 32496 13484
rect 32548 13472 32554 13524
rect 22888 13416 31754 13444
rect 22888 13404 22894 13416
rect 23474 13376 23480 13388
rect 22756 13348 23480 13376
rect 23474 13336 23480 13348
rect 23532 13336 23538 13388
rect 23750 13336 23756 13388
rect 23808 13376 23814 13388
rect 24670 13376 24676 13388
rect 23808 13348 24676 13376
rect 23808 13336 23814 13348
rect 24670 13336 24676 13348
rect 24728 13336 24734 13388
rect 13998 13308 14004 13320
rect 8496 13280 11008 13308
rect 13386 13280 14004 13308
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 23014 13268 23020 13320
rect 23072 13308 23078 13320
rect 23072 13280 25452 13308
rect 23072 13268 23078 13280
rect 7006 13200 7012 13252
rect 7064 13200 7070 13252
rect 7098 13200 7104 13252
rect 7156 13240 7162 13252
rect 9674 13240 9680 13252
rect 7156 13212 7498 13240
rect 7156 13200 7162 13212
rect 9646 13200 9680 13240
rect 9732 13240 9738 13252
rect 10781 13243 10839 13249
rect 9732 13212 10548 13240
rect 9732 13200 9738 13212
rect 9646 13172 9674 13200
rect 6380 13144 9674 13172
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 10413 13175 10471 13181
rect 10413 13172 10425 13175
rect 9824 13144 10425 13172
rect 9824 13132 9830 13144
rect 10413 13141 10425 13144
rect 10459 13141 10471 13175
rect 10520 13172 10548 13212
rect 10781 13209 10793 13243
rect 10827 13240 10839 13243
rect 12253 13243 12311 13249
rect 10827 13212 12112 13240
rect 10827 13209 10839 13212
rect 10781 13203 10839 13209
rect 11606 13172 11612 13184
rect 10520 13144 11612 13172
rect 10413 13135 10471 13141
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 12084 13172 12112 13212
rect 12253 13209 12265 13243
rect 12299 13240 12311 13243
rect 12342 13240 12348 13252
rect 12299 13212 12348 13240
rect 12299 13209 12311 13212
rect 12253 13203 12311 13209
rect 12342 13200 12348 13212
rect 12400 13200 12406 13252
rect 13722 13200 13728 13252
rect 13780 13240 13786 13252
rect 14090 13240 14096 13252
rect 13780 13212 14096 13240
rect 13780 13200 13786 13212
rect 14090 13200 14096 13212
rect 14148 13200 14154 13252
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14826 13240 14832 13252
rect 14240 13212 14832 13240
rect 14240 13200 14246 13212
rect 14826 13200 14832 13212
rect 14884 13200 14890 13252
rect 15286 13200 15292 13252
rect 15344 13200 15350 13252
rect 17402 13240 17408 13252
rect 16132 13212 17408 13240
rect 13630 13172 13636 13184
rect 12084 13144 13636 13172
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 16132 13172 16160 13212
rect 17402 13200 17408 13212
rect 17460 13200 17466 13252
rect 17862 13200 17868 13252
rect 17920 13200 17926 13252
rect 18966 13240 18972 13252
rect 18708 13212 18972 13240
rect 13872 13144 16160 13172
rect 13872 13132 13878 13144
rect 16206 13132 16212 13184
rect 16264 13172 16270 13184
rect 18708 13172 18736 13212
rect 18966 13200 18972 13212
rect 19024 13240 19030 13252
rect 20625 13243 20683 13249
rect 20625 13240 20637 13243
rect 19024 13212 20637 13240
rect 19024 13200 19030 13212
rect 20625 13209 20637 13212
rect 20671 13209 20683 13243
rect 20625 13203 20683 13209
rect 21008 13212 21114 13240
rect 16264 13144 18736 13172
rect 19337 13175 19395 13181
rect 16264 13132 16270 13144
rect 19337 13141 19349 13175
rect 19383 13172 19395 13175
rect 19429 13175 19487 13181
rect 19429 13172 19441 13175
rect 19383 13144 19441 13172
rect 19383 13141 19395 13144
rect 19337 13135 19395 13141
rect 19429 13141 19441 13144
rect 19475 13172 19487 13175
rect 21008 13172 21036 13212
rect 22370 13200 22376 13252
rect 22428 13240 22434 13252
rect 22428 13212 22876 13240
rect 22428 13200 22434 13212
rect 21266 13172 21272 13184
rect 19475 13144 21272 13172
rect 19475 13141 19487 13144
rect 19429 13135 19487 13141
rect 21266 13132 21272 13144
rect 21324 13132 21330 13184
rect 22848 13181 22876 13212
rect 23106 13200 23112 13252
rect 23164 13240 23170 13252
rect 23201 13243 23259 13249
rect 23201 13240 23213 13243
rect 23164 13212 23213 13240
rect 23164 13200 23170 13212
rect 23201 13209 23213 13212
rect 23247 13209 23259 13243
rect 23201 13203 23259 13209
rect 23293 13243 23351 13249
rect 23293 13209 23305 13243
rect 23339 13240 23351 13243
rect 23750 13240 23756 13252
rect 23339 13212 23756 13240
rect 23339 13209 23351 13212
rect 23293 13203 23351 13209
rect 23750 13200 23756 13212
rect 23808 13200 23814 13252
rect 23934 13200 23940 13252
rect 23992 13240 23998 13252
rect 25424 13249 25452 13280
rect 24581 13243 24639 13249
rect 24581 13240 24593 13243
rect 23992 13212 24593 13240
rect 23992 13200 23998 13212
rect 24581 13209 24593 13212
rect 24627 13209 24639 13243
rect 24581 13203 24639 13209
rect 25409 13243 25467 13249
rect 25409 13209 25421 13243
rect 25455 13240 25467 13243
rect 27522 13240 27528 13252
rect 25455 13212 27528 13240
rect 25455 13209 25467 13212
rect 25409 13203 25467 13209
rect 27522 13200 27528 13212
rect 27580 13200 27586 13252
rect 22833 13175 22891 13181
rect 22833 13141 22845 13175
rect 22879 13141 22891 13175
rect 22833 13135 22891 13141
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 3602 12928 3608 12980
rect 3660 12928 3666 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 4801 12971 4859 12977
rect 4801 12968 4813 12971
rect 4580 12940 4813 12968
rect 4580 12928 4586 12940
rect 4801 12937 4813 12940
rect 4847 12968 4859 12971
rect 5626 12968 5632 12980
rect 4847 12940 5632 12968
rect 4847 12937 4859 12940
rect 4801 12931 4859 12937
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 5718 12928 5724 12980
rect 5776 12928 5782 12980
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 6236 12940 6469 12968
rect 6236 12928 6242 12940
rect 6457 12937 6469 12940
rect 6503 12968 6515 12971
rect 6822 12968 6828 12980
rect 6503 12940 6828 12968
rect 6503 12937 6515 12940
rect 6457 12931 6515 12937
rect 6822 12928 6828 12940
rect 6880 12968 6886 12980
rect 7098 12968 7104 12980
rect 6880 12940 7104 12968
rect 6880 12928 6886 12940
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 10594 12968 10600 12980
rect 7331 12940 10600 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12529 12971 12587 12977
rect 12529 12968 12541 12971
rect 12492 12940 12541 12968
rect 12492 12928 12498 12940
rect 12529 12937 12541 12940
rect 12575 12937 12587 12971
rect 12529 12931 12587 12937
rect 13725 12971 13783 12977
rect 13725 12937 13737 12971
rect 13771 12968 13783 12971
rect 14550 12968 14556 12980
rect 13771 12940 14556 12968
rect 13771 12937 13783 12940
rect 13725 12931 13783 12937
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 16117 12971 16175 12977
rect 16117 12968 16129 12971
rect 15344 12940 16129 12968
rect 15344 12928 15350 12940
rect 16117 12937 16129 12940
rect 16163 12968 16175 12971
rect 16666 12968 16672 12980
rect 16163 12940 16672 12968
rect 16163 12937 16175 12940
rect 16117 12931 16175 12937
rect 16666 12928 16672 12940
rect 16724 12928 16730 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 17000 12940 17785 12968
rect 17000 12928 17006 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 18141 12971 18199 12977
rect 18141 12937 18153 12971
rect 18187 12968 18199 12971
rect 18782 12968 18788 12980
rect 18187 12940 18788 12968
rect 18187 12937 18199 12940
rect 18141 12931 18199 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 21085 12971 21143 12977
rect 21085 12937 21097 12971
rect 21131 12968 21143 12971
rect 21174 12968 21180 12980
rect 21131 12940 21180 12968
rect 21131 12937 21143 12940
rect 21085 12931 21143 12937
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 21266 12928 21272 12980
rect 21324 12968 21330 12980
rect 22002 12968 22008 12980
rect 21324 12940 22008 12968
rect 21324 12928 21330 12940
rect 22002 12928 22008 12940
rect 22060 12968 22066 12980
rect 22060 12940 22692 12968
rect 22060 12928 22066 12940
rect 2866 12860 2872 12912
rect 2924 12900 2930 12912
rect 3513 12903 3571 12909
rect 3513 12900 3525 12903
rect 2924 12872 3525 12900
rect 2924 12860 2930 12872
rect 3513 12869 3525 12872
rect 3559 12900 3571 12903
rect 3694 12900 3700 12912
rect 3559 12872 3700 12900
rect 3559 12869 3571 12872
rect 3513 12863 3571 12869
rect 3694 12860 3700 12872
rect 3752 12860 3758 12912
rect 3970 12860 3976 12912
rect 4028 12900 4034 12912
rect 4249 12903 4307 12909
rect 4249 12900 4261 12903
rect 4028 12872 4261 12900
rect 4028 12860 4034 12872
rect 4249 12869 4261 12872
rect 4295 12900 4307 12903
rect 4338 12900 4344 12912
rect 4295 12872 4344 12900
rect 4295 12869 4307 12872
rect 4249 12863 4307 12869
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 4430 12860 4436 12912
rect 4488 12900 4494 12912
rect 10318 12900 10324 12912
rect 4488 12872 7420 12900
rect 4488 12860 4494 12872
rect 1210 12792 1216 12844
rect 1268 12832 1274 12844
rect 1581 12835 1639 12841
rect 1581 12832 1593 12835
rect 1268 12804 1593 12832
rect 1268 12792 1274 12804
rect 1581 12801 1593 12804
rect 1627 12801 1639 12835
rect 1581 12795 1639 12801
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 2314 12832 2320 12844
rect 1903 12804 2320 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 2314 12792 2320 12804
rect 2372 12792 2378 12844
rect 2498 12792 2504 12844
rect 2556 12792 2562 12844
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 3878 12832 3884 12844
rect 2823 12804 3884 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 3878 12792 3884 12804
rect 3936 12792 3942 12844
rect 5074 12792 5080 12844
rect 5132 12832 5138 12844
rect 5442 12832 5448 12844
rect 5132 12804 5448 12832
rect 5132 12792 5138 12804
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 5626 12792 5632 12844
rect 5684 12792 5690 12844
rect 2516 12764 2544 12792
rect 2240 12736 2544 12764
rect 4433 12767 4491 12773
rect 2240 12640 2268 12736
rect 4433 12733 4445 12767
rect 4479 12764 4491 12767
rect 5350 12764 5356 12776
rect 4479 12736 5356 12764
rect 4479 12733 4491 12736
rect 4433 12727 4491 12733
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 6012 12764 6040 12872
rect 7193 12835 7251 12841
rect 7193 12801 7205 12835
rect 7239 12832 7251 12835
rect 7282 12832 7288 12844
rect 7239 12804 7288 12832
rect 7239 12801 7251 12804
rect 7193 12795 7251 12801
rect 5951 12736 6040 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 2498 12656 2504 12708
rect 2556 12696 2562 12708
rect 3145 12699 3203 12705
rect 3145 12696 3157 12699
rect 2556 12668 3157 12696
rect 2556 12656 2562 12668
rect 3145 12665 3157 12668
rect 3191 12696 3203 12699
rect 7208 12696 7236 12795
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 7392 12773 7420 12872
rect 9646 12872 10324 12900
rect 9398 12792 9404 12844
rect 9456 12792 9462 12844
rect 7377 12767 7435 12773
rect 7377 12733 7389 12767
rect 7423 12733 7435 12767
rect 7377 12727 7435 12733
rect 7466 12724 7472 12776
rect 7524 12764 7530 12776
rect 8021 12767 8079 12773
rect 8021 12764 8033 12767
rect 7524 12736 8033 12764
rect 7524 12724 7530 12736
rect 8021 12733 8033 12736
rect 8067 12733 8079 12767
rect 8021 12727 8079 12733
rect 3191 12668 7236 12696
rect 3191 12665 3203 12668
rect 3145 12659 3203 12665
rect 8036 12640 8064 12727
rect 8294 12724 8300 12776
rect 8352 12724 8358 12776
rect 9416 12764 9444 12792
rect 9646 12764 9674 12872
rect 10318 12860 10324 12872
rect 10376 12900 10382 12912
rect 11333 12903 11391 12909
rect 11333 12900 11345 12903
rect 10376 12872 11345 12900
rect 10376 12860 10382 12872
rect 11333 12869 11345 12872
rect 11379 12869 11391 12903
rect 11333 12863 11391 12869
rect 11885 12903 11943 12909
rect 11885 12869 11897 12903
rect 11931 12900 11943 12903
rect 13630 12900 13636 12912
rect 11931 12872 13636 12900
rect 11931 12869 11943 12872
rect 11885 12863 11943 12869
rect 13630 12860 13636 12872
rect 13688 12860 13694 12912
rect 13814 12860 13820 12912
rect 13872 12900 13878 12912
rect 14274 12900 14280 12912
rect 13872 12872 14280 12900
rect 13872 12860 13878 12872
rect 14274 12860 14280 12872
rect 14332 12900 14338 12912
rect 15657 12903 15715 12909
rect 15657 12900 15669 12903
rect 14332 12872 15669 12900
rect 14332 12860 14338 12872
rect 15657 12869 15669 12872
rect 15703 12869 15715 12903
rect 18414 12900 18420 12912
rect 15657 12863 15715 12869
rect 16316 12872 18420 12900
rect 9950 12792 9956 12844
rect 10008 12832 10014 12844
rect 10686 12832 10692 12844
rect 10008 12804 10692 12832
rect 10008 12792 10014 12804
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 12406 12804 12909 12832
rect 9416 12736 9674 12764
rect 10042 12724 10048 12776
rect 10100 12724 10106 12776
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 12406 12764 12434 12804
rect 12897 12801 12909 12804
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 13446 12832 13452 12844
rect 13136 12804 13452 12832
rect 13136 12792 13142 12804
rect 13446 12792 13452 12804
rect 13504 12832 13510 12844
rect 14093 12835 14151 12841
rect 14093 12832 14105 12835
rect 13504 12804 14105 12832
rect 13504 12792 13510 12804
rect 14093 12801 14105 12804
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 14734 12792 14740 12844
rect 14792 12832 14798 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14792 12804 14933 12832
rect 14792 12792 14798 12804
rect 14921 12801 14933 12804
rect 14967 12832 14979 12835
rect 15102 12832 15108 12844
rect 14967 12804 15108 12832
rect 14967 12801 14979 12804
rect 14921 12795 14979 12801
rect 15102 12792 15108 12804
rect 15160 12832 15166 12844
rect 16316 12841 16344 12872
rect 18414 12860 18420 12872
rect 18472 12900 18478 12912
rect 18874 12900 18880 12912
rect 18472 12872 18880 12900
rect 18472 12860 18478 12872
rect 18874 12860 18880 12872
rect 18932 12900 18938 12912
rect 18969 12903 19027 12909
rect 18969 12900 18981 12903
rect 18932 12872 18981 12900
rect 18932 12860 18938 12872
rect 18969 12869 18981 12872
rect 19015 12869 19027 12903
rect 22278 12900 22284 12912
rect 18969 12863 19027 12869
rect 20180 12872 22284 12900
rect 16301 12835 16359 12841
rect 16301 12832 16313 12835
rect 15160 12804 16313 12832
rect 15160 12792 15166 12804
rect 16301 12801 16313 12804
rect 16347 12801 16359 12835
rect 16301 12795 16359 12801
rect 17402 12792 17408 12844
rect 17460 12832 17466 12844
rect 18046 12832 18052 12844
rect 17460 12804 18052 12832
rect 17460 12792 17466 12804
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12832 18291 12835
rect 20180 12832 20208 12872
rect 22278 12860 22284 12872
rect 22336 12860 22342 12912
rect 18279 12804 20208 12832
rect 21177 12835 21235 12841
rect 18279 12801 18291 12804
rect 18233 12795 18291 12801
rect 21177 12801 21189 12835
rect 21223 12832 21235 12835
rect 21223 12804 22094 12832
rect 21223 12801 21235 12804
rect 21177 12795 21235 12801
rect 10192 12736 12434 12764
rect 12989 12767 13047 12773
rect 10192 12724 10198 12736
rect 12989 12733 13001 12767
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12764 13231 12767
rect 13219 12736 14136 12764
rect 13219 12733 13231 12736
rect 13173 12727 13231 12733
rect 10502 12656 10508 12708
rect 10560 12656 10566 12708
rect 11149 12699 11207 12705
rect 11149 12665 11161 12699
rect 11195 12696 11207 12699
rect 12250 12696 12256 12708
rect 11195 12668 12256 12696
rect 11195 12665 11207 12668
rect 11149 12659 11207 12665
rect 12250 12656 12256 12668
rect 12308 12656 12314 12708
rect 2222 12588 2228 12640
rect 2280 12588 2286 12640
rect 2958 12588 2964 12640
rect 3016 12628 3022 12640
rect 3510 12628 3516 12640
rect 3016 12600 3516 12628
rect 3016 12588 3022 12600
rect 3510 12588 3516 12600
rect 3568 12628 3574 12640
rect 4614 12628 4620 12640
rect 3568 12600 4620 12628
rect 3568 12588 3574 12600
rect 4614 12588 4620 12600
rect 4672 12628 4678 12640
rect 4893 12631 4951 12637
rect 4893 12628 4905 12631
rect 4672 12600 4905 12628
rect 4672 12588 4678 12600
rect 4893 12597 4905 12600
rect 4939 12597 4951 12631
rect 4893 12591 4951 12597
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5442 12628 5448 12640
rect 5307 12600 5448 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 6822 12588 6828 12640
rect 6880 12588 6886 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7466 12628 7472 12640
rect 6972 12600 7472 12628
rect 6972 12588 6978 12600
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 9306 12628 9312 12640
rect 8076 12600 9312 12628
rect 8076 12588 8082 12600
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 11422 12588 11428 12640
rect 11480 12628 11486 12640
rect 11609 12631 11667 12637
rect 11609 12628 11621 12631
rect 11480 12600 11621 12628
rect 11480 12588 11486 12600
rect 11609 12597 11621 12600
rect 11655 12628 11667 12631
rect 12158 12628 12164 12640
rect 11655 12600 12164 12628
rect 11655 12597 11667 12600
rect 11609 12591 11667 12597
rect 12158 12588 12164 12600
rect 12216 12628 12222 12640
rect 12894 12628 12900 12640
rect 12216 12600 12900 12628
rect 12216 12588 12222 12600
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 13004 12628 13032 12727
rect 14108 12696 14136 12736
rect 14182 12724 14188 12776
rect 14240 12724 14246 12776
rect 14369 12767 14427 12773
rect 14369 12733 14381 12767
rect 14415 12764 14427 12767
rect 15194 12764 15200 12776
rect 14415 12736 15200 12764
rect 14415 12733 14427 12736
rect 14369 12727 14427 12733
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 15286 12724 15292 12776
rect 15344 12764 15350 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 15344 12736 16865 12764
rect 15344 12724 15350 12736
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 18064 12764 18092 12792
rect 18064 12736 18368 12764
rect 16853 12727 16911 12733
rect 15102 12696 15108 12708
rect 14108 12668 15108 12696
rect 15102 12656 15108 12668
rect 15160 12696 15166 12708
rect 15470 12696 15476 12708
rect 15160 12668 15476 12696
rect 15160 12656 15166 12668
rect 15470 12656 15476 12668
rect 15528 12656 15534 12708
rect 18340 12696 18368 12736
rect 18414 12724 18420 12776
rect 18472 12724 18478 12776
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 20070 12764 20076 12776
rect 19843 12736 20076 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 21450 12764 21456 12776
rect 21407 12736 21456 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 22066 12764 22094 12804
rect 22462 12764 22468 12776
rect 22066 12736 22468 12764
rect 22462 12724 22468 12736
rect 22520 12724 22526 12776
rect 22664 12764 22692 12940
rect 22738 12928 22744 12980
rect 22796 12968 22802 12980
rect 23198 12968 23204 12980
rect 22796 12940 23204 12968
rect 22796 12928 22802 12940
rect 23198 12928 23204 12940
rect 23256 12928 23262 12980
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 24765 12971 24823 12977
rect 24765 12968 24777 12971
rect 23532 12940 24777 12968
rect 23532 12928 23538 12940
rect 24765 12937 24777 12940
rect 24811 12937 24823 12971
rect 24765 12931 24823 12937
rect 23293 12903 23351 12909
rect 23293 12869 23305 12903
rect 23339 12900 23351 12903
rect 23566 12900 23572 12912
rect 23339 12872 23572 12900
rect 23339 12869 23351 12872
rect 23293 12863 23351 12869
rect 23566 12860 23572 12872
rect 23624 12860 23630 12912
rect 23842 12860 23848 12912
rect 23900 12860 23906 12912
rect 23014 12792 23020 12844
rect 23072 12792 23078 12844
rect 23842 12764 23848 12776
rect 22664 12736 23848 12764
rect 23842 12724 23848 12736
rect 23900 12724 23906 12776
rect 21726 12696 21732 12708
rect 18340 12668 18460 12696
rect 18322 12628 18328 12640
rect 13004 12600 18328 12628
rect 18322 12588 18328 12600
rect 18380 12588 18386 12640
rect 18432 12628 18460 12668
rect 19306 12668 21732 12696
rect 19306 12628 19334 12668
rect 21726 12656 21732 12668
rect 21784 12656 21790 12708
rect 24394 12656 24400 12708
rect 24452 12696 24458 12708
rect 25041 12699 25099 12705
rect 25041 12696 25053 12699
rect 24452 12668 25053 12696
rect 24452 12656 24458 12668
rect 25041 12665 25053 12668
rect 25087 12665 25099 12699
rect 25041 12659 25099 12665
rect 18432 12600 19334 12628
rect 20717 12631 20775 12637
rect 20717 12597 20729 12631
rect 20763 12628 20775 12631
rect 20898 12628 20904 12640
rect 20763 12600 20904 12628
rect 20763 12597 20775 12600
rect 20717 12591 20775 12597
rect 20898 12588 20904 12600
rect 20956 12588 20962 12640
rect 22002 12588 22008 12640
rect 22060 12628 22066 12640
rect 22189 12631 22247 12637
rect 22189 12628 22201 12631
rect 22060 12600 22201 12628
rect 22060 12588 22066 12600
rect 22189 12597 22201 12600
rect 22235 12597 22247 12631
rect 22189 12591 22247 12597
rect 22278 12588 22284 12640
rect 22336 12628 22342 12640
rect 23014 12628 23020 12640
rect 22336 12600 23020 12628
rect 22336 12588 22342 12600
rect 23014 12588 23020 12600
rect 23072 12588 23078 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 3326 12384 3332 12436
rect 3384 12424 3390 12436
rect 3786 12424 3792 12436
rect 3384 12396 3792 12424
rect 3384 12384 3390 12396
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 3970 12384 3976 12436
rect 4028 12384 4034 12436
rect 4617 12427 4675 12433
rect 4617 12393 4629 12427
rect 4663 12424 4675 12427
rect 7742 12424 7748 12436
rect 4663 12396 7748 12424
rect 4663 12393 4675 12396
rect 4617 12387 4675 12393
rect 3145 12359 3203 12365
rect 3145 12325 3157 12359
rect 3191 12356 3203 12359
rect 4154 12356 4160 12368
rect 3191 12328 4160 12356
rect 3191 12325 3203 12328
rect 3145 12319 3203 12325
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12288 1915 12291
rect 1903 12260 2774 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 1486 12180 1492 12232
rect 1544 12220 1550 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1544 12192 1593 12220
rect 1544 12180 1550 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 2746 12152 2774 12260
rect 3418 12248 3424 12300
rect 3476 12288 3482 12300
rect 3970 12288 3976 12300
rect 3476 12260 3976 12288
rect 3476 12248 3482 12260
rect 3970 12248 3976 12260
rect 4028 12248 4034 12300
rect 4724 12297 4752 12396
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 7837 12427 7895 12433
rect 7837 12393 7849 12427
rect 7883 12424 7895 12427
rect 10870 12424 10876 12436
rect 7883 12396 10876 12424
rect 7883 12393 7895 12396
rect 7837 12387 7895 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 11793 12427 11851 12433
rect 11793 12393 11805 12427
rect 11839 12424 11851 12427
rect 12526 12424 12532 12436
rect 11839 12396 12532 12424
rect 11839 12393 11851 12396
rect 11793 12387 11851 12393
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 13035 12396 17632 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 7006 12316 7012 12368
rect 7064 12356 7070 12368
rect 7064 12328 7604 12356
rect 7064 12316 7070 12328
rect 4709 12291 4767 12297
rect 4709 12257 4721 12291
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 5166 12248 5172 12300
rect 5224 12288 5230 12300
rect 5353 12291 5411 12297
rect 5353 12288 5365 12291
rect 5224 12260 5365 12288
rect 5224 12248 5230 12260
rect 5353 12257 5365 12260
rect 5399 12288 5411 12291
rect 6086 12288 6092 12300
rect 5399 12260 6092 12288
rect 5399 12257 5411 12260
rect 5353 12251 5411 12257
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 6178 12248 6184 12300
rect 6236 12288 6242 12300
rect 7377 12291 7435 12297
rect 6236 12260 6684 12288
rect 6236 12248 6242 12260
rect 2958 12180 2964 12232
rect 3016 12180 3022 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4246 12220 4252 12232
rect 4203 12192 4252 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 4246 12180 4252 12192
rect 4304 12180 4310 12232
rect 6656 12164 6684 12260
rect 7377 12257 7389 12291
rect 7423 12288 7435 12291
rect 7466 12288 7472 12300
rect 7423 12260 7472 12288
rect 7423 12257 7435 12260
rect 7377 12251 7435 12257
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 7576 12288 7604 12328
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 15286 12356 15292 12368
rect 13780 12328 15292 12356
rect 13780 12316 13786 12328
rect 15286 12316 15292 12328
rect 15344 12316 15350 12368
rect 15470 12316 15476 12368
rect 15528 12316 15534 12368
rect 17604 12356 17632 12396
rect 18046 12384 18052 12436
rect 18104 12384 18110 12436
rect 18874 12384 18880 12436
rect 18932 12384 18938 12436
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21821 12427 21879 12433
rect 21821 12424 21833 12427
rect 20772 12396 21833 12424
rect 20772 12384 20778 12396
rect 21821 12393 21833 12396
rect 21867 12424 21879 12427
rect 21910 12424 21916 12436
rect 21867 12396 21916 12424
rect 21867 12393 21879 12396
rect 21821 12387 21879 12393
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 25590 12424 25596 12436
rect 22066 12396 25596 12424
rect 19426 12356 19432 12368
rect 17604 12328 19432 12356
rect 19426 12316 19432 12328
rect 19484 12316 19490 12368
rect 22066 12356 22094 12396
rect 25590 12384 25596 12396
rect 25648 12384 25654 12436
rect 19536 12328 20208 12356
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 7576 12260 8401 12288
rect 8389 12257 8401 12260
rect 8435 12257 8447 12291
rect 8389 12251 8447 12257
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 9364 12260 9873 12288
rect 9364 12248 9370 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12288 11299 12291
rect 12066 12288 12072 12300
rect 11287 12260 12072 12288
rect 11287 12257 11299 12260
rect 11241 12251 11299 12257
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12250 12248 12256 12300
rect 12308 12248 12314 12300
rect 12342 12248 12348 12300
rect 12400 12248 12406 12300
rect 13633 12291 13691 12297
rect 13280 12260 13492 12288
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 10410 12220 10416 12232
rect 8343 12192 10416 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 10965 12223 11023 12229
rect 10965 12220 10977 12223
rect 10520 12192 10977 12220
rect 5629 12155 5687 12161
rect 2746 12124 3648 12152
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 3513 12087 3571 12093
rect 3513 12084 3525 12087
rect 3476 12056 3525 12084
rect 3476 12044 3482 12056
rect 3513 12053 3525 12056
rect 3559 12053 3571 12087
rect 3620 12084 3648 12124
rect 5629 12121 5641 12155
rect 5675 12152 5687 12155
rect 5718 12152 5724 12164
rect 5675 12124 5724 12152
rect 5675 12121 5687 12124
rect 5629 12115 5687 12121
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 6638 12112 6644 12164
rect 6696 12112 6702 12164
rect 7742 12112 7748 12164
rect 7800 12152 7806 12164
rect 8018 12152 8024 12164
rect 7800 12124 8024 12152
rect 7800 12112 7806 12124
rect 8018 12112 8024 12124
rect 8076 12112 8082 12164
rect 8386 12112 8392 12164
rect 8444 12152 8450 12164
rect 8570 12152 8576 12164
rect 8444 12124 8576 12152
rect 8444 12112 8450 12124
rect 8570 12112 8576 12124
rect 8628 12112 8634 12164
rect 8662 12112 8668 12164
rect 8720 12152 8726 12164
rect 9030 12152 9036 12164
rect 8720 12124 9036 12152
rect 8720 12112 8726 12124
rect 9030 12112 9036 12124
rect 9088 12112 9094 12164
rect 9122 12112 9128 12164
rect 9180 12112 9186 12164
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 10520 12152 10548 12192
rect 10965 12189 10977 12192
rect 11011 12189 11023 12223
rect 10965 12183 11023 12189
rect 11057 12223 11115 12229
rect 11057 12189 11069 12223
rect 11103 12220 11115 12223
rect 13170 12220 13176 12232
rect 11103 12192 13176 12220
rect 11103 12189 11115 12192
rect 11057 12183 11115 12189
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 9732 12124 10548 12152
rect 9732 12112 9738 12124
rect 11606 12112 11612 12164
rect 11664 12152 11670 12164
rect 13280 12152 13308 12260
rect 13464 12229 13492 12260
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 15194 12288 15200 12300
rect 13679 12260 15200 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 15488 12288 15516 12316
rect 16577 12291 16635 12297
rect 16577 12288 16589 12291
rect 15488 12260 16589 12288
rect 16577 12257 16589 12260
rect 16623 12257 16635 12291
rect 16577 12251 16635 12257
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 19536 12288 19564 12328
rect 16724 12260 19564 12288
rect 16724 12248 16730 12260
rect 19610 12248 19616 12300
rect 19668 12248 19674 12300
rect 20070 12248 20076 12300
rect 20128 12248 20134 12300
rect 20180 12288 20208 12328
rect 21744 12328 22094 12356
rect 20806 12288 20812 12300
rect 20180 12260 20812 12288
rect 20806 12248 20812 12260
rect 20864 12288 20870 12300
rect 21744 12288 21772 12328
rect 20864 12260 21772 12288
rect 20864 12248 20870 12260
rect 21910 12248 21916 12300
rect 21968 12288 21974 12300
rect 22557 12291 22615 12297
rect 22557 12288 22569 12291
rect 21968 12260 22569 12288
rect 21968 12248 21974 12260
rect 22557 12257 22569 12260
rect 22603 12257 22615 12291
rect 22557 12251 22615 12257
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 14458 12180 14464 12232
rect 14516 12220 14522 12232
rect 15473 12223 15531 12229
rect 15473 12220 15485 12223
rect 14516 12192 15485 12220
rect 14516 12180 14522 12192
rect 15473 12189 15485 12192
rect 15519 12220 15531 12223
rect 16301 12223 16359 12229
rect 16301 12220 16313 12223
rect 15519 12192 16313 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 16301 12189 16313 12192
rect 16347 12189 16359 12223
rect 16301 12183 16359 12189
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 22281 12223 22339 12229
rect 22281 12220 22293 12223
rect 22244 12192 22293 12220
rect 22244 12180 22250 12192
rect 22281 12189 22293 12192
rect 22327 12189 22339 12223
rect 22281 12183 22339 12189
rect 11664 12124 13308 12152
rect 13357 12155 13415 12161
rect 11664 12112 11670 12124
rect 13357 12121 13369 12155
rect 13403 12152 13415 12155
rect 13722 12152 13728 12164
rect 13403 12124 13728 12152
rect 13403 12121 13415 12124
rect 13357 12115 13415 12121
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 14734 12112 14740 12164
rect 14792 12112 14798 12164
rect 14826 12112 14832 12164
rect 14884 12152 14890 12164
rect 16666 12152 16672 12164
rect 14884 12124 16672 12152
rect 14884 12112 14890 12124
rect 16666 12112 16672 12124
rect 16724 12112 16730 12164
rect 16868 12124 17066 12152
rect 4338 12084 4344 12096
rect 3620 12056 4344 12084
rect 3513 12047 3571 12053
rect 4338 12044 4344 12056
rect 4396 12084 4402 12096
rect 6270 12084 6276 12096
rect 4396 12056 6276 12084
rect 4396 12044 4402 12056
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 7156 12056 8217 12084
rect 7156 12044 7162 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 8205 12047 8263 12053
rect 10594 12044 10600 12096
rect 10652 12044 10658 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 12161 12087 12219 12093
rect 12161 12084 12173 12087
rect 11112 12056 12173 12084
rect 11112 12044 11118 12056
rect 12161 12053 12173 12056
rect 12207 12053 12219 12087
rect 12161 12047 12219 12053
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13906 12084 13912 12096
rect 13228 12056 13912 12084
rect 13228 12044 13234 12056
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 14090 12044 14096 12096
rect 14148 12044 14154 12096
rect 14182 12044 14188 12096
rect 14240 12084 14246 12096
rect 14369 12087 14427 12093
rect 14369 12084 14381 12087
rect 14240 12056 14381 12084
rect 14240 12044 14246 12056
rect 14369 12053 14381 12056
rect 14415 12053 14427 12087
rect 14752 12084 14780 12112
rect 15933 12087 15991 12093
rect 15933 12084 15945 12087
rect 14752 12056 15945 12084
rect 14369 12047 14427 12053
rect 15933 12053 15945 12056
rect 15979 12053 15991 12087
rect 15933 12047 15991 12053
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 16868 12084 16896 12124
rect 17862 12112 17868 12164
rect 17920 12152 17926 12164
rect 18509 12155 18567 12161
rect 18509 12152 18521 12155
rect 17920 12124 18521 12152
rect 17920 12112 17926 12124
rect 18509 12121 18521 12124
rect 18555 12152 18567 12155
rect 18690 12152 18696 12164
rect 18555 12124 18696 12152
rect 18555 12121 18567 12124
rect 18509 12115 18567 12121
rect 18690 12112 18696 12124
rect 18748 12112 18754 12164
rect 18874 12112 18880 12164
rect 18932 12152 18938 12164
rect 18932 12124 19288 12152
rect 18932 12112 18938 12124
rect 18325 12087 18383 12093
rect 18325 12084 18337 12087
rect 16632 12056 18337 12084
rect 16632 12044 16638 12056
rect 18325 12053 18337 12056
rect 18371 12084 18383 12087
rect 18969 12087 19027 12093
rect 18969 12084 18981 12087
rect 18371 12056 18981 12084
rect 18371 12053 18383 12056
rect 18325 12047 18383 12053
rect 18969 12053 18981 12056
rect 19015 12053 19027 12087
rect 19260 12084 19288 12124
rect 20346 12112 20352 12164
rect 20404 12112 20410 12164
rect 21818 12152 21824 12164
rect 21574 12124 21824 12152
rect 21818 12112 21824 12124
rect 21876 12152 21882 12164
rect 23014 12152 23020 12164
rect 21876 12124 23020 12152
rect 21876 12112 21882 12124
rect 23014 12112 23020 12124
rect 23072 12112 23078 12164
rect 19337 12087 19395 12093
rect 19337 12084 19349 12087
rect 19260 12056 19349 12084
rect 18969 12047 19027 12053
rect 19337 12053 19349 12056
rect 19383 12053 19395 12087
rect 19337 12047 19395 12053
rect 24026 12044 24032 12096
rect 24084 12044 24090 12096
rect 24394 12044 24400 12096
rect 24452 12044 24458 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 1489 11883 1547 11889
rect 1489 11849 1501 11883
rect 1535 11880 1547 11883
rect 1762 11880 1768 11892
rect 1535 11852 1768 11880
rect 1535 11849 1547 11852
rect 1489 11843 1547 11849
rect 1762 11840 1768 11852
rect 1820 11840 1826 11892
rect 1857 11883 1915 11889
rect 1857 11849 1869 11883
rect 1903 11880 1915 11883
rect 1946 11880 1952 11892
rect 1903 11852 1952 11880
rect 1903 11849 1915 11852
rect 1857 11843 1915 11849
rect 1946 11840 1952 11852
rect 2004 11840 2010 11892
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 3602 11880 3608 11892
rect 3467 11852 3608 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 4433 11883 4491 11889
rect 4433 11849 4445 11883
rect 4479 11880 4491 11883
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 4479 11852 5273 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 5500 11852 5641 11880
rect 5500 11840 5506 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 5629 11843 5687 11849
rect 6733 11883 6791 11889
rect 6733 11849 6745 11883
rect 6779 11880 6791 11883
rect 6779 11852 9720 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11812 1731 11815
rect 4246 11812 4252 11824
rect 1719 11784 4252 11812
rect 1719 11781 1731 11784
rect 1673 11775 1731 11781
rect 4246 11772 4252 11784
rect 4304 11772 4310 11824
rect 5721 11815 5779 11821
rect 4448 11784 5672 11812
rect 4448 11756 4476 11784
rect 2406 11704 2412 11756
rect 2464 11704 2470 11756
rect 4430 11704 4436 11756
rect 4488 11704 4494 11756
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 5258 11744 5264 11756
rect 4571 11716 5264 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 5644 11744 5672 11784
rect 5721 11781 5733 11815
rect 5767 11812 5779 11815
rect 6822 11812 6828 11824
rect 5767 11784 6828 11812
rect 5767 11781 5779 11784
rect 5721 11775 5779 11781
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 7742 11812 7748 11824
rect 7392 11784 7748 11812
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 5644 11716 6377 11744
rect 6365 11713 6377 11716
rect 6411 11744 6423 11747
rect 6914 11744 6920 11756
rect 6411 11716 6920 11744
rect 6411 11713 6423 11716
rect 6365 11707 6423 11713
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 7392 11753 7420 11784
rect 7742 11772 7748 11784
rect 7800 11772 7806 11824
rect 8202 11772 8208 11824
rect 8260 11772 8266 11824
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 1946 11636 1952 11688
rect 2004 11676 2010 11688
rect 2133 11679 2191 11685
rect 2133 11676 2145 11679
rect 2004 11648 2145 11676
rect 2004 11636 2010 11648
rect 2133 11645 2145 11648
rect 2179 11645 2191 11679
rect 2133 11639 2191 11645
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11645 4767 11679
rect 4709 11639 4767 11645
rect 4724 11608 4752 11639
rect 5166 11636 5172 11688
rect 5224 11676 5230 11688
rect 5813 11679 5871 11685
rect 5813 11676 5825 11679
rect 5224 11648 5825 11676
rect 5224 11636 5230 11648
rect 5813 11645 5825 11648
rect 5859 11676 5871 11679
rect 5902 11676 5908 11688
rect 5859 11648 5908 11676
rect 5859 11645 5871 11648
rect 5813 11639 5871 11645
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 6086 11636 6092 11688
rect 6144 11676 6150 11688
rect 7392 11676 7420 11707
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 9180 11716 9597 11744
rect 9180 11704 9186 11716
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 9692 11744 9720 11852
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 12437 11883 12495 11889
rect 12437 11880 12449 11883
rect 10652 11852 12449 11880
rect 10652 11840 10658 11852
rect 12437 11849 12449 11852
rect 12483 11849 12495 11883
rect 13814 11880 13820 11892
rect 12437 11843 12495 11849
rect 13188 11852 13820 11880
rect 9858 11772 9864 11824
rect 9916 11812 9922 11824
rect 10502 11812 10508 11824
rect 9916 11784 10508 11812
rect 9916 11772 9922 11784
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 11606 11772 11612 11824
rect 11664 11772 11670 11824
rect 11790 11772 11796 11824
rect 11848 11812 11854 11824
rect 11848 11784 12572 11812
rect 11848 11772 11854 11784
rect 12345 11747 12403 11753
rect 12345 11744 12357 11747
rect 9692 11716 12357 11744
rect 9585 11707 9643 11713
rect 12345 11713 12357 11716
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 6144 11648 7420 11676
rect 7653 11679 7711 11685
rect 6144 11636 6150 11648
rect 7653 11645 7665 11679
rect 7699 11676 7711 11679
rect 8386 11676 8392 11688
rect 7699 11648 8392 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 9858 11636 9864 11688
rect 9916 11676 9922 11688
rect 12544 11685 12572 11784
rect 13188 11753 13216 11852
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 15562 11840 15568 11892
rect 15620 11840 15626 11892
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 17862 11880 17868 11892
rect 17368 11852 17868 11880
rect 17368 11840 17374 11852
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 18141 11883 18199 11889
rect 18141 11849 18153 11883
rect 18187 11880 18199 11883
rect 18322 11880 18328 11892
rect 18187 11852 18328 11880
rect 18187 11849 18199 11852
rect 18141 11843 18199 11849
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 20898 11880 20904 11892
rect 19260 11852 20904 11880
rect 15197 11815 15255 11821
rect 15197 11812 15209 11815
rect 14674 11784 15209 11812
rect 15197 11781 15209 11784
rect 15243 11812 15255 11815
rect 15470 11812 15476 11824
rect 15243 11784 15476 11812
rect 15243 11781 15255 11784
rect 15197 11775 15255 11781
rect 15470 11772 15476 11784
rect 15528 11772 15534 11824
rect 17126 11772 17132 11824
rect 17184 11812 17190 11824
rect 18509 11815 18567 11821
rect 18509 11812 18521 11815
rect 17184 11784 18521 11812
rect 17184 11772 17190 11784
rect 18509 11781 18521 11784
rect 18555 11812 18567 11815
rect 19153 11815 19211 11821
rect 19153 11812 19165 11815
rect 18555 11784 19165 11812
rect 18555 11781 18567 11784
rect 18509 11775 18567 11781
rect 19153 11781 19165 11784
rect 19199 11781 19211 11815
rect 19153 11775 19211 11781
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 15930 11704 15936 11756
rect 15988 11704 15994 11756
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11744 16083 11747
rect 19260 11744 19288 11852
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 24026 11880 24032 11892
rect 22066 11852 24032 11880
rect 21818 11812 21824 11824
rect 21206 11784 21824 11812
rect 21818 11772 21824 11784
rect 21876 11772 21882 11824
rect 16071 11716 19288 11744
rect 16071 11713 16083 11716
rect 16025 11707 16083 11713
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 9916 11648 10333 11676
rect 9916 11636 9922 11648
rect 10321 11645 10333 11648
rect 10367 11645 10379 11679
rect 10321 11639 10379 11645
rect 10965 11679 11023 11685
rect 10965 11645 10977 11679
rect 11011 11676 11023 11679
rect 12529 11679 12587 11685
rect 11011 11648 12434 11676
rect 11011 11645 11023 11648
rect 10965 11639 11023 11645
rect 4724 11580 5764 11608
rect 5736 11552 5764 11580
rect 8662 11568 8668 11620
rect 8720 11608 8726 11620
rect 10226 11608 10232 11620
rect 8720 11580 10232 11608
rect 8720 11568 8726 11580
rect 10226 11568 10232 11580
rect 10284 11568 10290 11620
rect 12406 11608 12434 11648
rect 12529 11645 12541 11679
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11676 13507 11679
rect 15010 11676 15016 11688
rect 13495 11648 15016 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 16209 11679 16267 11685
rect 16209 11645 16221 11679
rect 16255 11676 16267 11679
rect 17034 11676 17040 11688
rect 16255 11648 17040 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 17034 11636 17040 11648
rect 17092 11636 17098 11688
rect 17405 11679 17463 11685
rect 17405 11645 17417 11679
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 13170 11608 13176 11620
rect 12406 11580 13176 11608
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 14550 11568 14556 11620
rect 14608 11608 14614 11620
rect 17420 11608 17448 11639
rect 17586 11636 17592 11688
rect 17644 11636 17650 11688
rect 18598 11636 18604 11688
rect 18656 11636 18662 11688
rect 18690 11636 18696 11688
rect 18748 11636 18754 11688
rect 19702 11636 19708 11688
rect 19760 11636 19766 11688
rect 19981 11679 20039 11685
rect 19981 11645 19993 11679
rect 20027 11676 20039 11679
rect 22066 11676 22094 11852
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 22649 11815 22707 11821
rect 22649 11781 22661 11815
rect 22695 11812 22707 11815
rect 22738 11812 22744 11824
rect 22695 11784 22744 11812
rect 22695 11781 22707 11784
rect 22649 11775 22707 11781
rect 22738 11772 22744 11784
rect 22796 11772 22802 11824
rect 23106 11772 23112 11824
rect 23164 11772 23170 11824
rect 20027 11648 22094 11676
rect 20027 11645 20039 11648
rect 19981 11639 20039 11645
rect 22186 11636 22192 11688
rect 22244 11676 22250 11688
rect 22373 11679 22431 11685
rect 22373 11676 22385 11679
rect 22244 11648 22385 11676
rect 22244 11636 22250 11648
rect 22373 11645 22385 11648
rect 22419 11645 22431 11679
rect 23658 11676 23664 11688
rect 22373 11639 22431 11645
rect 22480 11648 23664 11676
rect 19610 11608 19616 11620
rect 14608 11580 19616 11608
rect 14608 11568 14614 11580
rect 19610 11568 19616 11580
rect 19668 11568 19674 11620
rect 22480 11608 22508 11648
rect 23658 11636 23664 11648
rect 23716 11636 23722 11688
rect 24394 11608 24400 11620
rect 21008 11580 22508 11608
rect 23676 11580 24400 11608
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 5258 11540 5264 11552
rect 4111 11512 5264 11540
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 5718 11500 5724 11552
rect 5776 11500 5782 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 8352 11512 9137 11540
rect 8352 11500 8358 11512
rect 9125 11509 9137 11512
rect 9171 11540 9183 11543
rect 9398 11540 9404 11552
rect 9171 11512 9404 11540
rect 9171 11509 9183 11512
rect 9125 11503 9183 11509
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 10318 11540 10324 11552
rect 9548 11512 10324 11540
rect 9548 11500 9554 11512
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 11974 11500 11980 11552
rect 12032 11500 12038 11552
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 14921 11543 14979 11549
rect 14921 11540 14933 11543
rect 12124 11512 14933 11540
rect 12124 11500 12130 11512
rect 14921 11509 14933 11512
rect 14967 11509 14979 11543
rect 14921 11503 14979 11509
rect 16942 11500 16948 11552
rect 17000 11500 17006 11552
rect 18598 11500 18604 11552
rect 18656 11540 18662 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 18656 11512 19441 11540
rect 18656 11500 18662 11512
rect 19429 11509 19441 11512
rect 19475 11540 19487 11543
rect 21008 11540 21036 11580
rect 19475 11512 21036 11540
rect 19475 11509 19487 11512
rect 19429 11503 19487 11509
rect 21450 11500 21456 11552
rect 21508 11500 21514 11552
rect 21818 11500 21824 11552
rect 21876 11540 21882 11552
rect 21913 11543 21971 11549
rect 21913 11540 21925 11543
rect 21876 11512 21925 11540
rect 21876 11500 21882 11512
rect 21913 11509 21925 11512
rect 21959 11509 21971 11543
rect 21913 11503 21971 11509
rect 23106 11500 23112 11552
rect 23164 11540 23170 11552
rect 23676 11540 23704 11580
rect 24394 11568 24400 11580
rect 24452 11568 24458 11620
rect 23164 11512 23704 11540
rect 23164 11500 23170 11512
rect 23750 11500 23756 11552
rect 23808 11540 23814 11552
rect 24121 11543 24179 11549
rect 24121 11540 24133 11543
rect 23808 11512 24133 11540
rect 23808 11500 23814 11512
rect 24121 11509 24133 11512
rect 24167 11540 24179 11543
rect 25130 11540 25136 11552
rect 24167 11512 25136 11540
rect 24167 11509 24179 11512
rect 24121 11503 24179 11509
rect 25130 11500 25136 11512
rect 25188 11500 25194 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 3418 11296 3424 11348
rect 3476 11296 3482 11348
rect 3605 11339 3663 11345
rect 3605 11305 3617 11339
rect 3651 11336 3663 11339
rect 3694 11336 3700 11348
rect 3651 11308 3700 11336
rect 3651 11305 3663 11308
rect 3605 11299 3663 11305
rect 3694 11296 3700 11308
rect 3752 11296 3758 11348
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 5776 11308 6561 11336
rect 5776 11296 5782 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 7837 11339 7895 11345
rect 7837 11305 7849 11339
rect 7883 11336 7895 11339
rect 10594 11336 10600 11348
rect 7883 11308 10600 11336
rect 7883 11305 7895 11308
rect 7837 11299 7895 11305
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 11606 11336 11612 11348
rect 11296 11308 11612 11336
rect 11296 11296 11302 11308
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 12400 11308 13277 11336
rect 12400 11296 12406 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 13354 11296 13360 11348
rect 13412 11296 13418 11348
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 13541 11339 13599 11345
rect 13541 11336 13553 11339
rect 13504 11308 13553 11336
rect 13504 11296 13510 11308
rect 13541 11305 13553 11308
rect 13587 11305 13599 11339
rect 14826 11336 14832 11348
rect 13541 11299 13599 11305
rect 14108 11308 14832 11336
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 8662 11268 8668 11280
rect 1627 11240 4108 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11200 2283 11203
rect 2271 11172 2636 11200
rect 2271 11169 2283 11172
rect 2225 11163 2283 11169
rect 1762 11092 1768 11144
rect 1820 11092 1826 11144
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11101 2559 11135
rect 2608 11132 2636 11172
rect 3694 11132 3700 11144
rect 2608 11104 3700 11132
rect 2501 11095 2559 11101
rect 1578 11024 1584 11076
rect 1636 11064 1642 11076
rect 2516 11064 2544 11095
rect 3694 11092 3700 11104
rect 3752 11092 3758 11144
rect 4080 11141 4108 11240
rect 7024 11240 8668 11268
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 6822 11200 6828 11212
rect 4847 11172 6828 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 7024 11209 7052 11240
rect 8662 11228 8668 11240
rect 8720 11228 8726 11280
rect 9398 11228 9404 11280
rect 9456 11268 9462 11280
rect 10321 11271 10379 11277
rect 9456 11240 9720 11268
rect 9456 11228 9462 11240
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11169 7067 11203
rect 7009 11163 7067 11169
rect 7834 11160 7840 11212
rect 7892 11200 7898 11212
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 7892 11172 8309 11200
rect 7892 11160 7898 11172
rect 8297 11169 8309 11172
rect 8343 11169 8355 11203
rect 8297 11163 8355 11169
rect 8478 11160 8484 11212
rect 8536 11160 8542 11212
rect 9214 11160 9220 11212
rect 9272 11200 9278 11212
rect 9692 11209 9720 11240
rect 10321 11237 10333 11271
rect 10367 11268 10379 11271
rect 10870 11268 10876 11280
rect 10367 11240 10876 11268
rect 10367 11237 10379 11240
rect 10321 11231 10379 11237
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 13372 11268 13400 11296
rect 14108 11277 14136 11308
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 15102 11296 15108 11348
rect 15160 11336 15166 11348
rect 16485 11339 16543 11345
rect 16485 11336 16497 11339
rect 15160 11308 16497 11336
rect 15160 11296 15166 11308
rect 16485 11305 16497 11308
rect 16531 11305 16543 11339
rect 16485 11299 16543 11305
rect 18877 11339 18935 11345
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 18966 11336 18972 11348
rect 18923 11308 18972 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 22649 11339 22707 11345
rect 22649 11305 22661 11339
rect 22695 11336 22707 11339
rect 22830 11336 22836 11348
rect 22695 11308 22836 11336
rect 22695 11305 22707 11308
rect 22649 11299 22707 11305
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 31754 11336 31760 11348
rect 31726 11296 31760 11336
rect 31812 11336 31818 11348
rect 32033 11339 32091 11345
rect 32033 11336 32045 11339
rect 31812 11308 32045 11336
rect 31812 11296 31818 11308
rect 32033 11305 32045 11308
rect 32079 11305 32091 11339
rect 32033 11299 32091 11305
rect 14093 11271 14151 11277
rect 14093 11268 14105 11271
rect 13372 11240 14105 11268
rect 14093 11237 14105 11240
rect 14139 11237 14151 11271
rect 14093 11231 14151 11237
rect 9585 11203 9643 11209
rect 9585 11200 9597 11203
rect 9272 11172 9597 11200
rect 9272 11160 9278 11172
rect 9585 11169 9597 11172
rect 9631 11169 9643 11203
rect 9585 11163 9643 11169
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 10778 11160 10784 11212
rect 10836 11160 10842 11212
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 11011 11172 11805 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 11793 11169 11805 11172
rect 11839 11200 11851 11203
rect 13354 11200 13360 11212
rect 11839 11172 13360 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 15010 11160 15016 11212
rect 15068 11200 15074 11212
rect 18690 11200 18696 11212
rect 15068 11172 18696 11200
rect 15068 11160 15074 11172
rect 18690 11160 18696 11172
rect 18748 11160 18754 11212
rect 21818 11160 21824 11212
rect 21876 11200 21882 11212
rect 22925 11203 22983 11209
rect 22925 11200 22937 11203
rect 21876 11172 22937 11200
rect 21876 11160 21882 11172
rect 22925 11169 22937 11172
rect 22971 11169 22983 11203
rect 22925 11163 22983 11169
rect 27522 11160 27528 11212
rect 27580 11200 27586 11212
rect 29733 11203 29791 11209
rect 29733 11200 29745 11203
rect 27580 11172 29745 11200
rect 27580 11160 27586 11172
rect 29733 11169 29745 11172
rect 29779 11169 29791 11203
rect 29733 11163 29791 11169
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 6638 11132 6644 11144
rect 6210 11104 6644 11132
rect 4065 11095 4123 11101
rect 6638 11092 6644 11104
rect 6696 11132 6702 11144
rect 8205 11135 8263 11141
rect 6696 11104 7512 11132
rect 6696 11092 6702 11104
rect 4982 11064 4988 11076
rect 1636 11036 2544 11064
rect 2746 11036 4988 11064
rect 1636 11024 1642 11036
rect 1946 10956 1952 11008
rect 2004 10996 2010 11008
rect 2746 10996 2774 11036
rect 4982 11024 4988 11036
rect 5040 11024 5046 11076
rect 5077 11067 5135 11073
rect 5077 11033 5089 11067
rect 5123 11064 5135 11067
rect 5166 11064 5172 11076
rect 5123 11036 5172 11064
rect 5123 11033 5135 11036
rect 5077 11027 5135 11033
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 7190 11064 7196 11076
rect 6380 11036 7196 11064
rect 2004 10968 2774 10996
rect 4157 10999 4215 11005
rect 2004 10956 2010 10968
rect 4157 10965 4169 10999
rect 4203 10996 4215 10999
rect 6380 10996 6408 11036
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 7484 11073 7512 11104
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 8846 11132 8852 11144
rect 8251 11104 8852 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 8846 11092 8852 11104
rect 8904 11092 8910 11144
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9766 11132 9772 11144
rect 9539 11104 9772 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 11517 11135 11575 11141
rect 11517 11132 11529 11135
rect 9916 11104 11529 11132
rect 9916 11092 9922 11104
rect 11517 11101 11529 11104
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 14458 11092 14464 11144
rect 14516 11132 14522 11144
rect 14737 11135 14795 11141
rect 14737 11132 14749 11135
rect 14516 11104 14749 11132
rect 14516 11092 14522 11104
rect 14737 11101 14749 11104
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 16908 11104 17141 11132
rect 16908 11092 16914 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 18874 11092 18880 11144
rect 18932 11132 18938 11144
rect 19521 11135 19579 11141
rect 19521 11132 19533 11135
rect 18932 11104 19533 11132
rect 18932 11092 18938 11104
rect 19521 11101 19533 11104
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11101 20959 11135
rect 31726 11132 31754 11296
rect 31142 11104 31754 11132
rect 20901 11095 20959 11101
rect 7469 11067 7527 11073
rect 7469 11033 7481 11067
rect 7515 11064 7527 11067
rect 8294 11064 8300 11076
rect 7515 11036 8300 11064
rect 7515 11033 7527 11036
rect 7469 11027 7527 11033
rect 8294 11024 8300 11036
rect 8352 11024 8358 11076
rect 9048 11036 9352 11064
rect 4203 10968 6408 10996
rect 4203 10965 4215 10968
rect 4157 10959 4215 10965
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 9048 10996 9076 11036
rect 7156 10968 9076 10996
rect 9125 10999 9183 11005
rect 7156 10956 7162 10968
rect 9125 10965 9137 10999
rect 9171 10996 9183 10999
rect 9214 10996 9220 11008
rect 9171 10968 9220 10996
rect 9171 10965 9183 10968
rect 9125 10959 9183 10965
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 9324 10996 9352 11036
rect 9398 11024 9404 11076
rect 9456 11064 9462 11076
rect 10689 11067 10747 11073
rect 10689 11064 10701 11067
rect 9456 11036 10701 11064
rect 9456 11024 9462 11036
rect 10689 11033 10701 11036
rect 10735 11033 10747 11067
rect 10689 11027 10747 11033
rect 12250 11024 12256 11076
rect 12308 11024 12314 11076
rect 13740 11036 14228 11064
rect 13740 10996 13768 11036
rect 9324 10968 13768 10996
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14090 10996 14096 11008
rect 13872 10968 14096 10996
rect 13872 10956 13878 10968
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 14200 10996 14228 11036
rect 15010 11024 15016 11076
rect 15068 11024 15074 11076
rect 15470 11024 15476 11076
rect 15528 11024 15534 11076
rect 16482 11024 16488 11076
rect 16540 11064 16546 11076
rect 17405 11067 17463 11073
rect 17405 11064 17417 11067
rect 16540 11036 17417 11064
rect 16540 11024 16546 11036
rect 17405 11033 17417 11036
rect 17451 11064 17463 11067
rect 17451 11036 17816 11064
rect 17451 11033 17463 11036
rect 17405 11027 17463 11033
rect 15378 10996 15384 11008
rect 14200 10968 15384 10996
rect 15378 10956 15384 10968
rect 15436 10956 15442 11008
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 16761 10999 16819 11005
rect 16761 10996 16773 10999
rect 16632 10968 16773 10996
rect 16632 10956 16638 10968
rect 16761 10965 16773 10968
rect 16807 10965 16819 10999
rect 17788 10996 17816 11036
rect 17862 11024 17868 11076
rect 17920 11024 17926 11076
rect 19702 11024 19708 11076
rect 19760 11064 19766 11076
rect 20257 11067 20315 11073
rect 20257 11064 20269 11067
rect 19760 11036 20269 11064
rect 19760 11024 19766 11036
rect 20257 11033 20269 11036
rect 20303 11064 20315 11067
rect 20916 11064 20944 11095
rect 20303 11036 20944 11064
rect 20303 11033 20315 11036
rect 20257 11027 20315 11033
rect 21174 11024 21180 11076
rect 21232 11024 21238 11076
rect 21818 11024 21824 11076
rect 21876 11024 21882 11076
rect 27614 11024 27620 11076
rect 27672 11064 27678 11076
rect 30009 11067 30067 11073
rect 30009 11064 30021 11067
rect 27672 11036 30021 11064
rect 27672 11024 27678 11036
rect 30009 11033 30021 11036
rect 30055 11033 30067 11067
rect 30009 11027 30067 11033
rect 31294 11024 31300 11076
rect 31352 11064 31358 11076
rect 31757 11067 31815 11073
rect 31757 11064 31769 11067
rect 31352 11036 31769 11064
rect 31352 11024 31358 11036
rect 31757 11033 31769 11036
rect 31803 11064 31815 11067
rect 47854 11064 47860 11076
rect 31803 11036 47860 11064
rect 31803 11033 31815 11036
rect 31757 11027 31815 11033
rect 47854 11024 47860 11036
rect 47912 11024 47918 11076
rect 18414 10996 18420 11008
rect 17788 10968 18420 10996
rect 16761 10959 16819 10965
rect 18414 10956 18420 10968
rect 18472 10996 18478 11008
rect 21358 10996 21364 11008
rect 18472 10968 21364 10996
rect 18472 10956 18478 10968
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 1489 10795 1547 10801
rect 1489 10761 1501 10795
rect 1535 10792 1547 10795
rect 4430 10792 4436 10804
rect 1535 10764 4436 10792
rect 1535 10761 1547 10764
rect 1489 10755 1547 10761
rect 4430 10752 4436 10764
rect 4488 10792 4494 10804
rect 4617 10795 4675 10801
rect 4617 10792 4629 10795
rect 4488 10764 4629 10792
rect 4488 10752 4494 10764
rect 4617 10761 4629 10764
rect 4663 10761 4675 10795
rect 4617 10755 4675 10761
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 5859 10764 9076 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 4798 10684 4804 10736
rect 4856 10684 4862 10736
rect 4890 10684 4896 10736
rect 4948 10724 4954 10736
rect 4948 10696 7052 10724
rect 4948 10684 4954 10696
rect 2148 10628 5304 10656
rect 2148 10597 2176 10628
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2133 10591 2191 10597
rect 2133 10588 2145 10591
rect 1903 10560 2145 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2133 10557 2145 10560
rect 2179 10557 2191 10591
rect 2133 10551 2191 10557
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10557 2467 10591
rect 2409 10551 2467 10557
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 1118 10480 1124 10532
rect 1176 10520 1182 10532
rect 2424 10520 2452 10551
rect 1176 10492 2452 10520
rect 3436 10520 3464 10551
rect 3694 10548 3700 10600
rect 3752 10548 3758 10600
rect 4246 10548 4252 10600
rect 4304 10588 4310 10600
rect 5276 10588 5304 10628
rect 5350 10616 5356 10668
rect 5408 10616 5414 10668
rect 7024 10665 7052 10696
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 8846 10616 8852 10668
rect 8904 10616 8910 10668
rect 9048 10656 9076 10764
rect 9950 10752 9956 10804
rect 10008 10752 10014 10804
rect 10781 10795 10839 10801
rect 10781 10761 10793 10795
rect 10827 10792 10839 10795
rect 11146 10792 11152 10804
rect 10827 10764 11152 10792
rect 10827 10761 10839 10764
rect 10781 10755 10839 10761
rect 11146 10752 11152 10764
rect 11204 10792 11210 10804
rect 11882 10792 11888 10804
rect 11204 10764 11888 10792
rect 11204 10752 11210 10764
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 14734 10792 14740 10804
rect 12728 10764 14740 10792
rect 9490 10684 9496 10736
rect 9548 10684 9554 10736
rect 9861 10727 9919 10733
rect 9861 10693 9873 10727
rect 9907 10724 9919 10727
rect 12728 10724 12756 10764
rect 14734 10752 14740 10764
rect 14792 10752 14798 10804
rect 14829 10795 14887 10801
rect 14829 10761 14841 10795
rect 14875 10792 14887 10795
rect 16942 10792 16948 10804
rect 14875 10764 16948 10792
rect 14875 10761 14887 10764
rect 14829 10755 14887 10761
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 17034 10752 17040 10804
rect 17092 10792 17098 10804
rect 19245 10795 19303 10801
rect 19245 10792 19257 10795
rect 17092 10764 19257 10792
rect 17092 10752 17098 10764
rect 19245 10761 19257 10764
rect 19291 10761 19303 10795
rect 21450 10792 21456 10804
rect 19245 10755 19303 10761
rect 19628 10764 21456 10792
rect 9907 10696 12756 10724
rect 9907 10693 9919 10696
rect 9861 10687 9919 10693
rect 12894 10684 12900 10736
rect 12952 10684 12958 10736
rect 15746 10684 15752 10736
rect 15804 10724 15810 10736
rect 17773 10727 17831 10733
rect 17773 10724 17785 10727
rect 15804 10696 17785 10724
rect 15804 10684 15810 10696
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 9048 10628 10701 10656
rect 10689 10625 10701 10628
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 13630 10616 13636 10668
rect 13688 10656 13694 10668
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 13688 10628 14749 10656
rect 13688 10616 13694 10628
rect 14737 10625 14749 10628
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 15933 10659 15991 10665
rect 15933 10656 15945 10659
rect 14884 10628 15945 10656
rect 14884 10616 14890 10628
rect 15933 10625 15945 10628
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 6730 10588 6736 10600
rect 4304 10560 5212 10588
rect 5276 10560 6736 10588
rect 4304 10548 4310 10560
rect 4890 10520 4896 10532
rect 3436 10492 4896 10520
rect 1176 10480 1182 10492
rect 4890 10480 4896 10492
rect 4948 10480 4954 10532
rect 5184 10529 5212 10560
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 7745 10591 7803 10597
rect 7515 10560 7604 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 5169 10523 5227 10529
rect 5169 10489 5181 10523
rect 5215 10489 5227 10523
rect 7098 10520 7104 10532
rect 5169 10483 5227 10489
rect 6472 10492 7104 10520
rect 1673 10455 1731 10461
rect 1673 10421 1685 10455
rect 1719 10452 1731 10455
rect 1946 10452 1952 10464
rect 1719 10424 1952 10452
rect 1719 10421 1731 10424
rect 1673 10415 1731 10421
rect 1946 10412 1952 10424
rect 2004 10412 2010 10464
rect 2406 10412 2412 10464
rect 2464 10452 2470 10464
rect 6472 10461 6500 10492
rect 7098 10480 7104 10492
rect 7156 10480 7162 10532
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 2464 10424 6469 10452
rect 2464 10412 2470 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6457 10415 6515 10421
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 6825 10455 6883 10461
rect 6825 10452 6837 10455
rect 6788 10424 6837 10452
rect 6788 10412 6794 10424
rect 6825 10421 6837 10424
rect 6871 10421 6883 10455
rect 7576 10452 7604 10560
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 8110 10588 8116 10600
rect 7791 10560 8116 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 8260 10560 8800 10588
rect 8260 10548 8266 10560
rect 8772 10520 8800 10560
rect 10226 10548 10232 10600
rect 10284 10588 10290 10600
rect 10962 10588 10968 10600
rect 10284 10560 10968 10588
rect 10284 10548 10290 10560
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 11296 10560 12081 10588
rect 11296 10548 11302 10560
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 12345 10591 12403 10597
rect 12345 10588 12357 10591
rect 12069 10551 12127 10557
rect 12176 10560 12357 10588
rect 10321 10523 10379 10529
rect 10321 10520 10333 10523
rect 8772 10492 10333 10520
rect 10321 10489 10333 10492
rect 10367 10489 10379 10523
rect 10321 10483 10379 10489
rect 10410 10480 10416 10532
rect 10468 10520 10474 10532
rect 11882 10520 11888 10532
rect 10468 10492 11888 10520
rect 10468 10480 10474 10492
rect 11882 10480 11888 10492
rect 11940 10480 11946 10532
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 12176 10520 12204 10560
rect 12345 10557 12357 10560
rect 12391 10557 12403 10591
rect 12345 10551 12403 10557
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15194 10588 15200 10600
rect 15059 10560 15200 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 16025 10591 16083 10597
rect 16025 10557 16037 10591
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 12032 10492 12204 10520
rect 12032 10480 12038 10492
rect 14642 10480 14648 10532
rect 14700 10520 14706 10532
rect 15565 10523 15623 10529
rect 15565 10520 15577 10523
rect 14700 10492 15577 10520
rect 14700 10480 14706 10492
rect 15565 10489 15577 10492
rect 15611 10489 15623 10523
rect 16040 10520 16068 10551
rect 16114 10548 16120 10600
rect 16172 10548 16178 10600
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 16356 10560 16865 10588
rect 16356 10548 16362 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 17420 10588 17448 10696
rect 17773 10693 17785 10696
rect 17819 10693 17831 10727
rect 17773 10687 17831 10693
rect 17862 10684 17868 10736
rect 17920 10724 17926 10736
rect 17920 10696 18262 10724
rect 17920 10684 17926 10696
rect 17494 10616 17500 10668
rect 17552 10616 17558 10668
rect 19628 10588 19656 10764
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 20254 10684 20260 10736
rect 20312 10724 20318 10736
rect 20312 10696 20470 10724
rect 20312 10684 20318 10696
rect 17420 10560 19656 10588
rect 16853 10551 16911 10557
rect 19702 10548 19708 10600
rect 19760 10548 19766 10600
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 22830 10588 22836 10600
rect 20027 10560 22836 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 22830 10548 22836 10560
rect 22888 10548 22894 10600
rect 16040 10492 16160 10520
rect 15565 10483 15623 10489
rect 7834 10452 7840 10464
rect 7576 10424 7840 10452
rect 6825 10415 6883 10421
rect 7834 10412 7840 10424
rect 7892 10452 7898 10464
rect 9858 10452 9864 10464
rect 7892 10424 9864 10452
rect 7892 10412 7898 10424
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 11514 10412 11520 10464
rect 11572 10452 11578 10464
rect 11609 10455 11667 10461
rect 11609 10452 11621 10455
rect 11572 10424 11621 10452
rect 11572 10412 11578 10424
rect 11609 10421 11621 10424
rect 11655 10421 11667 10455
rect 11609 10415 11667 10421
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 11848 10424 13829 10452
rect 11848 10412 11854 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 14369 10455 14427 10461
rect 14369 10421 14381 10455
rect 14415 10452 14427 10455
rect 15654 10452 15660 10464
rect 14415 10424 15660 10452
rect 14415 10421 14427 10424
rect 14369 10415 14427 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 16132 10452 16160 10492
rect 21358 10480 21364 10532
rect 21416 10520 21422 10532
rect 21453 10523 21511 10529
rect 21453 10520 21465 10523
rect 21416 10492 21465 10520
rect 21416 10480 21422 10492
rect 21453 10489 21465 10492
rect 21499 10489 21511 10523
rect 21453 10483 21511 10489
rect 20530 10452 20536 10464
rect 16132 10424 20536 10452
rect 20530 10412 20536 10424
rect 20588 10412 20594 10464
rect 21818 10412 21824 10464
rect 21876 10452 21882 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21876 10424 22017 10452
rect 21876 10412 21882 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 22005 10415 22063 10421
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 1210 10208 1216 10260
rect 1268 10248 1274 10260
rect 2685 10251 2743 10257
rect 2685 10248 2697 10251
rect 1268 10220 2697 10248
rect 1268 10208 1274 10220
rect 2685 10217 2697 10220
rect 2731 10217 2743 10251
rect 2685 10211 2743 10217
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 3237 10251 3295 10257
rect 3237 10248 3249 10251
rect 2924 10220 3249 10248
rect 2924 10208 2930 10220
rect 3237 10217 3249 10220
rect 3283 10217 3295 10251
rect 3237 10211 3295 10217
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 8754 10248 8760 10260
rect 7800 10220 8760 10248
rect 7800 10208 7806 10220
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 9122 10208 9128 10260
rect 9180 10208 9186 10260
rect 10045 10251 10103 10257
rect 10045 10217 10057 10251
rect 10091 10248 10103 10251
rect 10778 10248 10784 10260
rect 10091 10220 10784 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 11514 10248 11520 10260
rect 11112 10220 11520 10248
rect 11112 10208 11118 10220
rect 11514 10208 11520 10220
rect 11572 10248 11578 10260
rect 11974 10248 11980 10260
rect 11572 10220 11980 10248
rect 11572 10208 11578 10220
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 13630 10248 13636 10260
rect 12124 10220 13636 10248
rect 12124 10208 12130 10220
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 15838 10248 15844 10260
rect 13740 10220 15844 10248
rect 2961 10183 3019 10189
rect 2961 10149 2973 10183
rect 3007 10180 3019 10183
rect 3326 10180 3332 10192
rect 3007 10152 3332 10180
rect 3007 10149 3019 10152
rect 2961 10143 3019 10149
rect 3326 10140 3332 10152
rect 3384 10140 3390 10192
rect 3973 10183 4031 10189
rect 3973 10149 3985 10183
rect 4019 10180 4031 10183
rect 4154 10180 4160 10192
rect 4019 10152 4160 10180
rect 4019 10149 4031 10152
rect 3973 10143 4031 10149
rect 4154 10140 4160 10152
rect 4212 10140 4218 10192
rect 4890 10140 4896 10192
rect 4948 10180 4954 10192
rect 5902 10180 5908 10192
rect 4948 10152 5908 10180
rect 4948 10140 4954 10152
rect 5902 10140 5908 10152
rect 5960 10140 5966 10192
rect 6365 10183 6423 10189
rect 6365 10149 6377 10183
rect 6411 10180 6423 10183
rect 6549 10183 6607 10189
rect 6549 10180 6561 10183
rect 6411 10152 6561 10180
rect 6411 10149 6423 10152
rect 6365 10143 6423 10149
rect 6549 10149 6561 10152
rect 6595 10180 6607 10183
rect 6638 10180 6644 10192
rect 6595 10152 6644 10180
rect 6595 10149 6607 10152
rect 6549 10143 6607 10149
rect 6638 10140 6644 10152
rect 6696 10140 6702 10192
rect 8110 10140 8116 10192
rect 8168 10180 8174 10192
rect 8573 10183 8631 10189
rect 8573 10180 8585 10183
rect 8168 10152 8585 10180
rect 8168 10140 8174 10152
rect 8573 10149 8585 10152
rect 8619 10180 8631 10183
rect 10962 10180 10968 10192
rect 8619 10152 10968 10180
rect 8619 10149 8631 10152
rect 8573 10143 8631 10149
rect 10962 10140 10968 10152
rect 11020 10140 11026 10192
rect 13740 10180 13768 10220
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 16761 10251 16819 10257
rect 16761 10248 16773 10251
rect 16632 10220 16773 10248
rect 16632 10208 16638 10220
rect 16761 10217 16773 10220
rect 16807 10217 16819 10251
rect 16761 10211 16819 10217
rect 18874 10208 18880 10260
rect 18932 10248 18938 10260
rect 20162 10248 20168 10260
rect 18932 10220 20168 10248
rect 18932 10208 18938 10220
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 20254 10208 20260 10260
rect 20312 10248 20318 10260
rect 21453 10251 21511 10257
rect 21453 10248 21465 10251
rect 20312 10220 21465 10248
rect 20312 10208 20318 10220
rect 21453 10217 21465 10220
rect 21499 10248 21511 10251
rect 21818 10248 21824 10260
rect 21499 10220 21824 10248
rect 21499 10217 21511 10220
rect 21453 10211 21511 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 13464 10152 13768 10180
rect 1394 10072 1400 10124
rect 1452 10112 1458 10124
rect 1581 10115 1639 10121
rect 1581 10112 1593 10115
rect 1452 10084 1593 10112
rect 1452 10072 1458 10084
rect 1581 10081 1593 10084
rect 1627 10081 1639 10115
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 1581 10075 1639 10081
rect 2884 10084 4537 10112
rect 1596 9976 1624 10075
rect 2682 10004 2688 10056
rect 2740 10044 2746 10056
rect 2884 10044 2912 10084
rect 4525 10081 4537 10084
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 5813 10115 5871 10121
rect 5813 10112 5825 10115
rect 5684 10084 5825 10112
rect 5684 10072 5690 10084
rect 5813 10081 5825 10084
rect 5859 10081 5871 10115
rect 5813 10075 5871 10081
rect 6822 10072 6828 10124
rect 6880 10112 6886 10124
rect 7834 10112 7840 10124
rect 6880 10084 7840 10112
rect 6880 10072 6886 10084
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 8294 10072 8300 10124
rect 8352 10072 8358 10124
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10112 10747 10115
rect 11882 10112 11888 10124
rect 10735 10084 11888 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 11974 10072 11980 10124
rect 12032 10112 12038 10124
rect 13464 10112 13492 10152
rect 13814 10140 13820 10192
rect 13872 10180 13878 10192
rect 14093 10183 14151 10189
rect 14093 10180 14105 10183
rect 13872 10152 14105 10180
rect 13872 10140 13878 10152
rect 14093 10149 14105 10152
rect 14139 10149 14151 10183
rect 14093 10143 14151 10149
rect 12032 10084 13492 10112
rect 12032 10072 12038 10084
rect 13538 10072 13544 10124
rect 13596 10072 13602 10124
rect 14829 10115 14887 10121
rect 14829 10081 14841 10115
rect 14875 10112 14887 10115
rect 15194 10112 15200 10124
rect 14875 10084 15200 10112
rect 14875 10081 14887 10084
rect 14829 10075 14887 10081
rect 15194 10072 15200 10084
rect 15252 10112 15258 10124
rect 16206 10112 16212 10124
rect 15252 10084 16212 10112
rect 15252 10072 15258 10084
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 19429 10115 19487 10121
rect 19429 10112 19441 10115
rect 17144 10084 19441 10112
rect 2740 10016 2912 10044
rect 3145 10047 3203 10053
rect 2740 10004 2746 10016
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3418 10044 3424 10056
rect 3191 10016 3424 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10044 4307 10047
rect 4338 10044 4344 10056
rect 4295 10016 4344 10044
rect 4295 10013 4307 10016
rect 4249 10007 4307 10013
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 8312 10044 8340 10072
rect 8846 10044 8852 10056
rect 8234 10016 8852 10044
rect 8846 10004 8852 10016
rect 8904 10044 8910 10056
rect 9306 10044 9312 10056
rect 8904 10016 9312 10044
rect 8904 10004 8910 10016
rect 9306 10004 9312 10016
rect 9364 10044 9370 10056
rect 9490 10044 9496 10056
rect 9364 10016 9496 10044
rect 9364 10004 9370 10016
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10044 10563 10047
rect 11054 10044 11060 10056
rect 10551 10016 11060 10044
rect 10551 10013 10563 10016
rect 10505 10007 10563 10013
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 11238 10004 11244 10056
rect 11296 10004 11302 10056
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 14553 10047 14611 10053
rect 14553 10044 14565 10047
rect 14516 10016 14565 10044
rect 14516 10004 14522 10016
rect 14553 10013 14565 10016
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 17144 10053 17172 10084
rect 19429 10081 19441 10084
rect 19475 10112 19487 10115
rect 19702 10112 19708 10124
rect 19475 10084 19708 10112
rect 19475 10081 19487 10084
rect 19429 10075 19487 10081
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16908 10016 17141 10044
rect 16908 10004 16914 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 21818 10004 21824 10056
rect 21876 10044 21882 10056
rect 23566 10044 23572 10056
rect 21876 10016 23572 10044
rect 21876 10004 21882 10016
rect 23566 10004 23572 10016
rect 23624 10004 23630 10056
rect 4154 9976 4160 9988
rect 1596 9948 4160 9976
rect 4154 9936 4160 9948
rect 4212 9936 4218 9988
rect 6362 9976 6368 9988
rect 5368 9948 6368 9976
rect 5368 9920 5396 9948
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 7101 9979 7159 9985
rect 7101 9945 7113 9979
rect 7147 9945 7159 9979
rect 7101 9939 7159 9945
rect 9401 9979 9459 9985
rect 9401 9945 9413 9979
rect 9447 9976 9459 9979
rect 11422 9976 11428 9988
rect 9447 9948 11428 9976
rect 9447 9945 9459 9948
rect 9401 9939 9459 9945
rect 1811 9911 1869 9917
rect 1811 9877 1823 9911
rect 1857 9908 1869 9911
rect 3694 9908 3700 9920
rect 1857 9880 3700 9908
rect 1857 9877 1869 9880
rect 1811 9871 1869 9877
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 5350 9868 5356 9920
rect 5408 9868 5414 9920
rect 7116 9908 7144 9939
rect 11422 9936 11428 9948
rect 11480 9936 11486 9988
rect 11517 9979 11575 9985
rect 11517 9945 11529 9979
rect 11563 9976 11575 9979
rect 11790 9976 11796 9988
rect 11563 9948 11796 9976
rect 11563 9945 11575 9948
rect 11517 9939 11575 9945
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 11974 9976 11980 9988
rect 11900 9948 11980 9976
rect 8478 9908 8484 9920
rect 7116 9880 8484 9908
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 8570 9868 8576 9920
rect 8628 9908 8634 9920
rect 10413 9911 10471 9917
rect 10413 9908 10425 9911
rect 8628 9880 10425 9908
rect 8628 9868 8634 9880
rect 10413 9877 10425 9880
rect 10459 9877 10471 9911
rect 10413 9871 10471 9877
rect 10778 9868 10784 9920
rect 10836 9908 10842 9920
rect 11900 9908 11928 9948
rect 11974 9936 11980 9948
rect 12032 9936 12038 9988
rect 15470 9936 15476 9988
rect 15528 9936 15534 9988
rect 17034 9936 17040 9988
rect 17092 9976 17098 9988
rect 17405 9979 17463 9985
rect 17405 9976 17417 9979
rect 17092 9948 17417 9976
rect 17092 9936 17098 9948
rect 17405 9945 17417 9948
rect 17451 9945 17463 9979
rect 17862 9976 17868 9988
rect 17405 9939 17463 9945
rect 17512 9948 17868 9976
rect 10836 9880 11928 9908
rect 10836 9868 10842 9880
rect 12158 9868 12164 9920
rect 12216 9908 12222 9920
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12216 9880 13001 9908
rect 12216 9868 12222 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 15010 9868 15016 9920
rect 15068 9908 15074 9920
rect 16301 9911 16359 9917
rect 16301 9908 16313 9911
rect 15068 9880 16313 9908
rect 15068 9868 15074 9880
rect 16301 9877 16313 9880
rect 16347 9877 16359 9911
rect 16301 9871 16359 9877
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 17512 9908 17540 9948
rect 17862 9936 17868 9948
rect 17920 9936 17926 9988
rect 19242 9936 19248 9988
rect 19300 9976 19306 9988
rect 19705 9979 19763 9985
rect 19705 9976 19717 9979
rect 19300 9948 19717 9976
rect 19300 9936 19306 9948
rect 19705 9945 19717 9948
rect 19751 9945 19763 9979
rect 19705 9939 19763 9945
rect 16632 9880 17540 9908
rect 19720 9908 19748 9939
rect 20162 9936 20168 9988
rect 20220 9936 20226 9988
rect 21637 9979 21695 9985
rect 21637 9976 21649 9979
rect 21008 9948 21649 9976
rect 21008 9908 21036 9948
rect 21637 9945 21649 9948
rect 21683 9976 21695 9979
rect 23382 9976 23388 9988
rect 21683 9948 23388 9976
rect 21683 9945 21695 9948
rect 21637 9939 21695 9945
rect 23382 9936 23388 9948
rect 23440 9936 23446 9988
rect 19720 9880 21036 9908
rect 16632 9868 16638 9880
rect 21174 9868 21180 9920
rect 21232 9868 21238 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 6549 9707 6607 9713
rect 6549 9673 6561 9707
rect 6595 9704 6607 9707
rect 6638 9704 6644 9716
rect 6595 9676 6644 9704
rect 6595 9673 6607 9676
rect 6549 9667 6607 9673
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 13630 9704 13636 9716
rect 6788 9676 13636 9704
rect 6788 9664 6794 9676
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 13814 9704 13820 9716
rect 13775 9676 13820 9704
rect 13814 9664 13820 9676
rect 13872 9704 13878 9716
rect 13909 9707 13967 9713
rect 13909 9704 13921 9707
rect 13872 9676 13921 9704
rect 13872 9664 13878 9676
rect 13909 9673 13921 9676
rect 13955 9704 13967 9707
rect 13955 9676 16068 9704
rect 13955 9673 13967 9676
rect 13909 9667 13967 9673
rect 1486 9596 1492 9648
rect 1544 9596 1550 9648
rect 1673 9639 1731 9645
rect 1673 9605 1685 9639
rect 1719 9636 1731 9639
rect 1762 9636 1768 9648
rect 1719 9608 1768 9636
rect 1719 9605 1731 9608
rect 1673 9599 1731 9605
rect 1762 9596 1768 9608
rect 1820 9596 1826 9648
rect 2590 9636 2596 9648
rect 1964 9608 2596 9636
rect 1964 9577 1992 9608
rect 2590 9596 2596 9608
rect 2648 9596 2654 9648
rect 3237 9639 3295 9645
rect 3237 9605 3249 9639
rect 3283 9636 3295 9639
rect 3602 9636 3608 9648
rect 3283 9608 3608 9636
rect 3283 9605 3295 9608
rect 3237 9599 3295 9605
rect 3602 9596 3608 9608
rect 3660 9596 3666 9648
rect 5442 9596 5448 9648
rect 5500 9636 5506 9648
rect 5629 9639 5687 9645
rect 5629 9636 5641 9639
rect 5500 9608 5641 9636
rect 5500 9596 5506 9608
rect 5629 9605 5641 9608
rect 5675 9636 5687 9639
rect 5813 9639 5871 9645
rect 5813 9636 5825 9639
rect 5675 9608 5825 9636
rect 5675 9605 5687 9608
rect 5629 9599 5687 9605
rect 5813 9605 5825 9608
rect 5859 9605 5871 9639
rect 8386 9636 8392 9648
rect 5813 9599 5871 9605
rect 6564 9608 8392 9636
rect 1949 9571 2007 9577
rect 1949 9568 1961 9571
rect 1504 9540 1961 9568
rect 1504 9512 1532 9540
rect 1949 9537 1961 9540
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 2222 9528 2228 9580
rect 2280 9528 2286 9580
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3789 9571 3847 9577
rect 3789 9568 3801 9571
rect 3384 9540 3801 9568
rect 3384 9528 3390 9540
rect 3789 9537 3801 9540
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 4246 9528 4252 9580
rect 4304 9528 4310 9580
rect 1486 9460 1492 9512
rect 1544 9460 1550 9512
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 6564 9500 6592 9608
rect 8386 9596 8392 9608
rect 8444 9596 8450 9648
rect 10594 9596 10600 9648
rect 10652 9636 10658 9648
rect 10781 9639 10839 9645
rect 10781 9636 10793 9639
rect 10652 9608 10793 9636
rect 10652 9596 10658 9608
rect 10781 9605 10793 9608
rect 10827 9605 10839 9639
rect 10781 9599 10839 9605
rect 11882 9596 11888 9648
rect 11940 9636 11946 9648
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 11940 9608 11989 9636
rect 11940 9596 11946 9608
rect 11977 9605 11989 9608
rect 12023 9605 12035 9639
rect 13832 9636 13860 9664
rect 16040 9636 16068 9676
rect 16206 9664 16212 9716
rect 16264 9664 16270 9716
rect 18414 9704 18420 9716
rect 17512 9676 18420 9704
rect 16390 9636 16396 9648
rect 13202 9608 13860 9636
rect 15962 9608 16396 9636
rect 11977 9599 12035 9605
rect 16390 9596 16396 9608
rect 16448 9596 16454 9648
rect 17129 9639 17187 9645
rect 17129 9605 17141 9639
rect 17175 9636 17187 9639
rect 17512 9636 17540 9676
rect 18414 9664 18420 9676
rect 18472 9704 18478 9716
rect 18874 9704 18880 9716
rect 18472 9676 18880 9704
rect 18472 9664 18478 9676
rect 18874 9664 18880 9676
rect 18932 9664 18938 9716
rect 18506 9636 18512 9648
rect 17175 9608 17540 9636
rect 18354 9608 18512 9636
rect 17175 9605 17187 9608
rect 17129 9599 17187 9605
rect 18506 9596 18512 9608
rect 18564 9596 18570 9648
rect 19521 9639 19579 9645
rect 19521 9605 19533 9639
rect 19567 9636 19579 9639
rect 24578 9636 24584 9648
rect 19567 9608 24584 9636
rect 19567 9605 19579 9608
rect 19521 9599 19579 9605
rect 24578 9596 24584 9608
rect 24636 9596 24642 9648
rect 28629 9639 28687 9645
rect 28629 9605 28641 9639
rect 28675 9636 28687 9639
rect 31294 9636 31300 9648
rect 28675 9608 31300 9636
rect 28675 9605 28687 9608
rect 28629 9599 28687 9605
rect 6638 9528 6644 9580
rect 6696 9568 6702 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6696 9540 7113 9568
rect 6696 9528 6702 9540
rect 7101 9537 7113 9540
rect 7147 9568 7159 9571
rect 7742 9568 7748 9580
rect 7147 9540 7748 9568
rect 7147 9537 7159 9540
rect 7101 9531 7159 9537
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 9490 9528 9496 9580
rect 9548 9528 9554 9580
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 9732 9540 10701 9568
rect 9732 9528 9738 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 4571 9472 6592 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 6822 9460 6828 9512
rect 6880 9460 6886 9512
rect 7834 9460 7840 9512
rect 7892 9500 7898 9512
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 7892 9472 8125 9500
rect 7892 9460 7898 9472
rect 8113 9469 8125 9472
rect 8159 9469 8171 9503
rect 8113 9463 8171 9469
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 10226 9500 10232 9512
rect 8435 9472 10232 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 10226 9460 10232 9472
rect 10284 9460 10290 9512
rect 10962 9460 10968 9512
rect 11020 9460 11026 9512
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 11296 9472 11713 9500
rect 11296 9460 11302 9472
rect 11701 9469 11713 9472
rect 11747 9500 11759 9503
rect 14458 9500 14464 9512
rect 11747 9472 14464 9500
rect 11747 9469 11759 9472
rect 11701 9463 11759 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 14734 9460 14740 9512
rect 14792 9460 14798 9512
rect 16850 9460 16856 9512
rect 16908 9460 16914 9512
rect 17494 9460 17500 9512
rect 17552 9500 17558 9512
rect 19444 9500 19472 9531
rect 23750 9528 23756 9580
rect 23808 9568 23814 9580
rect 27525 9571 27583 9577
rect 27525 9568 27537 9571
rect 23808 9540 27537 9568
rect 23808 9528 23814 9540
rect 27525 9537 27537 9540
rect 27571 9568 27583 9571
rect 28442 9568 28448 9580
rect 27571 9540 28448 9568
rect 27571 9537 27583 9540
rect 27525 9531 27583 9537
rect 28442 9528 28448 9540
rect 28500 9528 28506 9580
rect 17552 9472 19472 9500
rect 19705 9503 19763 9509
rect 17552 9460 17558 9472
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 21174 9500 21180 9512
rect 19751 9472 21180 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 21174 9460 21180 9472
rect 21232 9460 21238 9512
rect 23382 9460 23388 9512
rect 23440 9500 23446 9512
rect 27985 9503 28043 9509
rect 27985 9500 27997 9503
rect 23440 9472 27997 9500
rect 23440 9460 23446 9472
rect 27985 9469 27997 9472
rect 28031 9469 28043 9503
rect 27985 9463 28043 9469
rect 3602 9392 3608 9444
rect 3660 9392 3666 9444
rect 6638 9432 6644 9444
rect 5368 9404 6644 9432
rect 934 9324 940 9376
rect 992 9364 998 9376
rect 5368 9364 5396 9404
rect 6638 9392 6644 9404
rect 6696 9392 6702 9444
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 10778 9432 10784 9444
rect 9548 9404 10784 9432
rect 9548 9392 9554 9404
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 13354 9392 13360 9444
rect 13412 9432 13418 9444
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 13412 9404 13461 9432
rect 13412 9392 13418 9404
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 13449 9395 13507 9401
rect 14093 9435 14151 9441
rect 14093 9401 14105 9435
rect 14139 9401 14151 9435
rect 14093 9395 14151 9401
rect 992 9336 5396 9364
rect 5537 9367 5595 9373
rect 992 9324 998 9336
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5626 9364 5632 9376
rect 5583 9336 5632 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5626 9324 5632 9336
rect 5684 9364 5690 9376
rect 5994 9364 6000 9376
rect 5684 9336 6000 9364
rect 5684 9324 5690 9336
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 8478 9324 8484 9376
rect 8536 9364 8542 9376
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 8536 9336 9873 9364
rect 8536 9324 8542 9336
rect 9861 9333 9873 9336
rect 9907 9333 9919 9367
rect 9861 9327 9919 9333
rect 10318 9324 10324 9376
rect 10376 9324 10382 9376
rect 12158 9324 12164 9376
rect 12216 9364 12222 9376
rect 12526 9364 12532 9376
rect 12216 9336 12532 9364
rect 12216 9324 12222 9336
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 13722 9364 13728 9376
rect 12768 9336 13728 9364
rect 12768 9324 12774 9336
rect 13722 9324 13728 9336
rect 13780 9364 13786 9376
rect 14108 9364 14136 9395
rect 18506 9392 18512 9444
rect 18564 9432 18570 9444
rect 18564 9404 19012 9432
rect 18564 9392 18570 9404
rect 13780 9336 14136 9364
rect 13780 9324 13786 9336
rect 14182 9324 14188 9376
rect 14240 9364 14246 9376
rect 16022 9364 16028 9376
rect 14240 9336 16028 9364
rect 14240 9324 14246 9336
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 16114 9324 16120 9376
rect 16172 9364 16178 9376
rect 18601 9367 18659 9373
rect 18601 9364 18613 9367
rect 16172 9336 18613 9364
rect 16172 9324 16178 9336
rect 18601 9333 18613 9336
rect 18647 9333 18659 9367
rect 18984 9364 19012 9404
rect 19058 9392 19064 9444
rect 19116 9392 19122 9444
rect 28644 9432 28672 9599
rect 31294 9596 31300 9608
rect 31352 9596 31358 9648
rect 27816 9404 28672 9432
rect 20073 9367 20131 9373
rect 20073 9364 20085 9367
rect 18984 9336 20085 9364
rect 18601 9327 18659 9333
rect 20073 9333 20085 9336
rect 20119 9364 20131 9367
rect 20162 9364 20168 9376
rect 20119 9336 20168 9364
rect 20119 9333 20131 9336
rect 20073 9327 20131 9333
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 27816 9373 27844 9404
rect 27801 9367 27859 9373
rect 27801 9333 27813 9367
rect 27847 9333 27859 9367
rect 27801 9327 27859 9333
rect 28442 9324 28448 9376
rect 28500 9324 28506 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 3513 9163 3571 9169
rect 3513 9160 3525 9163
rect 3476 9132 3525 9160
rect 3476 9120 3482 9132
rect 3513 9129 3525 9132
rect 3559 9129 3571 9163
rect 3513 9123 3571 9129
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 4672 9132 4752 9160
rect 4672 9120 4678 9132
rect 2869 9095 2927 9101
rect 2869 9061 2881 9095
rect 2915 9061 2927 9095
rect 2869 9055 2927 9061
rect 1578 8984 1584 9036
rect 1636 8984 1642 9036
rect 1854 8984 1860 9036
rect 1912 8984 1918 9036
rect 2884 9024 2912 9055
rect 2958 9052 2964 9104
rect 3016 9092 3022 9104
rect 3878 9092 3884 9104
rect 3016 9064 3884 9092
rect 3016 9052 3022 9064
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 4522 9024 4528 9036
rect 2884 8996 4528 9024
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 4724 9033 4752 9132
rect 4982 9120 4988 9172
rect 5040 9160 5046 9172
rect 5169 9163 5227 9169
rect 5169 9160 5181 9163
rect 5040 9132 5181 9160
rect 5040 9120 5046 9132
rect 5169 9129 5181 9132
rect 5215 9129 5227 9163
rect 5169 9123 5227 9129
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 6638 9160 6644 9172
rect 5491 9132 6644 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 7193 9163 7251 9169
rect 7193 9129 7205 9163
rect 7239 9160 7251 9163
rect 7466 9160 7472 9172
rect 7239 9132 7472 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 7837 9163 7895 9169
rect 7837 9129 7849 9163
rect 7883 9160 7895 9163
rect 9674 9160 9680 9172
rect 7883 9132 9680 9160
rect 7883 9129 7895 9132
rect 7837 9123 7895 9129
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10134 9120 10140 9172
rect 10192 9120 10198 9172
rect 11054 9120 11060 9172
rect 11112 9160 11118 9172
rect 11606 9160 11612 9172
rect 11112 9132 11612 9160
rect 11112 9120 11118 9132
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 14182 9160 14188 9172
rect 12584 9132 14188 9160
rect 12584 9120 12590 9132
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 14277 9163 14335 9169
rect 14277 9129 14289 9163
rect 14323 9160 14335 9163
rect 15930 9160 15936 9172
rect 14323 9132 15936 9160
rect 14323 9129 14335 9132
rect 14277 9123 14335 9129
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 17586 9120 17592 9172
rect 17644 9160 17650 9172
rect 17773 9163 17831 9169
rect 17773 9160 17785 9163
rect 17644 9132 17785 9160
rect 17644 9120 17650 9132
rect 17773 9129 17785 9132
rect 17819 9129 17831 9163
rect 17773 9123 17831 9129
rect 28442 9120 28448 9172
rect 28500 9160 28506 9172
rect 36354 9160 36360 9172
rect 28500 9132 36360 9160
rect 28500 9120 28506 9132
rect 36354 9120 36360 9132
rect 36412 9120 36418 9172
rect 8938 9092 8944 9104
rect 5552 9064 8944 9092
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 1596 8956 1624 8984
rect 1596 8928 2774 8956
rect 2746 8888 2774 8928
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 2924 8928 3065 8956
rect 2924 8916 2930 8928
rect 3053 8925 3065 8928
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 3326 8916 3332 8968
rect 3384 8916 3390 8968
rect 3881 8959 3939 8965
rect 3881 8925 3893 8959
rect 3927 8956 3939 8959
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3927 8928 3985 8956
rect 3927 8925 3939 8928
rect 3881 8919 3939 8925
rect 3973 8925 3985 8928
rect 4019 8956 4031 8959
rect 5552 8956 5580 9064
rect 8938 9052 8944 9064
rect 8996 9052 9002 9104
rect 15010 9092 15016 9104
rect 10796 9064 15016 9092
rect 6178 8984 6184 9036
rect 6236 8984 6242 9036
rect 6822 8984 6828 9036
rect 6880 9024 6886 9036
rect 6880 8996 8340 9024
rect 6880 8984 6886 8996
rect 4019 8928 5580 8956
rect 5905 8959 5963 8965
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 7742 8956 7748 8968
rect 7423 8928 7748 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 3418 8888 3424 8900
rect 2746 8860 3424 8888
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 5534 8848 5540 8900
rect 5592 8848 5598 8900
rect 5920 8888 5948 8919
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 8202 8916 8208 8968
rect 8260 8916 8266 8968
rect 8312 8956 8340 8996
rect 8478 8984 8484 9036
rect 8536 8984 8542 9036
rect 9398 8984 9404 9036
rect 9456 8984 9462 9036
rect 10796 9033 10824 9064
rect 15010 9052 15016 9064
rect 15068 9052 15074 9104
rect 15378 9052 15384 9104
rect 15436 9092 15442 9104
rect 15838 9092 15844 9104
rect 15436 9064 15844 9092
rect 15436 9052 15442 9064
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 10781 9027 10839 9033
rect 10781 8993 10793 9027
rect 10827 8993 10839 9027
rect 10781 8987 10839 8993
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 10928 8996 11345 9024
rect 10928 8984 10934 8996
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 11333 8987 11391 8993
rect 12250 8984 12256 9036
rect 12308 9024 12314 9036
rect 12621 9027 12679 9033
rect 12621 9024 12633 9027
rect 12308 8996 12633 9024
rect 12308 8984 12314 8996
rect 12621 8993 12633 8996
rect 12667 8993 12679 9027
rect 12621 8987 12679 8993
rect 13722 8984 13728 9036
rect 13780 9024 13786 9036
rect 14737 9027 14795 9033
rect 14737 9024 14749 9027
rect 13780 8996 14749 9024
rect 13780 8984 13786 8996
rect 14737 8993 14749 8996
rect 14783 8993 14795 9027
rect 14737 8987 14795 8993
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 9024 14979 9027
rect 15746 9024 15752 9036
rect 14967 8996 15752 9024
rect 14967 8993 14979 8996
rect 14921 8987 14979 8993
rect 15746 8984 15752 8996
rect 15804 8984 15810 9036
rect 16025 9027 16083 9033
rect 16025 8993 16037 9027
rect 16071 9024 16083 9027
rect 16850 9024 16856 9036
rect 16071 8996 16856 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 11609 8959 11667 8965
rect 8312 8928 11100 8956
rect 9122 8888 9128 8900
rect 5920 8860 9128 8888
rect 9122 8848 9128 8860
rect 9180 8848 9186 8900
rect 10505 8891 10563 8897
rect 10505 8857 10517 8891
rect 10551 8888 10563 8891
rect 10962 8888 10968 8900
rect 10551 8860 10968 8888
rect 10551 8857 10563 8860
rect 10505 8851 10563 8857
rect 10962 8848 10968 8860
rect 11020 8848 11026 8900
rect 11072 8888 11100 8928
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 11655 8928 16068 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 12802 8888 12808 8900
rect 11072 8860 12808 8888
rect 12802 8848 12808 8860
rect 12860 8848 12866 8900
rect 13541 8891 13599 8897
rect 13541 8857 13553 8891
rect 13587 8888 13599 8891
rect 14645 8891 14703 8897
rect 14645 8888 14657 8891
rect 13587 8860 14657 8888
rect 13587 8857 13599 8860
rect 13541 8851 13599 8857
rect 14645 8857 14657 8860
rect 14691 8857 14703 8891
rect 14645 8851 14703 8857
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 7006 8820 7012 8832
rect 5224 8792 7012 8820
rect 5224 8780 5230 8792
rect 7006 8780 7012 8792
rect 7064 8780 7070 8832
rect 8294 8780 8300 8832
rect 8352 8780 8358 8832
rect 9033 8823 9091 8829
rect 9033 8789 9045 8823
rect 9079 8820 9091 8823
rect 9490 8820 9496 8832
rect 9079 8792 9496 8820
rect 9079 8789 9091 8792
rect 9033 8783 9091 8789
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 9732 8792 10609 8820
rect 9732 8780 9738 8792
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 10597 8783 10655 8789
rect 10686 8780 10692 8832
rect 10744 8820 10750 8832
rect 12434 8820 12440 8832
rect 10744 8792 12440 8820
rect 10744 8780 10750 8792
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 16040 8820 16068 8928
rect 16206 8848 16212 8900
rect 16264 8888 16270 8900
rect 16301 8891 16359 8897
rect 16301 8888 16313 8891
rect 16264 8860 16313 8888
rect 16264 8848 16270 8860
rect 16301 8857 16313 8860
rect 16347 8857 16359 8891
rect 17526 8860 18184 8888
rect 16301 8851 16359 8857
rect 17218 8820 17224 8832
rect 16040 8792 17224 8820
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 18156 8829 18184 8860
rect 18141 8823 18199 8829
rect 18141 8789 18153 8823
rect 18187 8820 18199 8823
rect 18506 8820 18512 8832
rect 18187 8792 18512 8820
rect 18187 8789 18199 8792
rect 18141 8783 18199 8789
rect 18506 8780 18512 8792
rect 18564 8820 18570 8832
rect 18693 8823 18751 8829
rect 18693 8820 18705 8823
rect 18564 8792 18705 8820
rect 18564 8780 18570 8792
rect 18693 8789 18705 8792
rect 18739 8820 18751 8823
rect 18969 8823 19027 8829
rect 18969 8820 18981 8823
rect 18739 8792 18981 8820
rect 18739 8789 18751 8792
rect 18693 8783 18751 8789
rect 18969 8789 18981 8792
rect 19015 8789 19027 8823
rect 18969 8783 19027 8789
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 2924 8588 3341 8616
rect 2924 8576 2930 8588
rect 3329 8585 3341 8588
rect 3375 8585 3387 8619
rect 3329 8579 3387 8585
rect 3605 8619 3663 8625
rect 3605 8585 3617 8619
rect 3651 8616 3663 8619
rect 3694 8616 3700 8628
rect 3651 8588 3700 8616
rect 3651 8585 3663 8588
rect 3605 8579 3663 8585
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 3786 8576 3792 8628
rect 3844 8616 3850 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3844 8588 3985 8616
rect 3844 8576 3850 8588
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 3973 8579 4031 8585
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8585 4675 8619
rect 4617 8579 4675 8585
rect 3510 8508 3516 8560
rect 3568 8508 3574 8560
rect 4632 8548 4660 8579
rect 5166 8576 5172 8628
rect 5224 8576 5230 8628
rect 5813 8619 5871 8625
rect 5813 8585 5825 8619
rect 5859 8616 5871 8619
rect 5902 8616 5908 8628
rect 5859 8588 5908 8616
rect 5859 8585 5871 8588
rect 5813 8579 5871 8585
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 6362 8576 6368 8628
rect 6420 8576 6426 8628
rect 6638 8576 6644 8628
rect 6696 8576 6702 8628
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7800 8588 8033 8616
rect 7800 8576 7806 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 10042 8616 10048 8628
rect 8168 8588 10048 8616
rect 8168 8576 8174 8588
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 10137 8619 10195 8625
rect 10137 8585 10149 8619
rect 10183 8616 10195 8619
rect 10410 8616 10416 8628
rect 10183 8588 10416 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 10502 8576 10508 8628
rect 10560 8576 10566 8628
rect 11146 8576 11152 8628
rect 11204 8576 11210 8628
rect 11514 8576 11520 8628
rect 11572 8576 11578 8628
rect 12158 8576 12164 8628
rect 12216 8576 12222 8628
rect 12250 8576 12256 8628
rect 12308 8616 12314 8628
rect 12529 8619 12587 8625
rect 12529 8616 12541 8619
rect 12308 8588 12541 8616
rect 12308 8576 12314 8588
rect 12529 8585 12541 8588
rect 12575 8585 12587 8619
rect 12529 8579 12587 8585
rect 14277 8619 14335 8625
rect 14277 8585 14289 8619
rect 14323 8616 14335 8619
rect 14826 8616 14832 8628
rect 14323 8588 14832 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 14826 8576 14832 8588
rect 14884 8576 14890 8628
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 15933 8619 15991 8625
rect 15611 8588 15792 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 6914 8548 6920 8560
rect 4632 8520 6920 8548
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 7193 8551 7251 8557
rect 7193 8517 7205 8551
rect 7239 8548 7251 8551
rect 7558 8548 7564 8560
rect 7239 8520 7564 8548
rect 7239 8517 7251 8520
rect 7193 8511 7251 8517
rect 7558 8508 7564 8520
rect 7616 8548 7622 8560
rect 10686 8548 10692 8560
rect 7616 8520 10692 8548
rect 7616 8508 7622 8520
rect 10686 8508 10692 8520
rect 10744 8508 10750 8560
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 1670 8480 1676 8492
rect 1627 8452 1676 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 1670 8440 1676 8452
rect 1728 8440 1734 8492
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2130 8480 2136 8492
rect 1903 8452 2136 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3326 8480 3332 8492
rect 3099 8452 3332 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3326 8440 3332 8452
rect 3384 8480 3390 8492
rect 3528 8480 3556 8508
rect 3384 8452 3556 8480
rect 4157 8483 4215 8489
rect 3384 8440 3390 8452
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4246 8480 4252 8492
rect 4203 8452 4252 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8480 4859 8483
rect 5166 8480 5172 8492
rect 4847 8452 5172 8480
rect 4847 8449 4859 8452
rect 4801 8443 4859 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8480 7803 8483
rect 7791 8452 8616 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 1688 8412 1716 8440
rect 3510 8412 3516 8424
rect 1688 8384 3516 8412
rect 3510 8372 3516 8384
rect 3568 8372 3574 8424
rect 1026 8304 1032 8356
rect 1084 8344 1090 8356
rect 6012 8344 6040 8443
rect 7377 8415 7435 8421
rect 7377 8381 7389 8415
rect 7423 8412 7435 8415
rect 8110 8412 8116 8424
rect 7423 8384 8116 8412
rect 7423 8381 7435 8384
rect 7377 8375 7435 8381
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8381 8447 8415
rect 8588 8412 8616 8452
rect 8662 8440 8668 8492
rect 8720 8440 8726 8492
rect 11054 8480 11060 8492
rect 9416 8452 11060 8480
rect 9416 8412 9444 8452
rect 11054 8440 11060 8452
rect 11112 8440 11118 8492
rect 12618 8440 12624 8492
rect 12676 8440 12682 8492
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8480 13691 8483
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 13679 8452 14657 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 15764 8480 15792 8588
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16298 8616 16304 8628
rect 15979 8588 16304 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 17218 8576 17224 8628
rect 17276 8616 17282 8628
rect 32398 8616 32404 8628
rect 17276 8588 32404 8616
rect 17276 8576 17282 8588
rect 32398 8576 32404 8588
rect 32456 8576 32462 8628
rect 15838 8508 15844 8560
rect 15896 8548 15902 8560
rect 16025 8551 16083 8557
rect 16025 8548 16037 8551
rect 15896 8520 16037 8548
rect 15896 8508 15902 8520
rect 16025 8517 16037 8520
rect 16071 8517 16083 8551
rect 16025 8511 16083 8517
rect 16114 8508 16120 8560
rect 16172 8548 16178 8560
rect 18414 8548 18420 8560
rect 16172 8520 18420 8548
rect 16172 8508 16178 8520
rect 18414 8508 18420 8520
rect 18472 8508 18478 8560
rect 20438 8480 20444 8492
rect 15764 8452 20444 8480
rect 14645 8443 14703 8449
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 8588 8384 9444 8412
rect 8389 8375 8447 8381
rect 1084 8316 6040 8344
rect 6825 8347 6883 8353
rect 1084 8304 1090 8316
rect 6825 8313 6837 8347
rect 6871 8344 6883 8347
rect 8404 8344 8432 8375
rect 9490 8372 9496 8424
rect 9548 8412 9554 8424
rect 9677 8415 9735 8421
rect 9677 8412 9689 8415
rect 9548 8384 9689 8412
rect 9548 8372 9554 8384
rect 9677 8381 9689 8384
rect 9723 8412 9735 8415
rect 10410 8412 10416 8424
rect 9723 8384 10416 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 10594 8372 10600 8424
rect 10652 8372 10658 8424
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 12066 8412 12072 8424
rect 10827 8384 12072 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 12342 8372 12348 8424
rect 12400 8412 12406 8424
rect 12713 8415 12771 8421
rect 12713 8412 12725 8415
rect 12400 8384 12725 8412
rect 12400 8372 12406 8384
rect 12713 8381 12725 8384
rect 12759 8381 12771 8415
rect 12713 8375 12771 8381
rect 12802 8372 12808 8424
rect 12860 8412 12866 8424
rect 14737 8415 14795 8421
rect 14737 8412 14749 8415
rect 12860 8384 14749 8412
rect 12860 8372 12866 8384
rect 14737 8381 14749 8384
rect 14783 8381 14795 8415
rect 14737 8375 14795 8381
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8412 14979 8415
rect 16114 8412 16120 8424
rect 14967 8384 16120 8412
rect 14967 8381 14979 8384
rect 14921 8375 14979 8381
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8412 16267 8415
rect 20346 8412 20352 8424
rect 16255 8384 20352 8412
rect 16255 8381 16267 8384
rect 16209 8375 16267 8381
rect 20346 8372 20352 8384
rect 20404 8372 20410 8424
rect 9861 8347 9919 8353
rect 9861 8344 9873 8347
rect 6871 8316 8340 8344
rect 8404 8316 9873 8344
rect 6871 8313 6883 8316
rect 6825 8307 6883 8313
rect 2869 8279 2927 8285
rect 2869 8245 2881 8279
rect 2915 8276 2927 8279
rect 2958 8276 2964 8288
rect 2915 8248 2964 8276
rect 2915 8245 2927 8248
rect 2869 8239 2927 8245
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 7837 8279 7895 8285
rect 7837 8276 7849 8279
rect 7432 8248 7849 8276
rect 7432 8236 7438 8248
rect 7837 8245 7849 8248
rect 7883 8245 7895 8279
rect 8312 8276 8340 8316
rect 9861 8313 9873 8316
rect 9907 8344 9919 8347
rect 32858 8344 32864 8356
rect 9907 8316 32864 8344
rect 9907 8313 9919 8316
rect 9861 8307 9919 8313
rect 32858 8304 32864 8316
rect 32916 8304 32922 8356
rect 8386 8276 8392 8288
rect 8312 8248 8392 8276
rect 7837 8239 7895 8245
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 16666 8276 16672 8288
rect 12492 8248 16672 8276
rect 12492 8236 12498 8248
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 1544 8044 1593 8072
rect 1544 8032 1550 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 1581 8035 1639 8041
rect 1780 8044 2774 8072
rect 1780 7877 1808 8044
rect 2746 8004 2774 8044
rect 3326 8032 3332 8084
rect 3384 8032 3390 8084
rect 3510 8032 3516 8084
rect 3568 8032 3574 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 3970 8072 3976 8084
rect 3927 8044 3976 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 3896 8004 3924 8035
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4617 8075 4675 8081
rect 4617 8072 4629 8075
rect 4212 8044 4629 8072
rect 4212 8032 4218 8044
rect 4617 8041 4629 8044
rect 4663 8041 4675 8075
rect 4617 8035 4675 8041
rect 7558 8032 7564 8084
rect 7616 8032 7622 8084
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 8352 8044 9597 8072
rect 8352 8032 8358 8044
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 11698 8072 11704 8084
rect 9585 8035 9643 8041
rect 9692 8044 11704 8072
rect 2746 7976 3924 8004
rect 4246 7964 4252 8016
rect 4304 7964 4310 8016
rect 7190 7964 7196 8016
rect 7248 8004 7254 8016
rect 7745 8007 7803 8013
rect 7745 8004 7757 8007
rect 7248 7976 7757 8004
rect 7248 7964 7254 7976
rect 7745 7973 7757 7976
rect 7791 7973 7803 8007
rect 7745 7967 7803 7973
rect 2590 7936 2596 7948
rect 2424 7908 2596 7936
rect 2424 7877 2452 7908
rect 2590 7896 2596 7908
rect 2648 7936 2654 7948
rect 3973 7939 4031 7945
rect 3973 7936 3985 7939
rect 2648 7908 3985 7936
rect 2648 7896 2654 7908
rect 3973 7905 3985 7908
rect 4019 7905 4031 7939
rect 9692 7936 9720 8044
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12434 8032 12440 8084
rect 12492 8032 12498 8084
rect 12989 8075 13047 8081
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 17494 8072 17500 8084
rect 13035 8044 17500 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 11330 8004 11336 8016
rect 10060 7976 11336 8004
rect 10060 7945 10088 7976
rect 11330 7964 11336 7976
rect 11388 7964 11394 8016
rect 14108 7976 15148 8004
rect 3973 7899 4031 7905
rect 5552 7908 9720 7936
rect 10045 7939 10103 7945
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 2866 7828 2872 7880
rect 2924 7868 2930 7880
rect 3053 7871 3111 7877
rect 3053 7868 3065 7871
rect 2924 7840 3065 7868
rect 2924 7828 2930 7840
rect 3053 7837 3065 7840
rect 3099 7868 3111 7871
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 3099 7840 4445 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 5350 7800 5356 7812
rect 2746 7772 5356 7800
rect 2225 7735 2283 7741
rect 2225 7701 2237 7735
rect 2271 7732 2283 7735
rect 2746 7732 2774 7772
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 2271 7704 2774 7732
rect 2869 7735 2927 7741
rect 2271 7701 2283 7704
rect 2225 7695 2283 7701
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 5552 7732 5580 7908
rect 10045 7905 10057 7939
rect 10091 7905 10103 7939
rect 10045 7899 10103 7905
rect 10226 7896 10232 7948
rect 10284 7896 10290 7948
rect 14108 7945 14136 7976
rect 11517 7939 11575 7945
rect 11517 7936 11529 7939
rect 10336 7908 11529 7936
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 10336 7868 10364 7908
rect 11517 7905 11529 7908
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 14093 7939 14151 7945
rect 14093 7936 14105 7939
rect 13679 7908 14105 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 14093 7905 14105 7908
rect 14139 7905 14151 7939
rect 15120 7936 15148 7976
rect 15194 7964 15200 8016
rect 15252 7964 15258 8016
rect 19242 7936 19248 7948
rect 14093 7899 14151 7905
rect 14752 7908 15056 7936
rect 15120 7908 19248 7936
rect 5684 7840 10364 7868
rect 11241 7871 11299 7877
rect 5684 7828 5690 7840
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 7558 7760 7564 7812
rect 7616 7800 7622 7812
rect 11256 7800 11284 7831
rect 12066 7828 12072 7880
rect 12124 7868 12130 7880
rect 14752 7868 14780 7908
rect 15028 7877 15056 7908
rect 19242 7896 19248 7908
rect 19300 7896 19306 7948
rect 12124 7840 14780 7868
rect 14829 7871 14887 7877
rect 12124 7828 12130 7840
rect 14829 7837 14841 7871
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7868 15071 7871
rect 15059 7840 15884 7868
rect 15059 7837 15071 7840
rect 15013 7831 15071 7837
rect 12434 7800 12440 7812
rect 7616 7772 9674 7800
rect 11256 7772 12440 7800
rect 7616 7760 7622 7772
rect 2915 7704 5580 7732
rect 9646 7732 9674 7772
rect 12434 7760 12440 7772
rect 12492 7760 12498 7812
rect 13630 7760 13636 7812
rect 13688 7800 13694 7812
rect 14844 7800 14872 7831
rect 13688 7772 14872 7800
rect 13688 7760 13694 7772
rect 9953 7735 10011 7741
rect 9953 7732 9965 7735
rect 9646 7704 9965 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 9953 7701 9965 7704
rect 9999 7732 10011 7735
rect 12802 7732 12808 7744
rect 9999 7704 12808 7732
rect 9999 7701 10011 7704
rect 9953 7695 10011 7701
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 13354 7692 13360 7744
rect 13412 7692 13418 7744
rect 13446 7692 13452 7744
rect 13504 7692 13510 7744
rect 15856 7741 15884 7840
rect 15841 7735 15899 7741
rect 15841 7701 15853 7735
rect 15887 7732 15899 7735
rect 22830 7732 22836 7744
rect 15887 7704 22836 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 22830 7692 22836 7704
rect 22888 7732 22894 7744
rect 23382 7732 23388 7744
rect 22888 7704 23388 7732
rect 22888 7692 22894 7704
rect 23382 7692 23388 7704
rect 23440 7692 23446 7744
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 1946 7528 1952 7540
rect 1627 7500 1952 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 2222 7488 2228 7540
rect 2280 7488 2286 7540
rect 4341 7531 4399 7537
rect 4341 7528 4353 7531
rect 2332 7500 4353 7528
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 2038 7392 2044 7404
rect 1811 7364 2044 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 2038 7352 2044 7364
rect 2096 7392 2102 7404
rect 2332 7392 2360 7500
rect 4341 7497 4353 7500
rect 4387 7497 4399 7531
rect 4341 7491 4399 7497
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 11885 7531 11943 7537
rect 11885 7528 11897 7531
rect 11020 7500 11897 7528
rect 11020 7488 11026 7500
rect 11885 7497 11897 7500
rect 11931 7497 11943 7531
rect 11885 7491 11943 7497
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 13412 7500 13461 7528
rect 13412 7488 13418 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 23934 7488 23940 7540
rect 23992 7528 23998 7540
rect 27614 7528 27620 7540
rect 23992 7500 27620 7528
rect 23992 7488 23998 7500
rect 27614 7488 27620 7500
rect 27672 7488 27678 7540
rect 2958 7420 2964 7472
rect 3016 7460 3022 7472
rect 8570 7460 8576 7472
rect 3016 7432 8576 7460
rect 3016 7420 3022 7432
rect 8570 7420 8576 7432
rect 8628 7420 8634 7472
rect 9214 7420 9220 7472
rect 9272 7460 9278 7472
rect 9272 7432 12434 7460
rect 9272 7420 9278 7432
rect 2096 7364 2360 7392
rect 2409 7395 2467 7401
rect 2096 7352 2102 7364
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 2590 7392 2596 7404
rect 2455 7364 2596 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 3602 7392 3608 7404
rect 3099 7364 3608 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 3694 7352 3700 7404
rect 3752 7352 3758 7404
rect 7650 7352 7656 7404
rect 7708 7392 7714 7404
rect 9309 7395 9367 7401
rect 9309 7392 9321 7395
rect 7708 7364 9321 7392
rect 7708 7352 7714 7364
rect 9309 7361 9321 7364
rect 9355 7361 9367 7395
rect 10781 7395 10839 7401
rect 10781 7392 10793 7395
rect 9309 7355 9367 7361
rect 9416 7364 10793 7392
rect 2608 7324 2636 7352
rect 4157 7327 4215 7333
rect 4157 7324 4169 7327
rect 2608 7296 4169 7324
rect 4157 7293 4169 7296
rect 4203 7293 4215 7327
rect 4157 7287 4215 7293
rect 5258 7284 5264 7336
rect 5316 7324 5322 7336
rect 9416 7324 9444 7364
rect 10781 7361 10793 7364
rect 10827 7361 10839 7395
rect 12406 7392 12434 7432
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 12406 7364 12725 7392
rect 10781 7355 10839 7361
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 5316 7296 9444 7324
rect 5316 7284 5322 7296
rect 10318 7284 10324 7336
rect 10376 7324 10382 7336
rect 14292 7324 14320 7355
rect 22186 7352 22192 7404
rect 22244 7352 22250 7404
rect 23566 7352 23572 7404
rect 23624 7392 23630 7404
rect 24213 7395 24271 7401
rect 24213 7392 24225 7395
rect 23624 7364 24225 7392
rect 23624 7352 23630 7364
rect 24213 7361 24225 7364
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 10376 7296 14320 7324
rect 10376 7284 10382 7296
rect 22462 7284 22468 7336
rect 22520 7284 22526 7336
rect 1302 7216 1308 7268
rect 1360 7256 1366 7268
rect 3694 7256 3700 7268
rect 1360 7228 3700 7256
rect 1360 7216 1366 7228
rect 3694 7216 3700 7228
rect 3752 7256 3758 7268
rect 3973 7259 4031 7265
rect 3973 7256 3985 7259
rect 3752 7228 3985 7256
rect 3752 7216 3758 7228
rect 3973 7225 3985 7228
rect 4019 7225 4031 7259
rect 3973 7219 4031 7225
rect 10597 7259 10655 7265
rect 10597 7225 10609 7259
rect 10643 7256 10655 7259
rect 15654 7256 15660 7268
rect 10643 7228 15660 7256
rect 10643 7225 10655 7228
rect 10597 7219 10655 7225
rect 15654 7216 15660 7228
rect 15712 7216 15718 7268
rect 2869 7191 2927 7197
rect 2869 7157 2881 7191
rect 2915 7188 2927 7191
rect 2958 7188 2964 7200
rect 2915 7160 2964 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3513 7191 3571 7197
rect 3513 7157 3525 7191
rect 3559 7188 3571 7191
rect 5718 7188 5724 7200
rect 3559 7160 5724 7188
rect 3559 7157 3571 7160
rect 3513 7151 3571 7157
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 12529 7191 12587 7197
rect 12529 7157 12541 7191
rect 12575 7188 12587 7191
rect 13998 7188 14004 7200
rect 12575 7160 14004 7188
rect 12575 7157 12587 7160
rect 12529 7151 12587 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 14093 7191 14151 7197
rect 14093 7157 14105 7191
rect 14139 7188 14151 7191
rect 17494 7188 17500 7200
rect 14139 7160 17500 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 3418 6944 3424 6996
rect 3476 6944 3482 6996
rect 23201 6987 23259 6993
rect 23201 6953 23213 6987
rect 23247 6984 23259 6987
rect 23934 6984 23940 6996
rect 23247 6956 23940 6984
rect 23247 6953 23259 6956
rect 23201 6947 23259 6953
rect 23934 6944 23940 6956
rect 23992 6944 23998 6996
rect 2774 6876 2780 6928
rect 2832 6916 2838 6928
rect 2832 6888 2912 6916
rect 2832 6876 2838 6888
rect 1302 6808 1308 6860
rect 1360 6848 1366 6860
rect 2884 6848 2912 6888
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 1360 6820 2774 6848
rect 2884 6820 3801 6848
rect 1360 6808 1366 6820
rect 1762 6740 1768 6792
rect 1820 6740 1826 6792
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2590 6780 2596 6792
rect 2455 6752 2596 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 2746 6780 2774 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 3789 6811 3847 6817
rect 3970 6808 3976 6860
rect 4028 6808 4034 6860
rect 10502 6808 10508 6860
rect 10560 6848 10566 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 10560 6820 10609 6848
rect 10560 6808 10566 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 20714 6848 20720 6860
rect 19392 6820 20720 6848
rect 19392 6808 19398 6820
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 23750 6848 23756 6860
rect 22940 6820 23756 6848
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 2746 6752 3065 6780
rect 3053 6749 3065 6752
rect 3099 6780 3111 6783
rect 3513 6783 3571 6789
rect 3513 6780 3525 6783
rect 3099 6752 3525 6780
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 3513 6749 3525 6752
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 3602 6740 3608 6792
rect 3660 6780 3666 6792
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 3660 6752 4169 6780
rect 3660 6740 3666 6752
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 21726 6740 21732 6792
rect 21784 6780 21790 6792
rect 22940 6789 22968 6820
rect 23750 6808 23756 6820
rect 23808 6808 23814 6860
rect 22925 6783 22983 6789
rect 22925 6780 22937 6783
rect 21784 6752 22937 6780
rect 21784 6740 21790 6752
rect 22925 6749 22937 6752
rect 22971 6749 22983 6783
rect 22925 6743 22983 6749
rect 7282 6712 7288 6724
rect 1596 6684 7288 6712
rect 1596 6653 1624 6684
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 2225 6647 2283 6653
rect 2225 6613 2237 6647
rect 2271 6644 2283 6647
rect 2314 6644 2320 6656
rect 2271 6616 2320 6644
rect 2271 6613 2283 6616
rect 2225 6607 2283 6613
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 9766 6644 9772 6656
rect 2915 6616 9772 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 23382 6604 23388 6656
rect 23440 6604 23446 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 2869 6443 2927 6449
rect 2869 6409 2881 6443
rect 2915 6440 2927 6443
rect 4430 6440 4436 6452
rect 2915 6412 4436 6440
rect 2915 6409 2927 6412
rect 2869 6403 2927 6409
rect 4430 6400 4436 6412
rect 4488 6400 4494 6452
rect 22830 6400 22836 6452
rect 22888 6400 22894 6452
rect 1762 6332 1768 6384
rect 1820 6372 1826 6384
rect 3970 6372 3976 6384
rect 1820 6344 3976 6372
rect 1820 6332 1826 6344
rect 3970 6332 3976 6344
rect 4028 6332 4034 6384
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2924 6276 3065 6304
rect 2924 6264 2930 6276
rect 3053 6273 3065 6276
rect 3099 6304 3111 6307
rect 3329 6307 3387 6313
rect 3329 6304 3341 6307
rect 3099 6276 3341 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3329 6273 3341 6276
rect 3375 6273 3387 6307
rect 3329 6267 3387 6273
rect 22440 6307 22498 6313
rect 22440 6273 22452 6307
rect 22486 6304 22498 6307
rect 22848 6304 22876 6400
rect 22486 6276 22876 6304
rect 22486 6273 22498 6276
rect 22440 6267 22498 6273
rect 1302 6196 1308 6248
rect 1360 6236 1366 6248
rect 1581 6239 1639 6245
rect 1581 6236 1593 6239
rect 1360 6208 1593 6236
rect 1360 6196 1366 6208
rect 1581 6205 1593 6208
rect 1627 6205 1639 6239
rect 1581 6199 1639 6205
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 11422 6236 11428 6248
rect 1903 6208 11428 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 11422 6196 11428 6208
rect 11480 6196 11486 6248
rect 22511 6103 22569 6109
rect 22511 6069 22523 6103
rect 22557 6100 22569 6103
rect 22738 6100 22744 6112
rect 22557 6072 22744 6100
rect 22557 6069 22569 6072
rect 22511 6063 22569 6069
rect 22738 6060 22744 6072
rect 22796 6060 22802 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 1302 5856 1308 5908
rect 1360 5896 1366 5908
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 1360 5868 2697 5896
rect 1360 5856 1366 5868
rect 2685 5865 2697 5868
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 18877 5899 18935 5905
rect 18877 5865 18889 5899
rect 18923 5896 18935 5899
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 18923 5868 21005 5896
rect 18923 5865 18935 5868
rect 18877 5859 18935 5865
rect 20993 5865 21005 5868
rect 21039 5896 21051 5899
rect 22462 5896 22468 5908
rect 21039 5868 22468 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 7742 5788 7748 5840
rect 7800 5828 7806 5840
rect 12618 5828 12624 5840
rect 7800 5800 12624 5828
rect 7800 5788 7806 5800
rect 12618 5788 12624 5800
rect 12676 5788 12682 5840
rect 21726 5788 21732 5840
rect 21784 5788 21790 5840
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 6546 5760 6552 5772
rect 1903 5732 6552 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 13998 5720 14004 5772
rect 14056 5760 14062 5772
rect 15565 5763 15623 5769
rect 15565 5760 15577 5763
rect 14056 5732 15577 5760
rect 14056 5720 14062 5732
rect 15565 5729 15577 5732
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 17129 5763 17187 5769
rect 17129 5760 17141 5763
rect 16908 5732 17141 5760
rect 16908 5720 16914 5732
rect 17129 5729 17141 5732
rect 17175 5729 17187 5763
rect 17129 5723 17187 5729
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1360 5664 1593 5692
rect 1360 5652 1366 5664
rect 1581 5661 1593 5664
rect 1627 5692 1639 5695
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 1627 5664 2881 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 15749 5695 15807 5701
rect 15749 5692 15761 5695
rect 12676 5664 15761 5692
rect 12676 5652 12682 5664
rect 15749 5661 15761 5664
rect 15795 5692 15807 5695
rect 15795 5664 17172 5692
rect 15795 5661 15807 5664
rect 15749 5655 15807 5661
rect 16209 5559 16267 5565
rect 16209 5525 16221 5559
rect 16255 5556 16267 5559
rect 17034 5556 17040 5568
rect 16255 5528 17040 5556
rect 16255 5525 16267 5528
rect 16209 5519 16267 5525
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 17144 5556 17172 5664
rect 18506 5652 18512 5704
rect 18564 5692 18570 5704
rect 19337 5695 19395 5701
rect 19337 5692 19349 5695
rect 18564 5664 19349 5692
rect 18564 5652 18570 5664
rect 19337 5661 19349 5664
rect 19383 5661 19395 5695
rect 19337 5655 19395 5661
rect 20898 5652 20904 5704
rect 20956 5692 20962 5704
rect 21744 5692 21772 5788
rect 22738 5720 22744 5772
rect 22796 5760 22802 5772
rect 24857 5763 24915 5769
rect 24857 5760 24869 5763
rect 22796 5732 24869 5760
rect 22796 5720 22802 5732
rect 24857 5729 24869 5732
rect 24903 5729 24915 5763
rect 24857 5723 24915 5729
rect 26973 5763 27031 5769
rect 26973 5729 26985 5763
rect 27019 5760 27031 5763
rect 28718 5760 28724 5772
rect 27019 5732 28724 5760
rect 27019 5729 27031 5732
rect 26973 5723 27031 5729
rect 28718 5720 28724 5732
rect 28776 5720 28782 5772
rect 28813 5763 28871 5769
rect 28813 5729 28825 5763
rect 28859 5760 28871 5763
rect 28902 5760 28908 5772
rect 28859 5732 28908 5760
rect 28859 5729 28871 5732
rect 28813 5723 28871 5729
rect 28902 5720 28908 5732
rect 28960 5720 28966 5772
rect 20956 5664 21772 5692
rect 24673 5695 24731 5701
rect 20956 5652 20962 5664
rect 24673 5661 24685 5695
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 17402 5584 17408 5636
rect 17460 5584 17466 5636
rect 22186 5624 22192 5636
rect 18708 5596 22192 5624
rect 18708 5556 18736 5596
rect 22186 5584 22192 5596
rect 22244 5624 22250 5636
rect 23382 5624 23388 5636
rect 22244 5596 23388 5624
rect 22244 5584 22250 5596
rect 23382 5584 23388 5596
rect 23440 5584 23446 5636
rect 24688 5624 24716 5655
rect 25498 5624 25504 5636
rect 24688 5596 25504 5624
rect 25498 5584 25504 5596
rect 25556 5584 25562 5636
rect 26513 5627 26571 5633
rect 26513 5593 26525 5627
rect 26559 5593 26571 5627
rect 26513 5587 26571 5593
rect 17144 5528 18736 5556
rect 21358 5516 21364 5568
rect 21416 5516 21422 5568
rect 26528 5556 26556 5587
rect 27154 5584 27160 5636
rect 27212 5584 27218 5636
rect 27614 5556 27620 5568
rect 26528 5528 27620 5556
rect 27614 5516 27620 5528
rect 27672 5516 27678 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 22879 5355 22937 5361
rect 22879 5321 22891 5355
rect 22925 5352 22937 5355
rect 27154 5352 27160 5364
rect 22925 5324 27160 5352
rect 22925 5321 22937 5324
rect 22879 5315 22937 5321
rect 27154 5312 27160 5324
rect 27212 5312 27218 5364
rect 28534 5244 28540 5296
rect 28592 5284 28598 5296
rect 28592 5256 30052 5284
rect 28592 5244 28598 5256
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1360 5188 1593 5216
rect 1360 5176 1366 5188
rect 1581 5185 1593 5188
rect 1627 5216 1639 5219
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 1627 5188 2697 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 15654 5176 15660 5228
rect 15712 5176 15718 5228
rect 17494 5176 17500 5228
rect 17552 5176 17558 5228
rect 21358 5216 21364 5228
rect 17604 5188 21364 5216
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5148 1915 5151
rect 9030 5148 9036 5160
rect 1903 5120 9036 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 9030 5108 9036 5120
rect 9088 5108 9094 5160
rect 15470 5108 15476 5160
rect 15528 5148 15534 5160
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 15528 5120 15853 5148
rect 15528 5108 15534 5120
rect 15841 5117 15853 5120
rect 15887 5148 15899 5151
rect 17604 5148 17632 5188
rect 21358 5176 21364 5188
rect 21416 5176 21422 5228
rect 22186 5225 22192 5228
rect 22164 5219 22192 5225
rect 22164 5185 22176 5219
rect 22164 5179 22192 5185
rect 22186 5176 22192 5179
rect 22244 5176 22250 5228
rect 22776 5219 22834 5225
rect 22776 5216 22788 5219
rect 22388 5188 22788 5216
rect 15887 5120 17632 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 17678 5108 17684 5160
rect 17736 5108 17742 5160
rect 21376 5148 21404 5176
rect 22388 5148 22416 5188
rect 22776 5185 22788 5188
rect 22822 5185 22834 5219
rect 22776 5179 22834 5185
rect 21376 5120 22416 5148
rect 28629 5151 28687 5157
rect 28629 5117 28641 5151
rect 28675 5117 28687 5151
rect 28629 5111 28687 5117
rect 28644 5080 28672 5111
rect 28810 5108 28816 5160
rect 28868 5108 28874 5160
rect 30024 5157 30052 5256
rect 30009 5151 30067 5157
rect 30009 5117 30021 5151
rect 30055 5148 30067 5151
rect 41414 5148 41420 5160
rect 30055 5120 41420 5148
rect 30055 5117 30067 5120
rect 30009 5111 30067 5117
rect 41414 5108 41420 5120
rect 41472 5108 41478 5160
rect 33502 5080 33508 5092
rect 28644 5052 33508 5080
rect 33502 5040 33508 5052
rect 33560 5040 33566 5092
rect 1854 4972 1860 5024
rect 1912 5012 1918 5024
rect 2869 5015 2927 5021
rect 2869 5012 2881 5015
rect 1912 4984 2881 5012
rect 1912 4972 1918 4984
rect 2869 4981 2881 4984
rect 2915 4981 2927 5015
rect 2869 4975 2927 4981
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 17862 5012 17868 5024
rect 16347 4984 17868 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 18141 5015 18199 5021
rect 18141 4981 18153 5015
rect 18187 5012 18199 5015
rect 20530 5012 20536 5024
rect 18187 4984 20536 5012
rect 18187 4981 18199 4984
rect 18141 4975 18199 4981
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 22235 5015 22293 5021
rect 22235 4981 22247 5015
rect 22281 5012 22293 5015
rect 25958 5012 25964 5024
rect 22281 4984 25964 5012
rect 22281 4981 22293 4984
rect 22235 4975 22293 4981
rect 25958 4972 25964 4984
rect 26016 4972 26022 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 7558 4808 7564 4820
rect 2915 4780 7564 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 17402 4768 17408 4820
rect 17460 4808 17466 4820
rect 19521 4811 19579 4817
rect 19521 4808 19533 4811
rect 17460 4780 19533 4808
rect 17460 4768 17466 4780
rect 19521 4777 19533 4780
rect 19567 4777 19579 4811
rect 19521 4771 19579 4777
rect 20257 4811 20315 4817
rect 20257 4777 20269 4811
rect 20303 4808 20315 4811
rect 20898 4808 20904 4820
rect 20303 4780 20904 4808
rect 20303 4777 20315 4780
rect 20257 4771 20315 4777
rect 1302 4632 1308 4684
rect 1360 4672 1366 4684
rect 1581 4675 1639 4681
rect 1581 4672 1593 4675
rect 1360 4644 1593 4672
rect 1360 4632 1366 4644
rect 1581 4641 1593 4644
rect 1627 4641 1639 4675
rect 1581 4635 1639 4641
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 10778 4672 10784 4684
rect 1903 4644 10784 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 2866 4564 2872 4616
rect 2924 4604 2930 4616
rect 3053 4607 3111 4613
rect 3053 4604 3065 4607
rect 2924 4576 3065 4604
rect 2924 4564 2930 4576
rect 3053 4573 3065 4576
rect 3099 4604 3111 4607
rect 3329 4607 3387 4613
rect 3329 4604 3341 4607
rect 3099 4576 3341 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3329 4573 3341 4576
rect 3375 4573 3387 4607
rect 3329 4567 3387 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 20272 4604 20300 4771
rect 20898 4768 20904 4780
rect 20956 4768 20962 4820
rect 24719 4811 24777 4817
rect 24719 4777 24731 4811
rect 24765 4808 24777 4811
rect 28810 4808 28816 4820
rect 24765 4780 28816 4808
rect 24765 4777 24777 4780
rect 24719 4771 24777 4777
rect 28810 4768 28816 4780
rect 28868 4768 28874 4820
rect 25777 4675 25835 4681
rect 25777 4641 25789 4675
rect 25823 4672 25835 4675
rect 27798 4672 27804 4684
rect 25823 4644 27804 4672
rect 25823 4641 25835 4644
rect 25777 4635 25835 4641
rect 27798 4632 27804 4644
rect 27856 4632 27862 4684
rect 24616 4607 24674 4613
rect 24616 4604 24628 4607
rect 19475 4576 20300 4604
rect 22066 4576 24628 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 19889 4471 19947 4477
rect 19889 4468 19901 4471
rect 17736 4440 19901 4468
rect 17736 4428 17742 4440
rect 19889 4437 19901 4440
rect 19935 4468 19947 4471
rect 22066 4468 22094 4576
rect 24616 4573 24628 4576
rect 24662 4573 24674 4607
rect 24616 4567 24674 4573
rect 25958 4496 25964 4548
rect 26016 4496 26022 4548
rect 26418 4496 26424 4548
rect 26476 4536 26482 4548
rect 27522 4536 27528 4548
rect 26476 4508 27528 4536
rect 26476 4496 26482 4508
rect 27522 4496 27528 4508
rect 27580 4536 27586 4548
rect 27617 4539 27675 4545
rect 27617 4536 27629 4539
rect 27580 4508 27629 4536
rect 27580 4496 27586 4508
rect 27617 4505 27629 4508
rect 27663 4505 27675 4539
rect 27617 4499 27675 4505
rect 19935 4440 22094 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 1302 4224 1308 4276
rect 1360 4264 1366 4276
rect 1397 4267 1455 4273
rect 1397 4264 1409 4267
rect 1360 4236 1409 4264
rect 1360 4224 1366 4236
rect 1397 4233 1409 4236
rect 1443 4233 1455 4267
rect 1397 4227 1455 4233
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 1854 4128 1860 4140
rect 1452 4100 1860 4128
rect 1452 4088 1458 4100
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 2961 4131 3019 4137
rect 2961 4128 2973 4131
rect 2547 4100 2973 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 2961 4097 2973 4100
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 4212 4100 4261 4128
rect 4212 4088 4218 4100
rect 4249 4097 4261 4100
rect 4295 4128 4307 4131
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 4295 4100 4537 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4525 4097 4537 4100
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 4065 3995 4123 4001
rect 4065 3961 4077 3995
rect 4111 3992 4123 3995
rect 9674 3992 9680 4004
rect 4111 3964 9680 3992
rect 4111 3961 4123 3964
rect 4065 3955 4123 3961
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 3605 3927 3663 3933
rect 3605 3924 3617 3927
rect 3384 3896 3617 3924
rect 3384 3884 3390 3896
rect 3605 3893 3617 3896
rect 3651 3893 3663 3927
rect 3605 3887 3663 3893
rect 15010 3884 15016 3936
rect 15068 3884 15074 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 3973 3723 4031 3729
rect 3973 3689 3985 3723
rect 4019 3720 4031 3723
rect 10594 3720 10600 3732
rect 4019 3692 10600 3720
rect 4019 3689 4031 3692
rect 3973 3683 4031 3689
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 12066 3680 12072 3732
rect 12124 3680 12130 3732
rect 2961 3655 3019 3661
rect 2961 3621 2973 3655
rect 3007 3652 3019 3655
rect 13446 3652 13452 3664
rect 3007 3624 13452 3652
rect 3007 3621 3019 3624
rect 2961 3615 3019 3621
rect 13446 3612 13452 3624
rect 13504 3612 13510 3664
rect 28902 3612 28908 3664
rect 28960 3652 28966 3664
rect 44082 3652 44088 3664
rect 28960 3624 44088 3652
rect 28960 3612 28966 3624
rect 44082 3612 44088 3624
rect 44140 3612 44146 3664
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 1596 3556 4629 3584
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1596 3525 1624 3556
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 27522 3544 27528 3596
rect 27580 3584 27586 3596
rect 46750 3584 46756 3596
rect 27580 3556 46756 3584
rect 27580 3544 27586 3556
rect 46750 3544 46756 3556
rect 46808 3544 46814 3596
rect 1581 3519 1639 3525
rect 1581 3516 1593 3519
rect 1360 3488 1593 3516
rect 1360 3476 1366 3488
rect 1581 3485 1593 3488
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 2498 3516 2504 3528
rect 1903 3488 2504 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3145 3519 3203 3525
rect 3145 3516 3157 3519
rect 2924 3488 3157 3516
rect 2924 3476 2930 3488
rect 3145 3485 3157 3488
rect 3191 3516 3203 3519
rect 3421 3519 3479 3525
rect 3421 3516 3433 3519
rect 3191 3488 3433 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 3421 3485 3433 3488
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4157 3519 4215 3525
rect 4157 3516 4169 3519
rect 4120 3488 4169 3516
rect 4120 3476 4126 3488
rect 4157 3485 4169 3488
rect 4203 3516 4215 3519
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 4203 3488 4445 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 4433 3485 4445 3488
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 12066 3516 12072 3528
rect 11563 3488 12072 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 49418 3516 49424 3528
rect 27672 3488 49424 3516
rect 27672 3476 27678 3488
rect 49418 3476 49424 3488
rect 49476 3476 49482 3528
rect 20714 3408 20720 3460
rect 20772 3448 20778 3460
rect 38746 3448 38752 3460
rect 20772 3420 38752 3448
rect 20772 3408 20778 3420
rect 38746 3408 38752 3420
rect 38804 3408 38810 3460
rect 11606 3340 11612 3392
rect 11664 3340 11670 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 14001 3179 14059 3185
rect 14001 3176 14013 3179
rect 9824 3148 14013 3176
rect 9824 3136 9830 3148
rect 14001 3145 14013 3148
rect 14047 3145 14059 3179
rect 14001 3139 14059 3145
rect 10410 3108 10416 3120
rect 10258 3080 10416 3108
rect 10410 3068 10416 3080
rect 10468 3108 10474 3120
rect 10781 3111 10839 3117
rect 10781 3108 10793 3111
rect 10468 3080 10793 3108
rect 10468 3068 10474 3080
rect 10781 3077 10793 3080
rect 10827 3077 10839 3111
rect 10781 3071 10839 3077
rect 12618 3068 12624 3120
rect 12676 3068 12682 3120
rect 13909 3111 13967 3117
rect 13909 3077 13921 3111
rect 13955 3108 13967 3111
rect 15470 3108 15476 3120
rect 13955 3080 15476 3108
rect 13955 3077 13967 3080
rect 13909 3071 13967 3077
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 15565 3111 15623 3117
rect 15565 3077 15577 3111
rect 15611 3108 15623 3111
rect 17678 3108 17684 3120
rect 15611 3080 17684 3108
rect 15611 3077 15623 3080
rect 15565 3071 15623 3077
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 2774 3040 2780 3052
rect 1596 3012 2780 3040
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 1596 2981 1624 3012
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 3326 3040 3332 3052
rect 2915 3012 3332 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 3559 3012 4169 3040
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 1581 2975 1639 2981
rect 1581 2972 1593 2975
rect 1360 2944 1593 2972
rect 1360 2932 1366 2944
rect 1581 2941 1593 2944
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 2406 2972 2412 2984
rect 1903 2944 2412 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 6564 2972 6592 3003
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 7892 3012 8769 3040
rect 7892 3000 7898 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18325 3043 18383 3049
rect 18325 3040 18337 3043
rect 17920 3012 18337 3040
rect 17920 3000 17926 3012
rect 18325 3009 18337 3012
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 20530 3000 20536 3052
rect 20588 3000 20594 3052
rect 3988 2944 6592 2972
rect 7193 2975 7251 2981
rect 3988 2913 4016 2944
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 7239 2944 9045 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 17402 2972 17408 2984
rect 10551 2944 17408 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 3973 2907 4031 2913
rect 3973 2873 3985 2907
rect 4019 2873 4031 2907
rect 3973 2867 4031 2873
rect 10060 2876 10916 2904
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 10060 2836 10088 2876
rect 8352 2808 10088 2836
rect 10888 2836 10916 2876
rect 12434 2864 12440 2916
rect 12492 2904 12498 2916
rect 15749 2907 15807 2913
rect 15749 2904 15761 2907
rect 12492 2876 15761 2904
rect 12492 2864 12498 2876
rect 15749 2873 15761 2876
rect 15795 2873 15807 2907
rect 15749 2867 15807 2873
rect 12713 2839 12771 2845
rect 12713 2836 12725 2839
rect 10888 2808 12725 2836
rect 8352 2796 8358 2808
rect 12713 2805 12725 2808
rect 12759 2805 12771 2839
rect 12713 2799 12771 2805
rect 16853 2839 16911 2845
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 17494 2836 17500 2848
rect 16899 2808 17500 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 18141 2839 18199 2845
rect 18141 2805 18153 2839
rect 18187 2836 18199 2839
rect 20070 2836 20076 2848
rect 18187 2808 20076 2836
rect 18187 2805 18199 2808
rect 18141 2799 18199 2805
rect 20070 2796 20076 2808
rect 20128 2796 20134 2848
rect 20349 2839 20407 2845
rect 20349 2805 20361 2839
rect 20395 2836 20407 2839
rect 22002 2836 22008 2848
rect 20395 2808 22008 2836
rect 20395 2805 20407 2808
rect 20349 2799 20407 2805
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 7742 2632 7748 2644
rect 2915 2604 7748 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 25498 2592 25504 2644
rect 25556 2592 25562 2644
rect 27798 2592 27804 2644
rect 27856 2632 27862 2644
rect 28169 2635 28227 2641
rect 28169 2632 28181 2635
rect 27856 2604 28181 2632
rect 27856 2592 27862 2604
rect 28169 2601 28181 2604
rect 28215 2601 28227 2635
rect 28169 2595 28227 2601
rect 28718 2592 28724 2644
rect 28776 2632 28782 2644
rect 30837 2635 30895 2641
rect 30837 2632 30849 2635
rect 28776 2604 30849 2632
rect 28776 2592 28782 2604
rect 30837 2601 30849 2604
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 33502 2592 33508 2644
rect 33560 2592 33566 2644
rect 2774 2524 2780 2576
rect 2832 2564 2838 2576
rect 3513 2567 3571 2573
rect 3513 2564 3525 2567
rect 2832 2536 3525 2564
rect 2832 2524 2838 2536
rect 3513 2533 3525 2536
rect 3559 2533 3571 2567
rect 11606 2564 11612 2576
rect 3513 2527 3571 2533
rect 4816 2536 11612 2564
rect 1210 2456 1216 2508
rect 1268 2496 1274 2508
rect 1581 2499 1639 2505
rect 1581 2496 1593 2499
rect 1268 2468 1593 2496
rect 1268 2456 1274 2468
rect 1581 2465 1593 2468
rect 1627 2496 1639 2499
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 1627 2468 3801 2496
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 3789 2465 3801 2468
rect 3835 2465 3847 2499
rect 3789 2459 3847 2465
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4120 2468 4629 2496
rect 4120 2456 4126 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4816 2428 4844 2536
rect 11606 2524 11612 2536
rect 11664 2524 11670 2576
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6788 2468 7297 2496
rect 6788 2456 6794 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9456 2468 9965 2496
rect 9456 2456 9462 2468
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12124 2468 12633 2496
rect 12124 2456 12130 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 14734 2456 14740 2508
rect 14792 2496 14798 2508
rect 15289 2499 15347 2505
rect 15289 2496 15301 2499
rect 14792 2468 15301 2496
rect 14792 2456 14798 2468
rect 15289 2465 15301 2468
rect 15335 2465 15347 2499
rect 15289 2459 15347 2465
rect 17402 2456 17408 2508
rect 17460 2496 17466 2508
rect 17957 2499 18015 2505
rect 17957 2496 17969 2499
rect 17460 2468 17969 2496
rect 17460 2456 17466 2468
rect 17957 2465 17969 2468
rect 18003 2465 18015 2499
rect 17957 2459 18015 2465
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20220 2468 20545 2496
rect 20220 2456 20226 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22738 2456 22744 2508
rect 22796 2496 22802 2508
rect 23109 2499 23167 2505
rect 23109 2496 23121 2499
rect 22796 2468 23121 2496
rect 22796 2456 22802 2468
rect 23109 2465 23121 2468
rect 23155 2465 23167 2499
rect 23109 2459 23167 2465
rect 36354 2456 36360 2508
rect 36412 2456 36418 2508
rect 4387 2400 4844 2428
rect 7009 2431 7067 2437
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 8294 2428 8300 2440
rect 7055 2400 8300 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 3068 2360 3096 2391
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 9766 2428 9772 2440
rect 9631 2400 9772 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 12434 2428 12440 2440
rect 12391 2400 12440 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 15010 2388 15016 2440
rect 15068 2388 15074 2440
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 22002 2388 22008 2440
rect 22060 2428 22066 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22060 2400 22661 2428
rect 22060 2388 22066 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 25406 2388 25412 2440
rect 25464 2428 25470 2440
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25464 2400 25697 2428
rect 25464 2388 25470 2400
rect 25685 2397 25697 2400
rect 25731 2428 25743 2431
rect 25961 2431 26019 2437
rect 25961 2428 25973 2431
rect 25731 2400 25973 2428
rect 25731 2397 25743 2400
rect 25685 2391 25743 2397
rect 25961 2397 25973 2400
rect 26007 2397 26019 2431
rect 25961 2391 26019 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28629 2431 28687 2437
rect 28629 2428 28641 2431
rect 28408 2400 28641 2428
rect 28408 2388 28414 2400
rect 28629 2397 28641 2400
rect 28675 2397 28687 2431
rect 28629 2391 28687 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2428 31079 2431
rect 31297 2431 31355 2437
rect 31297 2428 31309 2431
rect 31067 2400 31309 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 31297 2397 31309 2400
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 33689 2431 33747 2437
rect 33689 2428 33701 2431
rect 33468 2400 33701 2428
rect 33468 2388 33474 2400
rect 33689 2397 33701 2400
rect 33735 2428 33747 2431
rect 33965 2431 34023 2437
rect 33965 2428 33977 2431
rect 33735 2400 33977 2428
rect 33735 2397 33747 2400
rect 33689 2391 33747 2397
rect 33965 2397 33977 2400
rect 34011 2397 34023 2431
rect 33965 2391 34023 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36136 2400 37289 2428
rect 36136 2388 36142 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 3329 2363 3387 2369
rect 3329 2360 3341 2363
rect 1360 2332 3341 2360
rect 1360 2320 1366 2332
rect 3329 2329 3341 2332
rect 3375 2329 3387 2363
rect 3329 2323 3387 2329
rect 1811 2295 1869 2301
rect 1811 2261 1823 2295
rect 1857 2292 1869 2295
rect 4890 2292 4896 2304
rect 1857 2264 4896 2292
rect 1857 2261 1869 2264
rect 1811 2255 1869 2261
rect 4890 2252 4896 2264
rect 4948 2252 4954 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
<< via1 >>
rect 22836 25848 22888 25900
rect 26792 25848 26844 25900
rect 25596 25780 25648 25832
rect 29184 25780 29236 25832
rect 12164 25712 12216 25764
rect 33692 25712 33744 25764
rect 10140 25644 10192 25696
rect 26884 25644 26936 25696
rect 12808 25576 12860 25628
rect 34796 25576 34848 25628
rect 10048 25508 10100 25560
rect 33600 25508 33652 25560
rect 10784 25440 10836 25492
rect 35624 25440 35676 25492
rect 15844 25372 15896 25424
rect 32864 25372 32916 25424
rect 12256 25304 12308 25356
rect 32220 25304 32272 25356
rect 13452 25236 13504 25288
rect 32588 25236 32640 25288
rect 10232 25168 10284 25220
rect 30288 25168 30340 25220
rect 15660 25100 15712 25152
rect 27620 25100 27672 25152
rect 28264 25100 28316 25152
rect 28724 25100 28776 25152
rect 3700 25032 3752 25084
rect 7564 25032 7616 25084
rect 15476 25032 15528 25084
rect 28448 25032 28500 25084
rect 15016 24964 15068 25016
rect 25596 24964 25648 25016
rect 26148 24964 26200 25016
rect 29000 24964 29052 25016
rect 14832 24896 14884 24948
rect 39304 24896 39356 24948
rect 15200 24828 15252 24880
rect 33508 24828 33560 24880
rect 25044 24760 25096 24812
rect 30472 24760 30524 24812
rect 14280 24692 14332 24744
rect 26240 24692 26292 24744
rect 27344 24692 27396 24744
rect 29552 24692 29604 24744
rect 3056 24624 3108 24676
rect 7288 24624 7340 24676
rect 14740 24624 14792 24676
rect 30012 24624 30064 24676
rect 32496 24624 32548 24676
rect 36268 24624 36320 24676
rect 3424 24556 3476 24608
rect 12256 24556 12308 24608
rect 15936 24556 15988 24608
rect 25688 24556 25740 24608
rect 27620 24556 27672 24608
rect 34152 24556 34204 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 1492 24284 1544 24336
rect 9680 24352 9732 24404
rect 3516 24216 3568 24268
rect 2412 24148 2464 24200
rect 4252 24148 4304 24200
rect 6828 24216 6880 24268
rect 9220 24216 9272 24268
rect 6644 24148 6696 24200
rect 8576 24148 8628 24200
rect 13176 24216 13228 24268
rect 10140 24148 10192 24200
rect 12440 24148 12492 24200
rect 12624 24148 12676 24200
rect 12808 24148 12860 24200
rect 14464 24284 14516 24336
rect 16212 24216 16264 24268
rect 18696 24216 18748 24268
rect 14188 24148 14240 24200
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 2780 24080 2832 24132
rect 4436 24080 4488 24132
rect 13820 24080 13872 24132
rect 3516 24012 3568 24064
rect 3700 24012 3752 24064
rect 8760 24012 8812 24064
rect 12072 24012 12124 24064
rect 12440 24012 12492 24064
rect 15384 24080 15436 24132
rect 14280 24055 14332 24064
rect 14280 24021 14289 24055
rect 14289 24021 14323 24055
rect 14323 24021 14332 24055
rect 14280 24012 14332 24021
rect 19064 24148 19116 24200
rect 19156 24148 19208 24200
rect 19800 24148 19852 24200
rect 25688 24352 25740 24404
rect 25872 24352 25924 24404
rect 29092 24352 29144 24404
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 21548 24216 21600 24268
rect 25044 24259 25096 24268
rect 25044 24225 25053 24259
rect 25053 24225 25087 24259
rect 25087 24225 25096 24259
rect 25044 24216 25096 24225
rect 24032 24191 24084 24200
rect 24032 24157 24041 24191
rect 24041 24157 24075 24191
rect 24075 24157 24084 24191
rect 24032 24148 24084 24157
rect 24952 24148 25004 24200
rect 25320 24216 25372 24268
rect 26516 24284 26568 24336
rect 27896 24284 27948 24336
rect 25872 24148 25924 24200
rect 25964 24148 26016 24200
rect 26240 24191 26292 24200
rect 26240 24157 26249 24191
rect 26249 24157 26283 24191
rect 26283 24157 26292 24191
rect 26240 24148 26292 24157
rect 26424 24148 26476 24200
rect 27804 24216 27856 24268
rect 34152 24395 34204 24404
rect 34152 24361 34161 24395
rect 34161 24361 34195 24395
rect 34195 24361 34204 24395
rect 34152 24352 34204 24361
rect 29276 24216 29328 24268
rect 30012 24259 30064 24268
rect 30012 24225 30021 24259
rect 30021 24225 30055 24259
rect 30055 24225 30064 24259
rect 30012 24216 30064 24225
rect 30380 24284 30432 24336
rect 35808 24284 35860 24336
rect 36912 24284 36964 24336
rect 38660 24327 38712 24336
rect 38660 24293 38669 24327
rect 38669 24293 38703 24327
rect 38703 24293 38712 24327
rect 38660 24284 38712 24293
rect 39304 24395 39356 24404
rect 39304 24361 39313 24395
rect 39313 24361 39347 24395
rect 39347 24361 39356 24395
rect 39304 24352 39356 24361
rect 44732 24395 44784 24404
rect 44732 24361 44741 24395
rect 44741 24361 44775 24395
rect 44775 24361 44784 24395
rect 44732 24352 44784 24361
rect 40684 24284 40736 24336
rect 39580 24216 39632 24268
rect 40132 24216 40184 24268
rect 17224 24080 17276 24132
rect 18788 24080 18840 24132
rect 25320 24080 25372 24132
rect 25504 24080 25556 24132
rect 27436 24080 27488 24132
rect 27528 24123 27580 24132
rect 27528 24089 27537 24123
rect 27537 24089 27571 24123
rect 27571 24089 27580 24123
rect 27528 24080 27580 24089
rect 27620 24080 27672 24132
rect 29000 24148 29052 24200
rect 30196 24148 30248 24200
rect 30564 24148 30616 24200
rect 31576 24148 31628 24200
rect 31852 24148 31904 24200
rect 32680 24148 32732 24200
rect 33324 24191 33376 24200
rect 33324 24157 33333 24191
rect 33333 24157 33367 24191
rect 33367 24157 33376 24191
rect 33324 24148 33376 24157
rect 34060 24191 34112 24200
rect 34060 24157 34069 24191
rect 34069 24157 34103 24191
rect 34103 24157 34112 24191
rect 34060 24148 34112 24157
rect 16948 24012 17000 24064
rect 17040 24012 17092 24064
rect 20352 24012 20404 24064
rect 24308 24012 24360 24064
rect 24952 24055 25004 24064
rect 24952 24021 24961 24055
rect 24961 24021 24995 24055
rect 24995 24021 25004 24055
rect 24952 24012 25004 24021
rect 25136 24012 25188 24064
rect 28356 24055 28408 24064
rect 28356 24021 28365 24055
rect 28365 24021 28399 24055
rect 28399 24021 28408 24055
rect 28356 24012 28408 24021
rect 34520 24080 34572 24132
rect 34980 24123 35032 24132
rect 34980 24089 34989 24123
rect 34989 24089 35023 24123
rect 35023 24089 35032 24123
rect 34980 24080 35032 24089
rect 35164 24080 35216 24132
rect 35716 24123 35768 24132
rect 35716 24089 35725 24123
rect 35725 24089 35759 24123
rect 35759 24089 35768 24123
rect 35716 24080 35768 24089
rect 35900 24148 35952 24200
rect 36820 24148 36872 24200
rect 37280 24148 37332 24200
rect 38476 24191 38528 24200
rect 38476 24157 38485 24191
rect 38485 24157 38519 24191
rect 38519 24157 38528 24191
rect 38476 24148 38528 24157
rect 39212 24191 39264 24200
rect 39212 24157 39221 24191
rect 39221 24157 39255 24191
rect 39255 24157 39264 24191
rect 39212 24148 39264 24157
rect 41512 24148 41564 24200
rect 44364 24191 44416 24200
rect 44364 24157 44373 24191
rect 44373 24157 44407 24191
rect 44407 24157 44416 24191
rect 44364 24148 44416 24157
rect 44732 24148 44784 24200
rect 45560 24148 45612 24200
rect 45928 24191 45980 24200
rect 45928 24157 45937 24191
rect 45937 24157 45971 24191
rect 45971 24157 45980 24191
rect 45928 24148 45980 24157
rect 46020 24148 46072 24200
rect 47308 24148 47360 24200
rect 48596 24191 48648 24200
rect 48596 24157 48605 24191
rect 48605 24157 48639 24191
rect 48639 24157 48648 24191
rect 48596 24148 48648 24157
rect 38292 24080 38344 24132
rect 30380 24012 30432 24064
rect 31852 24055 31904 24064
rect 31852 24021 31861 24055
rect 31861 24021 31895 24055
rect 31895 24021 31904 24055
rect 31852 24012 31904 24021
rect 32312 24055 32364 24064
rect 32312 24021 32321 24055
rect 32321 24021 32355 24055
rect 32355 24021 32364 24055
rect 32312 24012 32364 24021
rect 33416 24055 33468 24064
rect 33416 24021 33425 24055
rect 33425 24021 33459 24055
rect 33459 24021 33468 24055
rect 33416 24012 33468 24021
rect 35072 24055 35124 24064
rect 35072 24021 35081 24055
rect 35081 24021 35115 24055
rect 35115 24021 35124 24055
rect 35072 24012 35124 24021
rect 35992 24012 36044 24064
rect 36452 24012 36504 24064
rect 42064 24055 42116 24064
rect 42064 24021 42073 24055
rect 42073 24021 42107 24055
rect 42107 24021 42116 24055
rect 42064 24012 42116 24021
rect 43720 24012 43772 24064
rect 45376 24055 45428 24064
rect 45376 24021 45385 24055
rect 45385 24021 45419 24055
rect 45419 24021 45428 24055
rect 45376 24012 45428 24021
rect 46848 24055 46900 24064
rect 46848 24021 46857 24055
rect 46857 24021 46891 24055
rect 46891 24021 46900 24055
rect 46848 24012 46900 24021
rect 47124 24012 47176 24064
rect 48688 24012 48740 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 3700 23808 3752 23860
rect 5724 23808 5776 23860
rect 7104 23808 7156 23860
rect 12256 23851 12308 23860
rect 12256 23817 12265 23851
rect 12265 23817 12299 23851
rect 12299 23817 12308 23851
rect 12256 23808 12308 23817
rect 15936 23808 15988 23860
rect 4160 23740 4212 23792
rect 2136 23715 2188 23724
rect 2136 23681 2145 23715
rect 2145 23681 2179 23715
rect 2179 23681 2188 23715
rect 2136 23672 2188 23681
rect 2688 23672 2740 23724
rect 3884 23672 3936 23724
rect 8484 23740 8536 23792
rect 9956 23740 10008 23792
rect 12532 23740 12584 23792
rect 15752 23740 15804 23792
rect 4804 23715 4856 23724
rect 4804 23681 4813 23715
rect 4813 23681 4847 23715
rect 4847 23681 4856 23715
rect 4804 23672 4856 23681
rect 6552 23672 6604 23724
rect 7748 23672 7800 23724
rect 7932 23715 7984 23724
rect 7932 23681 7941 23715
rect 7941 23681 7975 23715
rect 7975 23681 7984 23715
rect 7932 23672 7984 23681
rect 11428 23672 11480 23724
rect 11520 23672 11572 23724
rect 12256 23672 12308 23724
rect 12808 23672 12860 23724
rect 13544 23672 13596 23724
rect 17132 23808 17184 23860
rect 17224 23808 17276 23860
rect 18788 23808 18840 23860
rect 18328 23740 18380 23792
rect 18880 23740 18932 23792
rect 19064 23740 19116 23792
rect 21180 23783 21232 23792
rect 21180 23749 21189 23783
rect 21189 23749 21223 23783
rect 21223 23749 21232 23783
rect 21180 23740 21232 23749
rect 21824 23740 21876 23792
rect 23296 23740 23348 23792
rect 24952 23808 25004 23860
rect 26424 23808 26476 23860
rect 25412 23740 25464 23792
rect 26516 23740 26568 23792
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 16948 23672 17000 23724
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 1216 23536 1268 23588
rect 1768 23468 1820 23520
rect 7380 23647 7432 23656
rect 7380 23613 7389 23647
rect 7389 23613 7423 23647
rect 7423 23613 7432 23647
rect 7380 23604 7432 23613
rect 17040 23604 17092 23656
rect 17868 23647 17920 23656
rect 17868 23613 17877 23647
rect 17877 23613 17911 23647
rect 17911 23613 17920 23647
rect 17868 23604 17920 23613
rect 18696 23715 18748 23724
rect 18696 23681 18705 23715
rect 18705 23681 18739 23715
rect 18739 23681 18748 23715
rect 18696 23672 18748 23681
rect 20904 23672 20956 23724
rect 29552 23808 29604 23860
rect 33600 23808 33652 23860
rect 34796 23851 34848 23860
rect 34796 23817 34805 23851
rect 34805 23817 34839 23851
rect 34839 23817 34848 23851
rect 34796 23808 34848 23817
rect 27068 23740 27120 23792
rect 27712 23740 27764 23792
rect 30104 23783 30156 23792
rect 30104 23749 30113 23783
rect 30113 23749 30147 23783
rect 30147 23749 30156 23783
rect 30104 23740 30156 23749
rect 32864 23740 32916 23792
rect 38292 23808 38344 23860
rect 38476 23851 38528 23860
rect 38476 23817 38485 23851
rect 38485 23817 38519 23851
rect 38519 23817 38528 23851
rect 38476 23808 38528 23817
rect 39212 23808 39264 23860
rect 39580 23808 39632 23860
rect 40316 23851 40368 23860
rect 40316 23817 40325 23851
rect 40325 23817 40359 23851
rect 40359 23817 40368 23851
rect 40316 23808 40368 23817
rect 40684 23851 40736 23860
rect 40684 23817 40693 23851
rect 40693 23817 40727 23851
rect 40727 23817 40736 23851
rect 40684 23808 40736 23817
rect 45928 23808 45980 23860
rect 47308 23808 47360 23860
rect 19524 23604 19576 23656
rect 13728 23536 13780 23588
rect 22376 23604 22428 23656
rect 22836 23604 22888 23656
rect 24860 23647 24912 23656
rect 24860 23613 24869 23647
rect 24869 23613 24903 23647
rect 24903 23613 24912 23647
rect 24860 23604 24912 23613
rect 25136 23604 25188 23656
rect 25780 23604 25832 23656
rect 28540 23672 28592 23724
rect 29552 23715 29604 23724
rect 29552 23681 29561 23715
rect 29561 23681 29595 23715
rect 29595 23681 29604 23715
rect 29552 23672 29604 23681
rect 30288 23715 30340 23724
rect 30288 23681 30297 23715
rect 30297 23681 30331 23715
rect 30331 23681 30340 23715
rect 30288 23672 30340 23681
rect 31392 23672 31444 23724
rect 27160 23647 27212 23656
rect 6552 23511 6604 23520
rect 6552 23477 6561 23511
rect 6561 23477 6595 23511
rect 6595 23477 6604 23511
rect 6552 23468 6604 23477
rect 9588 23468 9640 23520
rect 11520 23511 11572 23520
rect 11520 23477 11529 23511
rect 11529 23477 11563 23511
rect 11563 23477 11572 23511
rect 11520 23468 11572 23477
rect 11612 23468 11664 23520
rect 12716 23468 12768 23520
rect 13176 23468 13228 23520
rect 17776 23468 17828 23520
rect 18696 23468 18748 23520
rect 20076 23468 20128 23520
rect 20444 23511 20496 23520
rect 20444 23477 20453 23511
rect 20453 23477 20487 23511
rect 20487 23477 20496 23511
rect 20444 23468 20496 23477
rect 22284 23468 22336 23520
rect 23756 23511 23808 23520
rect 23756 23477 23765 23511
rect 23765 23477 23799 23511
rect 23799 23477 23808 23511
rect 23756 23468 23808 23477
rect 24860 23468 24912 23520
rect 27160 23613 27169 23647
rect 27169 23613 27203 23647
rect 27203 23613 27212 23647
rect 27160 23604 27212 23613
rect 26608 23511 26660 23520
rect 26608 23477 26617 23511
rect 26617 23477 26651 23511
rect 26651 23477 26660 23511
rect 26608 23468 26660 23477
rect 27252 23468 27304 23520
rect 30564 23604 30616 23656
rect 32036 23672 32088 23724
rect 31668 23604 31720 23656
rect 32220 23604 32272 23656
rect 30840 23536 30892 23588
rect 31024 23536 31076 23588
rect 34704 23715 34756 23724
rect 34704 23681 34713 23715
rect 34713 23681 34747 23715
rect 34747 23681 34756 23715
rect 34704 23672 34756 23681
rect 34520 23604 34572 23656
rect 28816 23468 28868 23520
rect 31300 23511 31352 23520
rect 31300 23477 31309 23511
rect 31309 23477 31343 23511
rect 31343 23477 31352 23511
rect 31300 23468 31352 23477
rect 31392 23468 31444 23520
rect 32220 23468 32272 23520
rect 32496 23468 32548 23520
rect 35624 23783 35676 23792
rect 35624 23749 35633 23783
rect 35633 23749 35667 23783
rect 35667 23749 35676 23783
rect 35624 23740 35676 23749
rect 35716 23740 35768 23792
rect 36268 23715 36320 23724
rect 36268 23681 36277 23715
rect 36277 23681 36311 23715
rect 36311 23681 36320 23715
rect 36268 23672 36320 23681
rect 36360 23672 36412 23724
rect 37648 23672 37700 23724
rect 44180 23740 44232 23792
rect 40960 23672 41012 23724
rect 42064 23672 42116 23724
rect 43720 23715 43772 23724
rect 43720 23681 43729 23715
rect 43729 23681 43763 23715
rect 43763 23681 43772 23715
rect 43720 23672 43772 23681
rect 43812 23672 43864 23724
rect 44640 23672 44692 23724
rect 46664 23672 46716 23724
rect 47768 23672 47820 23724
rect 48320 23672 48372 23724
rect 48688 23715 48740 23724
rect 48688 23681 48697 23715
rect 48697 23681 48731 23715
rect 48731 23681 48740 23715
rect 48688 23672 48740 23681
rect 38568 23604 38620 23656
rect 37188 23536 37240 23588
rect 41420 23536 41472 23588
rect 36084 23511 36136 23520
rect 36084 23477 36093 23511
rect 36093 23477 36127 23511
rect 36127 23477 36136 23511
rect 36084 23468 36136 23477
rect 37372 23468 37424 23520
rect 43352 23468 43404 23520
rect 45744 23511 45796 23520
rect 45744 23477 45753 23511
rect 45753 23477 45787 23511
rect 45787 23477 45796 23511
rect 45744 23468 45796 23477
rect 46940 23511 46992 23520
rect 46940 23477 46949 23511
rect 46949 23477 46983 23511
rect 46983 23477 46992 23511
rect 46940 23468 46992 23477
rect 47032 23468 47084 23520
rect 48688 23468 48740 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 1860 23264 1912 23316
rect 17868 23264 17920 23316
rect 19616 23264 19668 23316
rect 21456 23264 21508 23316
rect 22376 23264 22428 23316
rect 23296 23264 23348 23316
rect 23572 23264 23624 23316
rect 28816 23264 28868 23316
rect 29092 23264 29144 23316
rect 31300 23264 31352 23316
rect 33048 23264 33100 23316
rect 36268 23264 36320 23316
rect 36820 23307 36872 23316
rect 36820 23273 36829 23307
rect 36829 23273 36863 23307
rect 36863 23273 36872 23307
rect 36820 23264 36872 23273
rect 37280 23307 37332 23316
rect 37280 23273 37289 23307
rect 37289 23273 37323 23307
rect 37323 23273 37332 23307
rect 37280 23264 37332 23273
rect 44364 23264 44416 23316
rect 44640 23307 44692 23316
rect 44640 23273 44649 23307
rect 44649 23273 44683 23307
rect 44683 23273 44692 23307
rect 44640 23264 44692 23273
rect 48596 23264 48648 23316
rect 2872 23128 2924 23180
rect 4344 23128 4396 23180
rect 4712 23171 4764 23180
rect 4712 23137 4721 23171
rect 4721 23137 4755 23171
rect 4755 23137 4764 23171
rect 4712 23128 4764 23137
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 12900 23196 12952 23248
rect 13452 23196 13504 23248
rect 18880 23239 18932 23248
rect 18880 23205 18889 23239
rect 18889 23205 18923 23239
rect 18923 23205 18932 23239
rect 18880 23196 18932 23205
rect 19340 23196 19392 23248
rect 11428 23128 11480 23180
rect 12440 23128 12492 23180
rect 13636 23128 13688 23180
rect 17408 23128 17460 23180
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 20076 23128 20128 23137
rect 23756 23196 23808 23248
rect 21824 23171 21876 23180
rect 21824 23137 21833 23171
rect 21833 23137 21867 23171
rect 21867 23137 21876 23171
rect 21824 23128 21876 23137
rect 25136 23171 25188 23180
rect 25136 23137 25145 23171
rect 25145 23137 25179 23171
rect 25179 23137 25188 23171
rect 25136 23128 25188 23137
rect 25688 23196 25740 23248
rect 28632 23196 28684 23248
rect 28724 23196 28776 23248
rect 29736 23196 29788 23248
rect 32588 23239 32640 23248
rect 32588 23205 32597 23239
rect 32597 23205 32631 23239
rect 32631 23205 32640 23239
rect 32588 23196 32640 23205
rect 33508 23196 33560 23248
rect 33692 23196 33744 23248
rect 34888 23239 34940 23248
rect 34888 23205 34897 23239
rect 34897 23205 34931 23239
rect 34931 23205 34940 23239
rect 34888 23196 34940 23205
rect 34980 23196 35032 23248
rect 27160 23128 27212 23180
rect 27620 23128 27672 23180
rect 3424 23103 3476 23112
rect 3424 23069 3433 23103
rect 3433 23069 3467 23103
rect 3467 23069 3476 23103
rect 3424 23060 3476 23069
rect 3608 23103 3660 23112
rect 3608 23069 3617 23103
rect 3617 23069 3651 23103
rect 3651 23069 3660 23103
rect 3608 23060 3660 23069
rect 4252 23060 4304 23112
rect 7196 23103 7248 23112
rect 7196 23069 7205 23103
rect 7205 23069 7239 23103
rect 7239 23069 7248 23103
rect 7196 23060 7248 23069
rect 8944 23060 8996 23112
rect 13912 23103 13964 23112
rect 13912 23069 13921 23103
rect 13921 23069 13955 23103
rect 13955 23069 13964 23103
rect 13912 23060 13964 23069
rect 14372 23103 14424 23112
rect 14372 23069 14381 23103
rect 14381 23069 14415 23103
rect 14415 23069 14424 23103
rect 14372 23060 14424 23069
rect 15476 23103 15528 23112
rect 15476 23069 15485 23103
rect 15485 23069 15519 23103
rect 15519 23069 15528 23103
rect 15476 23060 15528 23069
rect 16856 23060 16908 23112
rect 19984 23060 20036 23112
rect 21916 23060 21968 23112
rect 25044 23060 25096 23112
rect 2780 23035 2832 23044
rect 2780 23001 2789 23035
rect 2789 23001 2823 23035
rect 2823 23001 2832 23035
rect 2780 22992 2832 23001
rect 3516 22992 3568 23044
rect 8852 22992 8904 23044
rect 4160 22967 4212 22976
rect 4160 22933 4169 22967
rect 4169 22933 4203 22967
rect 4203 22933 4212 22967
rect 4160 22924 4212 22933
rect 4528 22967 4580 22976
rect 4528 22933 4537 22967
rect 4537 22933 4571 22967
rect 4571 22933 4580 22967
rect 4528 22924 4580 22933
rect 6276 22924 6328 22976
rect 9036 22967 9088 22976
rect 9036 22933 9045 22967
rect 9045 22933 9079 22967
rect 9079 22933 9088 22967
rect 9036 22924 9088 22933
rect 9404 22924 9456 22976
rect 9588 23035 9640 23044
rect 9588 23001 9597 23035
rect 9597 23001 9631 23035
rect 9631 23001 9640 23035
rect 9588 22992 9640 23001
rect 9680 22992 9732 23044
rect 12256 22992 12308 23044
rect 17040 22992 17092 23044
rect 19064 22992 19116 23044
rect 21364 22992 21416 23044
rect 23296 22992 23348 23044
rect 11704 22924 11756 22976
rect 12624 22924 12676 22976
rect 12808 22924 12860 22976
rect 14556 22924 14608 22976
rect 15476 22924 15528 22976
rect 19340 22924 19392 22976
rect 20628 22924 20680 22976
rect 21088 22924 21140 22976
rect 23940 22924 23992 22976
rect 28540 23060 28592 23112
rect 25964 22924 26016 22976
rect 27804 22992 27856 23044
rect 28356 22924 28408 22976
rect 28908 23060 28960 23112
rect 31392 23128 31444 23180
rect 31944 23128 31996 23180
rect 36084 23128 36136 23180
rect 31484 23060 31536 23112
rect 31852 23103 31904 23112
rect 31852 23069 31861 23103
rect 31861 23069 31895 23103
rect 31895 23069 31904 23103
rect 31852 23060 31904 23069
rect 30288 22992 30340 23044
rect 32404 23035 32456 23044
rect 32404 23001 32413 23035
rect 32413 23001 32447 23035
rect 32447 23001 32456 23035
rect 32404 22992 32456 23001
rect 35072 23103 35124 23112
rect 35072 23069 35081 23103
rect 35081 23069 35115 23103
rect 35115 23069 35124 23103
rect 35072 23060 35124 23069
rect 35716 23103 35768 23112
rect 35716 23069 35725 23103
rect 35725 23069 35759 23103
rect 35759 23069 35768 23103
rect 35716 23060 35768 23069
rect 41420 23060 41472 23112
rect 43352 23103 43404 23112
rect 43352 23069 43361 23103
rect 43361 23069 43395 23103
rect 43395 23069 43404 23103
rect 43352 23060 43404 23069
rect 47860 23060 47912 23112
rect 48504 23060 48556 23112
rect 33324 22992 33376 23044
rect 33508 22992 33560 23044
rect 29828 22924 29880 22976
rect 30840 22924 30892 22976
rect 31852 22924 31904 22976
rect 32956 22924 33008 22976
rect 35532 22967 35584 22976
rect 35532 22933 35541 22967
rect 35541 22933 35575 22967
rect 35575 22933 35584 22967
rect 35532 22924 35584 22933
rect 36176 22967 36228 22976
rect 36176 22933 36185 22967
rect 36185 22933 36219 22967
rect 36219 22933 36228 22967
rect 36176 22924 36228 22933
rect 39948 22924 40000 22976
rect 47492 22924 47544 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 1032 22720 1084 22772
rect 11796 22720 11848 22772
rect 11888 22720 11940 22772
rect 12532 22720 12584 22772
rect 1952 22652 2004 22704
rect 1860 22584 1912 22636
rect 1124 22516 1176 22568
rect 4252 22584 4304 22636
rect 4804 22627 4856 22636
rect 4804 22593 4813 22627
rect 4813 22593 4847 22627
rect 4847 22593 4856 22627
rect 4804 22584 4856 22593
rect 2872 22516 2924 22568
rect 3516 22516 3568 22568
rect 2596 22380 2648 22432
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 6736 22652 6788 22704
rect 7932 22652 7984 22704
rect 10692 22695 10744 22704
rect 10692 22661 10701 22695
rect 10701 22661 10735 22695
rect 10735 22661 10744 22695
rect 10692 22652 10744 22661
rect 13636 22720 13688 22772
rect 14556 22763 14608 22772
rect 14556 22729 14565 22763
rect 14565 22729 14599 22763
rect 14599 22729 14608 22763
rect 14556 22720 14608 22729
rect 18788 22720 18840 22772
rect 19064 22720 19116 22772
rect 12808 22652 12860 22704
rect 16120 22695 16172 22704
rect 16120 22661 16129 22695
rect 16129 22661 16163 22695
rect 16163 22661 16172 22695
rect 16120 22652 16172 22661
rect 16764 22652 16816 22704
rect 6828 22584 6880 22636
rect 7840 22584 7892 22636
rect 8300 22584 8352 22636
rect 10048 22584 10100 22636
rect 11796 22627 11848 22636
rect 11796 22593 11805 22627
rect 11805 22593 11839 22627
rect 11839 22593 11848 22627
rect 11796 22584 11848 22593
rect 15016 22627 15068 22636
rect 15016 22593 15025 22627
rect 15025 22593 15059 22627
rect 15059 22593 15068 22627
rect 15016 22584 15068 22593
rect 6000 22448 6052 22500
rect 7012 22516 7064 22568
rect 8668 22559 8720 22568
rect 8668 22525 8677 22559
rect 8677 22525 8711 22559
rect 8711 22525 8720 22559
rect 8668 22516 8720 22525
rect 16856 22559 16908 22568
rect 16856 22525 16865 22559
rect 16865 22525 16899 22559
rect 16899 22525 16908 22559
rect 16856 22516 16908 22525
rect 18144 22516 18196 22568
rect 18512 22584 18564 22636
rect 19432 22584 19484 22636
rect 20076 22652 20128 22704
rect 21456 22763 21508 22772
rect 21456 22729 21465 22763
rect 21465 22729 21499 22763
rect 21499 22729 21508 22763
rect 21456 22720 21508 22729
rect 25136 22720 25188 22772
rect 25688 22763 25740 22772
rect 25688 22729 25697 22763
rect 25697 22729 25731 22763
rect 25731 22729 25740 22763
rect 25688 22720 25740 22729
rect 25780 22763 25832 22772
rect 25780 22729 25789 22763
rect 25789 22729 25823 22763
rect 25823 22729 25832 22763
rect 25780 22720 25832 22729
rect 21364 22652 21416 22704
rect 22376 22652 22428 22704
rect 23664 22652 23716 22704
rect 24400 22652 24452 22704
rect 24768 22652 24820 22704
rect 28816 22720 28868 22772
rect 27620 22652 27672 22704
rect 28632 22652 28684 22704
rect 30564 22763 30616 22772
rect 30564 22729 30573 22763
rect 30573 22729 30607 22763
rect 30607 22729 30616 22763
rect 30564 22720 30616 22729
rect 32956 22763 33008 22772
rect 32956 22729 32965 22763
rect 32965 22729 32999 22763
rect 32999 22729 33008 22763
rect 32956 22720 33008 22729
rect 33048 22720 33100 22772
rect 34704 22720 34756 22772
rect 35072 22763 35124 22772
rect 35072 22729 35081 22763
rect 35081 22729 35115 22763
rect 35115 22729 35124 22763
rect 35072 22720 35124 22729
rect 39948 22763 40000 22772
rect 39948 22729 39957 22763
rect 39957 22729 39991 22763
rect 39991 22729 40000 22763
rect 39948 22720 40000 22729
rect 47768 22763 47820 22772
rect 47768 22729 47777 22763
rect 47777 22729 47811 22763
rect 47811 22729 47820 22763
rect 47768 22720 47820 22729
rect 21916 22584 21968 22636
rect 22836 22584 22888 22636
rect 19064 22516 19116 22568
rect 20076 22516 20128 22568
rect 20444 22516 20496 22568
rect 22652 22516 22704 22568
rect 23940 22516 23992 22568
rect 25136 22516 25188 22568
rect 26608 22584 26660 22636
rect 25964 22516 26016 22568
rect 26424 22516 26476 22568
rect 27344 22584 27396 22636
rect 30932 22627 30984 22636
rect 30932 22593 30941 22627
rect 30941 22593 30975 22627
rect 30975 22593 30984 22627
rect 30932 22584 30984 22593
rect 27252 22516 27304 22568
rect 6368 22380 6420 22432
rect 7104 22380 7156 22432
rect 10048 22380 10100 22432
rect 12440 22380 12492 22432
rect 13452 22380 13504 22432
rect 18696 22380 18748 22432
rect 19248 22380 19300 22432
rect 21916 22423 21968 22432
rect 21916 22389 21925 22423
rect 21925 22389 21959 22423
rect 21959 22389 21968 22423
rect 21916 22380 21968 22389
rect 23480 22380 23532 22432
rect 23940 22380 23992 22432
rect 25320 22423 25372 22432
rect 25320 22389 25329 22423
rect 25329 22389 25363 22423
rect 25363 22389 25372 22423
rect 25320 22380 25372 22389
rect 25688 22380 25740 22432
rect 26240 22380 26292 22432
rect 26516 22380 26568 22432
rect 27436 22448 27488 22500
rect 30840 22516 30892 22568
rect 32220 22652 32272 22704
rect 31300 22584 31352 22636
rect 31208 22516 31260 22568
rect 32312 22584 32364 22636
rect 33876 22627 33928 22636
rect 33876 22593 33885 22627
rect 33885 22593 33919 22627
rect 33919 22593 33928 22627
rect 33876 22584 33928 22593
rect 34980 22627 35032 22636
rect 34980 22593 34989 22627
rect 34989 22593 35023 22627
rect 35023 22593 35032 22627
rect 34980 22584 35032 22593
rect 44732 22584 44784 22636
rect 48320 22627 48372 22636
rect 48320 22593 48329 22627
rect 48329 22593 48363 22627
rect 48363 22593 48372 22627
rect 48320 22584 48372 22593
rect 49056 22627 49108 22636
rect 49056 22593 49065 22627
rect 49065 22593 49099 22627
rect 49099 22593 49108 22627
rect 49056 22584 49108 22593
rect 31944 22448 31996 22500
rect 33600 22559 33652 22568
rect 33600 22525 33609 22559
rect 33609 22525 33643 22559
rect 33643 22525 33652 22559
rect 33600 22516 33652 22525
rect 28816 22380 28868 22432
rect 29000 22380 29052 22432
rect 32496 22423 32548 22432
rect 32496 22389 32505 22423
rect 32505 22389 32539 22423
rect 32539 22389 32548 22423
rect 32496 22380 32548 22389
rect 33416 22448 33468 22500
rect 47400 22448 47452 22500
rect 35716 22380 35768 22432
rect 37740 22380 37792 22432
rect 48504 22423 48556 22432
rect 48504 22389 48513 22423
rect 48513 22389 48547 22423
rect 48547 22389 48556 22423
rect 48504 22380 48556 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 2780 22176 2832 22228
rect 2964 22176 3016 22228
rect 4804 22176 4856 22228
rect 16120 22176 16172 22228
rect 16396 22176 16448 22228
rect 2228 22108 2280 22160
rect 3792 22108 3844 22160
rect 9496 22108 9548 22160
rect 11796 22108 11848 22160
rect 11980 22108 12032 22160
rect 14740 22108 14792 22160
rect 19892 22176 19944 22228
rect 20076 22176 20128 22228
rect 24584 22219 24636 22228
rect 24584 22185 24593 22219
rect 24593 22185 24627 22219
rect 24627 22185 24636 22219
rect 24584 22176 24636 22185
rect 22652 22108 22704 22160
rect 23204 22108 23256 22160
rect 1308 22040 1360 22092
rect 4620 22083 4672 22092
rect 4620 22049 4629 22083
rect 4629 22049 4663 22083
rect 4663 22049 4672 22083
rect 4620 22040 4672 22049
rect 1952 21972 2004 22024
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 3608 21879 3660 21888
rect 3608 21845 3617 21879
rect 3617 21845 3651 21879
rect 3651 21845 3660 21879
rect 3608 21836 3660 21845
rect 6092 21879 6144 21888
rect 6092 21845 6101 21879
rect 6101 21845 6135 21879
rect 6135 21845 6144 21879
rect 6092 21836 6144 21845
rect 6460 21972 6512 22024
rect 7380 22040 7432 22092
rect 7656 22040 7708 22092
rect 7932 22083 7984 22092
rect 7932 22049 7941 22083
rect 7941 22049 7975 22083
rect 7975 22049 7984 22083
rect 7932 22040 7984 22049
rect 8392 22040 8444 22092
rect 9036 22040 9088 22092
rect 6920 22015 6972 22024
rect 6920 21981 6929 22015
rect 6929 21981 6963 22015
rect 6963 21981 6972 22015
rect 6920 21972 6972 21981
rect 9864 22083 9916 22092
rect 9864 22049 9873 22083
rect 9873 22049 9907 22083
rect 9907 22049 9916 22083
rect 9864 22040 9916 22049
rect 10784 22040 10836 22092
rect 11244 22083 11296 22092
rect 11244 22049 11253 22083
rect 11253 22049 11287 22083
rect 11287 22049 11296 22083
rect 11244 22040 11296 22049
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 15108 22040 15160 22092
rect 19432 22040 19484 22092
rect 21916 22040 21968 22092
rect 25136 22108 25188 22160
rect 27804 22176 27856 22228
rect 28448 22176 28500 22228
rect 28908 22176 28960 22228
rect 31668 22176 31720 22228
rect 33232 22176 33284 22228
rect 27436 22108 27488 22160
rect 26792 22040 26844 22092
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 12808 21972 12860 22024
rect 15200 22015 15252 22024
rect 15200 21981 15209 22015
rect 15209 21981 15243 22015
rect 15243 21981 15252 22015
rect 15200 21972 15252 21981
rect 19524 22015 19576 22024
rect 19524 21981 19533 22015
rect 19533 21981 19567 22015
rect 19567 21981 19576 22015
rect 19524 21972 19576 21981
rect 20352 22015 20404 22024
rect 20352 21981 20361 22015
rect 20361 21981 20395 22015
rect 20395 21981 20404 22015
rect 20352 21972 20404 21981
rect 22008 21972 22060 22024
rect 22376 21972 22428 22024
rect 23664 22015 23716 22024
rect 23664 21981 23673 22015
rect 23673 21981 23707 22015
rect 23707 21981 23716 22015
rect 23664 21972 23716 21981
rect 24768 21972 24820 22024
rect 25688 21972 25740 22024
rect 29828 22040 29880 22092
rect 30748 22083 30800 22092
rect 30748 22049 30757 22083
rect 30757 22049 30791 22083
rect 30791 22049 30800 22083
rect 30748 22040 30800 22049
rect 31852 22108 31904 22160
rect 32404 22108 32456 22160
rect 8484 21836 8536 21888
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 9680 21879 9732 21888
rect 9680 21845 9689 21879
rect 9689 21845 9723 21879
rect 9723 21845 9732 21879
rect 9680 21836 9732 21845
rect 9772 21879 9824 21888
rect 9772 21845 9781 21879
rect 9781 21845 9815 21879
rect 9815 21845 9824 21879
rect 9772 21836 9824 21845
rect 12256 21836 12308 21888
rect 14096 21904 14148 21956
rect 14372 21947 14424 21956
rect 14372 21913 14381 21947
rect 14381 21913 14415 21947
rect 14415 21913 14424 21947
rect 14372 21904 14424 21913
rect 14924 21947 14976 21956
rect 14924 21913 14933 21947
rect 14933 21913 14967 21947
rect 14967 21913 14976 21947
rect 14924 21904 14976 21913
rect 17500 21904 17552 21956
rect 18144 21904 18196 21956
rect 18972 21904 19024 21956
rect 12624 21836 12676 21888
rect 16764 21836 16816 21888
rect 19340 21836 19392 21888
rect 20260 21904 20312 21956
rect 22192 21836 22244 21888
rect 22376 21879 22428 21888
rect 22376 21845 22385 21879
rect 22385 21845 22419 21879
rect 22419 21845 22428 21879
rect 22376 21836 22428 21845
rect 26332 21904 26384 21956
rect 26516 21904 26568 21956
rect 27344 21904 27396 21956
rect 25872 21836 25924 21888
rect 25964 21836 26016 21888
rect 28632 21879 28684 21888
rect 28632 21845 28641 21879
rect 28641 21845 28675 21879
rect 28675 21845 28684 21879
rect 28632 21836 28684 21845
rect 29276 21947 29328 21956
rect 29276 21913 29285 21947
rect 29285 21913 29319 21947
rect 29319 21913 29328 21947
rect 29276 21904 29328 21913
rect 30104 21879 30156 21888
rect 30104 21845 30113 21879
rect 30113 21845 30147 21879
rect 30147 21845 30156 21879
rect 30104 21836 30156 21845
rect 30472 21879 30524 21888
rect 30472 21845 30481 21879
rect 30481 21845 30515 21879
rect 30515 21845 30524 21879
rect 30472 21836 30524 21845
rect 30748 21904 30800 21956
rect 32404 21972 32456 22024
rect 32772 22040 32824 22092
rect 32864 22015 32916 22024
rect 32864 21981 32873 22015
rect 32873 21981 32907 22015
rect 32907 21981 32916 22015
rect 32864 21972 32916 21981
rect 33324 21972 33376 22024
rect 48688 21972 48740 22024
rect 49056 22015 49108 22024
rect 49056 21981 49065 22015
rect 49065 21981 49099 22015
rect 49099 21981 49108 22015
rect 49056 21972 49108 21981
rect 35808 21904 35860 21956
rect 31668 21836 31720 21888
rect 32312 21836 32364 21888
rect 44732 21836 44784 21888
rect 49240 21879 49292 21888
rect 49240 21845 49249 21879
rect 49249 21845 49283 21879
rect 49283 21845 49292 21879
rect 49240 21836 49292 21845
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 9312 21632 9364 21684
rect 2504 21496 2556 21548
rect 4344 21607 4396 21616
rect 4344 21573 4353 21607
rect 4353 21573 4387 21607
rect 4387 21573 4396 21607
rect 4344 21564 4396 21573
rect 5724 21564 5776 21616
rect 6736 21564 6788 21616
rect 7564 21564 7616 21616
rect 8024 21564 8076 21616
rect 8392 21564 8444 21616
rect 10968 21675 11020 21684
rect 10968 21641 10977 21675
rect 10977 21641 11011 21675
rect 11011 21641 11020 21675
rect 10968 21632 11020 21641
rect 16028 21675 16080 21684
rect 16028 21641 16037 21675
rect 16037 21641 16071 21675
rect 16071 21641 16080 21675
rect 16028 21632 16080 21641
rect 9588 21564 9640 21616
rect 5540 21496 5592 21548
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 7380 21496 7432 21548
rect 9496 21496 9548 21548
rect 2044 21471 2096 21480
rect 2044 21437 2053 21471
rect 2053 21437 2087 21471
rect 2087 21437 2096 21471
rect 2044 21428 2096 21437
rect 5080 21428 5132 21480
rect 6552 21428 6604 21480
rect 4896 21360 4948 21412
rect 5172 21292 5224 21344
rect 6184 21292 6236 21344
rect 8484 21428 8536 21480
rect 10324 21471 10376 21480
rect 10324 21437 10333 21471
rect 10333 21437 10367 21471
rect 10367 21437 10376 21471
rect 10324 21428 10376 21437
rect 11612 21496 11664 21548
rect 11980 21496 12032 21548
rect 10600 21428 10652 21480
rect 12256 21539 12308 21548
rect 12256 21505 12265 21539
rect 12265 21505 12299 21539
rect 12299 21505 12308 21539
rect 12256 21496 12308 21505
rect 15108 21564 15160 21616
rect 15936 21607 15988 21616
rect 15936 21573 15945 21607
rect 15945 21573 15979 21607
rect 15979 21573 15988 21607
rect 15936 21564 15988 21573
rect 12440 21496 12492 21548
rect 14648 21496 14700 21548
rect 19892 21632 19944 21684
rect 17592 21564 17644 21616
rect 18972 21564 19024 21616
rect 21364 21632 21416 21684
rect 22836 21632 22888 21684
rect 13360 21471 13412 21480
rect 13360 21437 13369 21471
rect 13369 21437 13403 21471
rect 13403 21437 13412 21471
rect 13360 21428 13412 21437
rect 14096 21428 14148 21480
rect 8944 21292 8996 21344
rect 9588 21292 9640 21344
rect 11060 21292 11112 21344
rect 11520 21292 11572 21344
rect 11796 21335 11848 21344
rect 11796 21301 11805 21335
rect 11805 21301 11839 21335
rect 11839 21301 11848 21335
rect 11796 21292 11848 21301
rect 15568 21403 15620 21412
rect 15568 21369 15577 21403
rect 15577 21369 15611 21403
rect 15611 21369 15620 21403
rect 15568 21360 15620 21369
rect 17316 21471 17368 21480
rect 17316 21437 17325 21471
rect 17325 21437 17359 21471
rect 17359 21437 17368 21471
rect 17316 21428 17368 21437
rect 17224 21360 17276 21412
rect 13544 21292 13596 21344
rect 14740 21292 14792 21344
rect 14924 21292 14976 21344
rect 18604 21292 18656 21344
rect 18972 21471 19024 21480
rect 18972 21437 18981 21471
rect 18981 21437 19015 21471
rect 19015 21437 19024 21471
rect 18972 21428 19024 21437
rect 19064 21428 19116 21480
rect 22928 21564 22980 21616
rect 25044 21632 25096 21684
rect 23940 21564 23992 21616
rect 24400 21564 24452 21616
rect 23388 21539 23440 21548
rect 23388 21505 23397 21539
rect 23397 21505 23431 21539
rect 23431 21505 23440 21539
rect 23388 21496 23440 21505
rect 25964 21675 26016 21684
rect 25964 21641 25973 21675
rect 25973 21641 26007 21675
rect 26007 21641 26016 21675
rect 25964 21632 26016 21641
rect 26332 21632 26384 21684
rect 20260 21360 20312 21412
rect 19432 21292 19484 21344
rect 19708 21292 19760 21344
rect 24676 21428 24728 21480
rect 26608 21428 26660 21480
rect 26884 21496 26936 21548
rect 27344 21496 27396 21548
rect 27896 21496 27948 21548
rect 24768 21360 24820 21412
rect 27620 21360 27672 21412
rect 28724 21564 28776 21616
rect 29000 21564 29052 21616
rect 33232 21675 33284 21684
rect 33232 21641 33241 21675
rect 33241 21641 33275 21675
rect 33275 21641 33284 21675
rect 33232 21632 33284 21641
rect 29828 21496 29880 21548
rect 28448 21471 28500 21480
rect 28448 21437 28457 21471
rect 28457 21437 28491 21471
rect 28491 21437 28500 21471
rect 28448 21428 28500 21437
rect 28724 21471 28776 21480
rect 28724 21437 28733 21471
rect 28733 21437 28767 21471
rect 28767 21437 28776 21471
rect 28724 21428 28776 21437
rect 28816 21428 28868 21480
rect 25320 21292 25372 21344
rect 30104 21292 30156 21344
rect 30196 21335 30248 21344
rect 30196 21301 30205 21335
rect 30205 21301 30239 21335
rect 30239 21301 30248 21335
rect 30196 21292 30248 21301
rect 30656 21335 30708 21344
rect 30656 21301 30665 21335
rect 30665 21301 30699 21335
rect 30699 21301 30708 21335
rect 30656 21292 30708 21301
rect 31484 21496 31536 21548
rect 32220 21496 32272 21548
rect 34520 21564 34572 21616
rect 35532 21496 35584 21548
rect 47860 21496 47912 21548
rect 31576 21428 31628 21480
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 31392 21360 31444 21412
rect 32404 21360 32456 21412
rect 31760 21292 31812 21344
rect 32496 21335 32548 21344
rect 32496 21301 32505 21335
rect 32505 21301 32539 21335
rect 32539 21301 32548 21335
rect 32496 21292 32548 21301
rect 33416 21335 33468 21344
rect 33416 21301 33425 21335
rect 33425 21301 33459 21335
rect 33459 21301 33468 21335
rect 33416 21292 33468 21301
rect 47860 21292 47912 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 7104 21088 7156 21140
rect 3332 21020 3384 21072
rect 6736 21020 6788 21072
rect 10324 21088 10376 21140
rect 15200 21088 15252 21140
rect 7656 21020 7708 21072
rect 2136 20952 2188 21004
rect 4160 20952 4212 21004
rect 4252 20995 4304 21004
rect 4252 20961 4261 20995
rect 4261 20961 4295 20995
rect 4295 20961 4304 20995
rect 4252 20952 4304 20961
rect 7012 20952 7064 21004
rect 7380 20952 7432 21004
rect 11796 21020 11848 21072
rect 8852 20952 8904 21004
rect 1860 20884 1912 20936
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 5448 20927 5500 20936
rect 5448 20893 5457 20927
rect 5457 20893 5491 20927
rect 5491 20893 5500 20927
rect 5448 20884 5500 20893
rect 8208 20927 8260 20936
rect 8208 20893 8217 20927
rect 8217 20893 8251 20927
rect 8251 20893 8260 20927
rect 8208 20884 8260 20893
rect 8576 20884 8628 20936
rect 11520 20952 11572 21004
rect 14648 21020 14700 21072
rect 12532 20995 12584 21004
rect 12532 20961 12541 20995
rect 12541 20961 12575 20995
rect 12575 20961 12584 20995
rect 12532 20952 12584 20961
rect 14924 20952 14976 21004
rect 15476 20952 15528 21004
rect 23572 21088 23624 21140
rect 23664 21088 23716 21140
rect 16396 20995 16448 21004
rect 16396 20961 16405 20995
rect 16405 20961 16439 20995
rect 16439 20961 16448 20995
rect 16396 20952 16448 20961
rect 21364 21020 21416 21072
rect 22376 21020 22428 21072
rect 19708 20995 19760 21004
rect 9036 20884 9088 20936
rect 11704 20884 11756 20936
rect 12072 20884 12124 20936
rect 2780 20859 2832 20868
rect 2780 20825 2789 20859
rect 2789 20825 2823 20859
rect 2823 20825 2832 20859
rect 2780 20816 2832 20825
rect 3516 20816 3568 20868
rect 5632 20816 5684 20868
rect 5264 20748 5316 20800
rect 6184 20816 6236 20868
rect 7104 20816 7156 20868
rect 10600 20816 10652 20868
rect 11336 20859 11388 20868
rect 11336 20825 11345 20859
rect 11345 20825 11379 20859
rect 11379 20825 11388 20859
rect 11336 20816 11388 20825
rect 14096 20816 14148 20868
rect 16580 20884 16632 20936
rect 17408 20927 17460 20936
rect 17408 20893 17417 20927
rect 17417 20893 17451 20927
rect 17451 20893 17460 20927
rect 17408 20884 17460 20893
rect 18604 20884 18656 20936
rect 19708 20961 19717 20995
rect 19717 20961 19751 20995
rect 19751 20961 19760 20995
rect 19708 20952 19760 20961
rect 21456 20952 21508 21004
rect 23572 20952 23624 21004
rect 23848 20995 23900 21004
rect 23848 20961 23857 20995
rect 23857 20961 23891 20995
rect 23891 20961 23900 20995
rect 23848 20952 23900 20961
rect 18880 20884 18932 20936
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 22284 20884 22336 20936
rect 24124 20884 24176 20936
rect 24768 20884 24820 20936
rect 27712 21088 27764 21140
rect 27804 21131 27856 21140
rect 27804 21097 27813 21131
rect 27813 21097 27847 21131
rect 27847 21097 27856 21131
rect 27804 21088 27856 21097
rect 27896 21088 27948 21140
rect 28908 21088 28960 21140
rect 30012 21088 30064 21140
rect 30104 21088 30156 21140
rect 31392 21088 31444 21140
rect 32588 21088 32640 21140
rect 44824 21088 44876 21140
rect 47492 21088 47544 21140
rect 49056 21088 49108 21140
rect 28264 21020 28316 21072
rect 25688 20995 25740 21004
rect 25688 20961 25697 20995
rect 25697 20961 25731 20995
rect 25731 20961 25740 20995
rect 26056 20995 26108 21004
rect 25688 20952 25740 20961
rect 26056 20961 26065 20995
rect 26065 20961 26099 20995
rect 26099 20961 26108 20995
rect 26056 20952 26108 20961
rect 27620 20952 27672 21004
rect 33416 21020 33468 21072
rect 29092 20952 29144 21004
rect 30472 20952 30524 21004
rect 31668 20952 31720 21004
rect 36452 20952 36504 21004
rect 25872 20884 25924 20936
rect 28448 20884 28500 20936
rect 29276 20884 29328 20936
rect 29552 20884 29604 20936
rect 31116 20927 31168 20936
rect 31116 20893 31125 20927
rect 31125 20893 31159 20927
rect 31159 20893 31168 20927
rect 31116 20884 31168 20893
rect 32680 20927 32732 20936
rect 32680 20893 32689 20927
rect 32689 20893 32723 20927
rect 32723 20893 32732 20927
rect 32680 20884 32732 20893
rect 5908 20748 5960 20800
rect 9220 20748 9272 20800
rect 11428 20791 11480 20800
rect 11428 20757 11437 20791
rect 11437 20757 11471 20791
rect 11471 20757 11480 20791
rect 11428 20748 11480 20757
rect 13912 20791 13964 20800
rect 13912 20757 13921 20791
rect 13921 20757 13955 20791
rect 13955 20757 13964 20791
rect 13912 20748 13964 20757
rect 14924 20791 14976 20800
rect 14924 20757 14933 20791
rect 14933 20757 14967 20791
rect 14967 20757 14976 20791
rect 14924 20748 14976 20757
rect 15752 20791 15804 20800
rect 15752 20757 15761 20791
rect 15761 20757 15795 20791
rect 15795 20757 15804 20791
rect 15752 20748 15804 20757
rect 16672 20748 16724 20800
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 17040 20748 17092 20800
rect 17592 20748 17644 20800
rect 17684 20748 17736 20800
rect 18420 20748 18472 20800
rect 26240 20816 26292 20868
rect 26608 20816 26660 20868
rect 31852 20859 31904 20868
rect 31852 20825 31861 20859
rect 31861 20825 31895 20859
rect 31895 20825 31904 20859
rect 31852 20816 31904 20825
rect 21088 20748 21140 20800
rect 21180 20791 21232 20800
rect 21180 20757 21189 20791
rect 21189 20757 21223 20791
rect 21223 20757 21232 20791
rect 21180 20748 21232 20757
rect 22468 20791 22520 20800
rect 22468 20757 22477 20791
rect 22477 20757 22511 20791
rect 22511 20757 22520 20791
rect 22468 20748 22520 20757
rect 22560 20791 22612 20800
rect 22560 20757 22569 20791
rect 22569 20757 22603 20791
rect 22603 20757 22612 20791
rect 22560 20748 22612 20757
rect 22652 20748 22704 20800
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 23940 20748 23992 20800
rect 30656 20748 30708 20800
rect 31208 20791 31260 20800
rect 31208 20757 31217 20791
rect 31217 20757 31251 20791
rect 31251 20757 31260 20791
rect 31208 20748 31260 20757
rect 31944 20791 31996 20800
rect 31944 20757 31953 20791
rect 31953 20757 31987 20791
rect 31987 20757 31996 20791
rect 31944 20748 31996 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 7012 20544 7064 20596
rect 8392 20544 8444 20596
rect 9496 20544 9548 20596
rect 3884 20476 3936 20528
rect 4252 20476 4304 20528
rect 5724 20476 5776 20528
rect 7104 20476 7156 20528
rect 8760 20519 8812 20528
rect 8760 20485 8769 20519
rect 8769 20485 8803 20519
rect 8803 20485 8812 20519
rect 8760 20476 8812 20485
rect 11336 20544 11388 20596
rect 11796 20519 11848 20528
rect 11796 20485 11805 20519
rect 11805 20485 11839 20519
rect 11839 20485 11848 20519
rect 11796 20476 11848 20485
rect 12440 20476 12492 20528
rect 13544 20476 13596 20528
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 3424 20451 3476 20460
rect 3424 20417 3433 20451
rect 3433 20417 3467 20451
rect 3467 20417 3476 20451
rect 3424 20408 3476 20417
rect 4988 20408 5040 20460
rect 2872 20340 2924 20392
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 5724 20383 5776 20392
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 5816 20383 5868 20392
rect 5816 20349 5825 20383
rect 5825 20349 5859 20383
rect 5859 20349 5868 20383
rect 5816 20340 5868 20349
rect 6092 20408 6144 20460
rect 7380 20408 7432 20460
rect 9128 20408 9180 20460
rect 15292 20476 15344 20528
rect 15568 20476 15620 20528
rect 16120 20587 16172 20596
rect 16120 20553 16129 20587
rect 16129 20553 16163 20587
rect 16163 20553 16172 20587
rect 16120 20544 16172 20553
rect 16580 20544 16632 20596
rect 16764 20544 16816 20596
rect 16948 20544 17000 20596
rect 18328 20544 18380 20596
rect 18604 20544 18656 20596
rect 19064 20544 19116 20596
rect 19432 20544 19484 20596
rect 8944 20340 8996 20392
rect 5632 20272 5684 20324
rect 7104 20204 7156 20256
rect 7380 20204 7432 20256
rect 8024 20204 8076 20256
rect 8392 20247 8444 20256
rect 8392 20213 8401 20247
rect 8401 20213 8435 20247
rect 8435 20213 8444 20247
rect 8392 20204 8444 20213
rect 10968 20340 11020 20392
rect 12532 20340 12584 20392
rect 16028 20451 16080 20460
rect 16028 20417 16037 20451
rect 16037 20417 16071 20451
rect 16071 20417 16080 20451
rect 16028 20408 16080 20417
rect 9680 20204 9732 20256
rect 11152 20247 11204 20256
rect 11152 20213 11161 20247
rect 11161 20213 11195 20247
rect 11195 20213 11204 20247
rect 11152 20204 11204 20213
rect 11244 20204 11296 20256
rect 12716 20204 12768 20256
rect 14004 20383 14056 20392
rect 14004 20349 14013 20383
rect 14013 20349 14047 20383
rect 14047 20349 14056 20383
rect 14004 20340 14056 20349
rect 14740 20340 14792 20392
rect 15200 20340 15252 20392
rect 17592 20408 17644 20460
rect 21456 20476 21508 20528
rect 22468 20544 22520 20596
rect 23756 20544 23808 20596
rect 24492 20476 24544 20528
rect 26056 20544 26108 20596
rect 27160 20544 27212 20596
rect 27252 20544 27304 20596
rect 29552 20544 29604 20596
rect 26148 20476 26200 20528
rect 30932 20587 30984 20596
rect 30932 20553 30941 20587
rect 30941 20553 30975 20587
rect 30975 20553 30984 20587
rect 30932 20544 30984 20553
rect 22008 20451 22060 20460
rect 22008 20417 22017 20451
rect 22017 20417 22051 20451
rect 22051 20417 22060 20451
rect 22008 20408 22060 20417
rect 23388 20408 23440 20460
rect 24216 20408 24268 20460
rect 25872 20408 25924 20460
rect 27528 20451 27580 20460
rect 27528 20417 27537 20451
rect 27537 20417 27571 20451
rect 27571 20417 27580 20451
rect 27528 20408 27580 20417
rect 18788 20340 18840 20392
rect 15108 20272 15160 20324
rect 16580 20272 16632 20324
rect 16764 20272 16816 20324
rect 17500 20272 17552 20324
rect 20628 20340 20680 20392
rect 24676 20340 24728 20392
rect 25964 20340 26016 20392
rect 29736 20408 29788 20460
rect 36912 20408 36964 20460
rect 28356 20383 28408 20392
rect 28356 20349 28365 20383
rect 28365 20349 28399 20383
rect 28399 20349 28408 20383
rect 28356 20340 28408 20349
rect 30196 20340 30248 20392
rect 30288 20340 30340 20392
rect 31484 20340 31536 20392
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 15568 20204 15620 20256
rect 16120 20204 16172 20256
rect 18328 20204 18380 20256
rect 22560 20272 22612 20324
rect 27620 20272 27672 20324
rect 27896 20272 27948 20324
rect 25688 20204 25740 20256
rect 26516 20204 26568 20256
rect 27712 20204 27764 20256
rect 28632 20204 28684 20256
rect 30196 20204 30248 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 3332 20043 3384 20052
rect 3332 20009 3341 20043
rect 3341 20009 3375 20043
rect 3375 20009 3384 20043
rect 3332 20000 3384 20009
rect 5264 20000 5316 20052
rect 7564 20000 7616 20052
rect 8024 20000 8076 20052
rect 8576 20000 8628 20052
rect 9864 20000 9916 20052
rect 11336 20043 11388 20052
rect 11336 20009 11345 20043
rect 11345 20009 11379 20043
rect 11379 20009 11388 20043
rect 11336 20000 11388 20009
rect 11888 20000 11940 20052
rect 13820 20000 13872 20052
rect 14188 20000 14240 20052
rect 17592 20000 17644 20052
rect 19800 20000 19852 20052
rect 21272 20000 21324 20052
rect 24584 20000 24636 20052
rect 3332 19864 3384 19916
rect 5448 19864 5500 19916
rect 8944 19864 8996 19916
rect 12440 19932 12492 19984
rect 17040 19932 17092 19984
rect 17224 19975 17276 19984
rect 17224 19941 17233 19975
rect 17233 19941 17267 19975
rect 17267 19941 17276 19975
rect 17224 19932 17276 19941
rect 13360 19864 13412 19916
rect 15476 19864 15528 19916
rect 16948 19907 17000 19916
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 16948 19864 17000 19873
rect 17684 19907 17736 19916
rect 17684 19873 17693 19907
rect 17693 19873 17727 19907
rect 17727 19873 17736 19907
rect 17684 19864 17736 19873
rect 18972 19932 19024 19984
rect 19248 19932 19300 19984
rect 22836 19932 22888 19984
rect 18788 19864 18840 19916
rect 21180 19864 21232 19916
rect 23848 19907 23900 19916
rect 4068 19796 4120 19848
rect 11060 19796 11112 19848
rect 14464 19796 14516 19848
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 3884 19728 3936 19780
rect 4804 19771 4856 19780
rect 4804 19737 4813 19771
rect 4813 19737 4847 19771
rect 4847 19737 4856 19771
rect 4804 19728 4856 19737
rect 5264 19728 5316 19780
rect 6736 19728 6788 19780
rect 7472 19728 7524 19780
rect 3700 19660 3752 19712
rect 6920 19660 6972 19712
rect 9496 19728 9548 19780
rect 11152 19728 11204 19780
rect 10968 19660 11020 19712
rect 13268 19728 13320 19780
rect 11796 19703 11848 19712
rect 11796 19669 11805 19703
rect 11805 19669 11839 19703
rect 11839 19669 11848 19703
rect 11796 19660 11848 19669
rect 11888 19660 11940 19712
rect 13176 19660 13228 19712
rect 13360 19703 13412 19712
rect 13360 19669 13369 19703
rect 13369 19669 13403 19703
rect 13403 19669 13412 19703
rect 13360 19660 13412 19669
rect 14188 19660 14240 19712
rect 15016 19660 15068 19712
rect 16120 19728 16172 19780
rect 18328 19728 18380 19780
rect 19064 19796 19116 19848
rect 19708 19796 19760 19848
rect 19432 19728 19484 19780
rect 19524 19728 19576 19780
rect 20444 19728 20496 19780
rect 21548 19728 21600 19780
rect 16396 19660 16448 19712
rect 18420 19703 18472 19712
rect 18420 19669 18429 19703
rect 18429 19669 18463 19703
rect 18463 19669 18472 19703
rect 18420 19660 18472 19669
rect 19892 19660 19944 19712
rect 21456 19660 21508 19712
rect 23848 19873 23857 19907
rect 23857 19873 23891 19907
rect 23891 19873 23900 19907
rect 23848 19864 23900 19873
rect 30840 20000 30892 20052
rect 49240 20000 49292 20052
rect 27988 19932 28040 19984
rect 29644 19932 29696 19984
rect 33508 19932 33560 19984
rect 25228 19907 25280 19916
rect 25228 19873 25237 19907
rect 25237 19873 25271 19907
rect 25271 19873 25280 19907
rect 25228 19864 25280 19873
rect 22284 19796 22336 19848
rect 23756 19839 23808 19848
rect 23756 19805 23765 19839
rect 23765 19805 23799 19839
rect 23799 19805 23808 19839
rect 23756 19796 23808 19805
rect 24768 19796 24820 19848
rect 28724 19864 28776 19916
rect 25780 19796 25832 19848
rect 27252 19796 27304 19848
rect 27988 19796 28040 19848
rect 28540 19796 28592 19848
rect 29920 19839 29972 19848
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 37188 19796 37240 19848
rect 22744 19771 22796 19780
rect 22744 19737 22753 19771
rect 22753 19737 22787 19771
rect 22787 19737 22796 19771
rect 22744 19728 22796 19737
rect 23572 19728 23624 19780
rect 26148 19771 26200 19780
rect 26148 19737 26157 19771
rect 26157 19737 26191 19771
rect 26191 19737 26200 19771
rect 26148 19728 26200 19737
rect 26608 19728 26660 19780
rect 23296 19703 23348 19712
rect 23296 19669 23305 19703
rect 23305 19669 23339 19703
rect 23339 19669 23348 19703
rect 23296 19660 23348 19669
rect 23664 19703 23716 19712
rect 23664 19669 23673 19703
rect 23673 19669 23707 19703
rect 23707 19669 23716 19703
rect 23664 19660 23716 19669
rect 25044 19703 25096 19712
rect 25044 19669 25053 19703
rect 25053 19669 25087 19703
rect 25087 19669 25096 19703
rect 25044 19660 25096 19669
rect 25872 19660 25924 19712
rect 30840 19728 30892 19780
rect 27896 19660 27948 19712
rect 28356 19660 28408 19712
rect 30472 19660 30524 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 4896 19456 4948 19508
rect 4988 19456 5040 19508
rect 6000 19456 6052 19508
rect 4160 19388 4212 19440
rect 10324 19456 10376 19508
rect 7564 19388 7616 19440
rect 10876 19499 10928 19508
rect 10876 19465 10885 19499
rect 10885 19465 10919 19499
rect 10919 19465 10928 19499
rect 10876 19456 10928 19465
rect 12164 19456 12216 19508
rect 14556 19456 14608 19508
rect 14832 19499 14884 19508
rect 14832 19465 14841 19499
rect 14841 19465 14875 19499
rect 14875 19465 14884 19499
rect 14832 19456 14884 19465
rect 17408 19456 17460 19508
rect 11428 19388 11480 19440
rect 2872 19320 2924 19372
rect 3608 19363 3660 19372
rect 3608 19329 3617 19363
rect 3617 19329 3651 19363
rect 3651 19329 3660 19363
rect 3608 19320 3660 19329
rect 5264 19320 5316 19372
rect 5448 19294 5500 19346
rect 6920 19320 6972 19372
rect 8668 19320 8720 19372
rect 10784 19363 10836 19372
rect 10784 19329 10793 19363
rect 10793 19329 10827 19363
rect 10827 19329 10836 19363
rect 10784 19320 10836 19329
rect 11888 19388 11940 19440
rect 14464 19388 14516 19440
rect 5908 19295 5960 19304
rect 5908 19261 5917 19295
rect 5917 19261 5951 19295
rect 5951 19261 5960 19295
rect 5908 19252 5960 19261
rect 5356 19184 5408 19236
rect 10968 19295 11020 19304
rect 10968 19261 10977 19295
rect 10977 19261 11011 19295
rect 11011 19261 11020 19295
rect 10968 19252 11020 19261
rect 12348 19252 12400 19304
rect 13268 19320 13320 19372
rect 13176 19252 13228 19304
rect 14096 19320 14148 19372
rect 15660 19363 15712 19372
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 17316 19320 17368 19372
rect 17500 19320 17552 19372
rect 18972 19456 19024 19508
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 19248 19456 19300 19508
rect 23296 19456 23348 19508
rect 23572 19456 23624 19508
rect 18052 19388 18104 19440
rect 18512 19388 18564 19440
rect 18788 19388 18840 19440
rect 21548 19388 21600 19440
rect 21824 19388 21876 19440
rect 22652 19388 22704 19440
rect 18144 19320 18196 19372
rect 19064 19320 19116 19372
rect 21916 19320 21968 19372
rect 25872 19456 25924 19508
rect 26240 19456 26292 19508
rect 27160 19456 27212 19508
rect 25504 19388 25556 19440
rect 26608 19388 26660 19440
rect 26976 19388 27028 19440
rect 27252 19431 27304 19440
rect 27252 19397 27261 19431
rect 27261 19397 27295 19431
rect 27295 19397 27304 19431
rect 27252 19388 27304 19397
rect 28632 19388 28684 19440
rect 32036 19388 32088 19440
rect 14648 19252 14700 19304
rect 14924 19295 14976 19304
rect 14924 19261 14933 19295
rect 14933 19261 14967 19295
rect 14967 19261 14976 19295
rect 14924 19252 14976 19261
rect 15108 19252 15160 19304
rect 6644 19184 6696 19236
rect 8392 19184 8444 19236
rect 9496 19184 9548 19236
rect 11704 19184 11756 19236
rect 4804 19116 4856 19168
rect 6368 19116 6420 19168
rect 11060 19116 11112 19168
rect 16304 19252 16356 19304
rect 16856 19252 16908 19304
rect 17592 19252 17644 19304
rect 18052 19252 18104 19304
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 20628 19252 20680 19304
rect 22652 19295 22704 19304
rect 22652 19261 22661 19295
rect 22661 19261 22695 19295
rect 22695 19261 22704 19295
rect 22652 19252 22704 19261
rect 23388 19252 23440 19304
rect 24860 19252 24912 19304
rect 16488 19184 16540 19236
rect 21824 19184 21876 19236
rect 13176 19116 13228 19168
rect 14188 19116 14240 19168
rect 14372 19159 14424 19168
rect 14372 19125 14381 19159
rect 14381 19125 14415 19159
rect 14415 19125 14424 19159
rect 14372 19116 14424 19125
rect 14464 19116 14516 19168
rect 16028 19116 16080 19168
rect 16120 19116 16172 19168
rect 16580 19116 16632 19168
rect 16856 19116 16908 19168
rect 17408 19116 17460 19168
rect 18144 19116 18196 19168
rect 18880 19116 18932 19168
rect 20996 19116 21048 19168
rect 22008 19159 22060 19168
rect 22008 19125 22017 19159
rect 22017 19125 22051 19159
rect 22051 19125 22060 19159
rect 22008 19116 22060 19125
rect 22192 19184 22244 19236
rect 29644 19320 29696 19372
rect 30656 19363 30708 19372
rect 30656 19329 30665 19363
rect 30665 19329 30699 19363
rect 30699 19329 30708 19363
rect 30656 19320 30708 19329
rect 25780 19295 25832 19304
rect 25780 19261 25789 19295
rect 25789 19261 25823 19295
rect 25823 19261 25832 19295
rect 25780 19252 25832 19261
rect 26884 19252 26936 19304
rect 27804 19252 27856 19304
rect 30840 19252 30892 19304
rect 25320 19184 25372 19236
rect 27436 19227 27488 19236
rect 27436 19193 27445 19227
rect 27445 19193 27479 19227
rect 27479 19193 27488 19227
rect 27436 19184 27488 19193
rect 22560 19116 22612 19168
rect 23756 19116 23808 19168
rect 25228 19116 25280 19168
rect 26608 19116 26660 19168
rect 27620 19116 27672 19168
rect 28356 19116 28408 19168
rect 28632 19116 28684 19168
rect 30288 19116 30340 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 9404 18955 9456 18964
rect 9404 18921 9413 18955
rect 9413 18921 9447 18955
rect 9447 18921 9456 18955
rect 9404 18912 9456 18921
rect 9772 18912 9824 18964
rect 12256 18912 12308 18964
rect 14372 18912 14424 18964
rect 14832 18912 14884 18964
rect 22008 18912 22060 18964
rect 22652 18912 22704 18964
rect 8484 18776 8536 18828
rect 4436 18708 4488 18760
rect 4620 18751 4672 18760
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 4620 18708 4672 18717
rect 9312 18776 9364 18828
rect 9772 18776 9824 18828
rect 9956 18819 10008 18828
rect 9956 18785 9965 18819
rect 9965 18785 9999 18819
rect 9999 18785 10008 18819
rect 9956 18776 10008 18785
rect 10232 18776 10284 18828
rect 10968 18776 11020 18828
rect 11152 18776 11204 18828
rect 14464 18844 14516 18896
rect 16488 18844 16540 18896
rect 15108 18776 15160 18828
rect 16212 18776 16264 18828
rect 16672 18776 16724 18828
rect 18328 18844 18380 18896
rect 19340 18844 19392 18896
rect 20720 18844 20772 18896
rect 25136 18887 25188 18896
rect 25136 18853 25145 18887
rect 25145 18853 25179 18887
rect 25179 18853 25188 18887
rect 25688 18912 25740 18964
rect 26148 18912 26200 18964
rect 27252 18912 27304 18964
rect 47032 18912 47084 18964
rect 25136 18844 25188 18853
rect 26792 18844 26844 18896
rect 19708 18776 19760 18828
rect 21456 18819 21508 18828
rect 21456 18785 21465 18819
rect 21465 18785 21499 18819
rect 21499 18785 21508 18819
rect 21456 18776 21508 18785
rect 21548 18776 21600 18828
rect 9128 18708 9180 18760
rect 10048 18708 10100 18760
rect 11336 18708 11388 18760
rect 11888 18708 11940 18760
rect 13360 18708 13412 18760
rect 14832 18708 14884 18760
rect 17040 18708 17092 18760
rect 18052 18708 18104 18760
rect 18604 18751 18656 18760
rect 18604 18717 18613 18751
rect 18613 18717 18647 18751
rect 18647 18717 18656 18751
rect 18604 18708 18656 18717
rect 18880 18708 18932 18760
rect 2780 18683 2832 18692
rect 2780 18649 2789 18683
rect 2789 18649 2823 18683
rect 2823 18649 2832 18683
rect 2780 18640 2832 18649
rect 3056 18640 3108 18692
rect 4068 18640 4120 18692
rect 4804 18640 4856 18692
rect 3332 18615 3384 18624
rect 3332 18581 3341 18615
rect 3341 18581 3375 18615
rect 3375 18581 3384 18615
rect 3332 18572 3384 18581
rect 5448 18640 5500 18692
rect 7196 18640 7248 18692
rect 7564 18640 7616 18692
rect 8576 18640 8628 18692
rect 6184 18572 6236 18624
rect 6368 18615 6420 18624
rect 6368 18581 6377 18615
rect 6377 18581 6411 18615
rect 6411 18581 6420 18615
rect 6368 18572 6420 18581
rect 8760 18572 8812 18624
rect 8944 18640 8996 18692
rect 9864 18572 9916 18624
rect 10692 18640 10744 18692
rect 11336 18572 11388 18624
rect 11612 18572 11664 18624
rect 12072 18615 12124 18624
rect 12072 18581 12081 18615
rect 12081 18581 12115 18615
rect 12115 18581 12124 18615
rect 12072 18572 12124 18581
rect 13176 18640 13228 18692
rect 13544 18683 13596 18692
rect 13544 18649 13553 18683
rect 13553 18649 13587 18683
rect 13587 18649 13596 18683
rect 13544 18640 13596 18649
rect 15292 18572 15344 18624
rect 16028 18640 16080 18692
rect 16396 18572 16448 18624
rect 20076 18640 20128 18692
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 16948 18572 17000 18581
rect 17592 18572 17644 18624
rect 18604 18572 18656 18624
rect 19524 18572 19576 18624
rect 19800 18572 19852 18624
rect 20812 18615 20864 18624
rect 20812 18581 20821 18615
rect 20821 18581 20855 18615
rect 20855 18581 20864 18615
rect 20812 18572 20864 18581
rect 22560 18708 22612 18760
rect 23664 18776 23716 18828
rect 25780 18776 25832 18828
rect 26240 18776 26292 18828
rect 30196 18819 30248 18828
rect 30196 18785 30205 18819
rect 30205 18785 30239 18819
rect 30239 18785 30248 18819
rect 30196 18776 30248 18785
rect 23572 18751 23624 18760
rect 23572 18717 23581 18751
rect 23581 18717 23615 18751
rect 23615 18717 23624 18751
rect 23572 18708 23624 18717
rect 23756 18708 23808 18760
rect 25136 18708 25188 18760
rect 27712 18708 27764 18760
rect 29828 18708 29880 18760
rect 30840 18819 30892 18828
rect 30840 18785 30849 18819
rect 30849 18785 30883 18819
rect 30883 18785 30892 18819
rect 30840 18776 30892 18785
rect 46940 18776 46992 18828
rect 22100 18572 22152 18624
rect 23388 18615 23440 18624
rect 23388 18581 23397 18615
rect 23397 18581 23431 18615
rect 23431 18581 23440 18615
rect 23388 18572 23440 18581
rect 23480 18572 23532 18624
rect 23848 18572 23900 18624
rect 25964 18640 26016 18692
rect 26976 18640 27028 18692
rect 30656 18640 30708 18692
rect 29736 18615 29788 18624
rect 29736 18581 29745 18615
rect 29745 18581 29779 18615
rect 29779 18581 29788 18615
rect 29736 18572 29788 18581
rect 30104 18615 30156 18624
rect 30104 18581 30113 18615
rect 30113 18581 30147 18615
rect 30147 18581 30156 18615
rect 30104 18572 30156 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 5632 18368 5684 18420
rect 6920 18368 6972 18420
rect 8944 18368 8996 18420
rect 10232 18368 10284 18420
rect 11888 18368 11940 18420
rect 5908 18300 5960 18352
rect 7472 18300 7524 18352
rect 9588 18300 9640 18352
rect 5632 18275 5684 18284
rect 5632 18241 5641 18275
rect 5641 18241 5675 18275
rect 5675 18241 5684 18275
rect 5632 18232 5684 18241
rect 6092 18232 6144 18284
rect 6644 18232 6696 18284
rect 6736 18275 6788 18284
rect 6736 18241 6745 18275
rect 6745 18241 6779 18275
rect 6779 18241 6788 18275
rect 6736 18232 6788 18241
rect 7012 18232 7064 18284
rect 7932 18232 7984 18284
rect 8392 18232 8444 18284
rect 10508 18300 10560 18352
rect 10232 18232 10284 18284
rect 11336 18232 11388 18284
rect 13728 18368 13780 18420
rect 19340 18368 19392 18420
rect 20720 18411 20772 18420
rect 20720 18377 20729 18411
rect 20729 18377 20763 18411
rect 20763 18377 20772 18411
rect 20720 18368 20772 18377
rect 20996 18368 21048 18420
rect 26976 18368 27028 18420
rect 30104 18368 30156 18420
rect 30656 18368 30708 18420
rect 38568 18368 38620 18420
rect 2044 18207 2096 18216
rect 2044 18173 2053 18207
rect 2053 18173 2087 18207
rect 2087 18173 2096 18207
rect 2044 18164 2096 18173
rect 3792 18164 3844 18216
rect 5908 18207 5960 18216
rect 5908 18173 5917 18207
rect 5917 18173 5951 18207
rect 5951 18173 5960 18207
rect 5908 18164 5960 18173
rect 7288 18207 7340 18216
rect 7288 18173 7297 18207
rect 7297 18173 7331 18207
rect 7331 18173 7340 18207
rect 7288 18164 7340 18173
rect 8576 18164 8628 18216
rect 9496 18164 9548 18216
rect 14004 18300 14056 18352
rect 14556 18300 14608 18352
rect 16028 18300 16080 18352
rect 6276 18096 6328 18148
rect 7012 18096 7064 18148
rect 7932 18096 7984 18148
rect 10692 18096 10744 18148
rect 11888 18096 11940 18148
rect 1124 18028 1176 18080
rect 6736 18028 6788 18080
rect 9864 18028 9916 18080
rect 10140 18028 10192 18080
rect 12072 18028 12124 18080
rect 13176 18207 13228 18216
rect 13176 18173 13185 18207
rect 13185 18173 13219 18207
rect 13219 18173 13228 18207
rect 15200 18232 15252 18284
rect 16580 18232 16632 18284
rect 19708 18300 19760 18352
rect 19800 18300 19852 18352
rect 21088 18343 21140 18352
rect 21088 18309 21097 18343
rect 21097 18309 21131 18343
rect 21131 18309 21140 18343
rect 21088 18300 21140 18309
rect 13176 18164 13228 18173
rect 15108 18164 15160 18216
rect 12808 18096 12860 18148
rect 15016 18139 15068 18148
rect 15016 18105 15025 18139
rect 15025 18105 15059 18139
rect 15059 18105 15068 18139
rect 15016 18096 15068 18105
rect 16948 18164 17000 18216
rect 17500 18207 17552 18216
rect 17500 18173 17509 18207
rect 17509 18173 17543 18207
rect 17543 18173 17552 18207
rect 17500 18164 17552 18173
rect 17592 18164 17644 18216
rect 19340 18164 19392 18216
rect 23480 18300 23532 18352
rect 25136 18300 25188 18352
rect 25320 18343 25372 18352
rect 25320 18309 25329 18343
rect 25329 18309 25363 18343
rect 25363 18309 25372 18343
rect 25320 18300 25372 18309
rect 26056 18343 26108 18352
rect 26056 18309 26065 18343
rect 26065 18309 26099 18343
rect 26099 18309 26108 18343
rect 26056 18300 26108 18309
rect 28632 18300 28684 18352
rect 29644 18300 29696 18352
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 27804 18232 27856 18284
rect 30656 18275 30708 18284
rect 30656 18241 30665 18275
rect 30665 18241 30699 18275
rect 30699 18241 30708 18275
rect 30656 18232 30708 18241
rect 31024 18232 31076 18284
rect 20076 18207 20128 18216
rect 20076 18173 20085 18207
rect 20085 18173 20119 18207
rect 20119 18173 20128 18207
rect 20076 18164 20128 18173
rect 20812 18164 20864 18216
rect 20720 18096 20772 18148
rect 22468 18164 22520 18216
rect 22928 18164 22980 18216
rect 12624 18028 12676 18080
rect 13544 18028 13596 18080
rect 15752 18028 15804 18080
rect 16396 18071 16448 18080
rect 16396 18037 16405 18071
rect 16405 18037 16439 18071
rect 16439 18037 16448 18071
rect 16396 18028 16448 18037
rect 17684 18028 17736 18080
rect 19708 18028 19760 18080
rect 22836 18028 22888 18080
rect 25228 18164 25280 18216
rect 27068 18164 27120 18216
rect 24492 18096 24544 18148
rect 26792 18096 26844 18148
rect 30380 18096 30432 18148
rect 37740 18164 37792 18216
rect 24676 18028 24728 18080
rect 27344 18028 27396 18080
rect 29828 18071 29880 18080
rect 29828 18037 29837 18071
rect 29837 18037 29871 18071
rect 29871 18037 29880 18071
rect 29828 18028 29880 18037
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 8392 17824 8444 17876
rect 8944 17824 8996 17876
rect 1860 17756 1912 17808
rect 6184 17756 6236 17808
rect 7196 17756 7248 17808
rect 7564 17756 7616 17808
rect 7840 17799 7892 17808
rect 7840 17765 7849 17799
rect 7849 17765 7883 17799
rect 7883 17765 7892 17799
rect 7840 17756 7892 17765
rect 10140 17824 10192 17876
rect 10324 17824 10376 17876
rect 12348 17824 12400 17876
rect 15200 17824 15252 17876
rect 16396 17824 16448 17876
rect 16672 17824 16724 17876
rect 21180 17824 21232 17876
rect 21272 17824 21324 17876
rect 21732 17824 21784 17876
rect 23756 17824 23808 17876
rect 1124 17688 1176 17740
rect 9772 17756 9824 17808
rect 11888 17756 11940 17808
rect 13268 17756 13320 17808
rect 16212 17756 16264 17808
rect 17592 17756 17644 17808
rect 9680 17688 9732 17740
rect 10048 17688 10100 17740
rect 12900 17688 12952 17740
rect 13636 17688 13688 17740
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 16948 17688 17000 17740
rect 18972 17688 19024 17740
rect 19616 17688 19668 17740
rect 20352 17688 20404 17740
rect 23756 17688 23808 17740
rect 3792 17663 3844 17672
rect 3792 17629 3801 17663
rect 3801 17629 3835 17663
rect 3835 17629 3844 17663
rect 3792 17620 3844 17629
rect 4160 17620 4212 17672
rect 4620 17620 4672 17672
rect 7104 17620 7156 17672
rect 8944 17620 8996 17672
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 9496 17620 9548 17672
rect 11704 17663 11756 17672
rect 11704 17629 11713 17663
rect 11713 17629 11747 17663
rect 11747 17629 11756 17663
rect 11704 17620 11756 17629
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 19340 17620 19392 17672
rect 22008 17620 22060 17672
rect 23664 17620 23716 17672
rect 1216 17552 1268 17604
rect 4068 17552 4120 17604
rect 4804 17552 4856 17604
rect 5448 17552 5500 17604
rect 7196 17595 7248 17604
rect 7196 17561 7205 17595
rect 7205 17561 7239 17595
rect 7239 17561 7248 17595
rect 7196 17552 7248 17561
rect 9404 17552 9456 17604
rect 12256 17552 12308 17604
rect 13544 17552 13596 17604
rect 14004 17552 14056 17604
rect 7380 17484 7432 17536
rect 8024 17484 8076 17536
rect 14280 17484 14332 17536
rect 14464 17527 14516 17536
rect 14464 17493 14473 17527
rect 14473 17493 14507 17527
rect 14507 17493 14516 17527
rect 14464 17484 14516 17493
rect 15016 17484 15068 17536
rect 15108 17527 15160 17536
rect 15108 17493 15117 17527
rect 15117 17493 15151 17527
rect 15151 17493 15160 17527
rect 15108 17484 15160 17493
rect 15384 17527 15436 17536
rect 15384 17493 15393 17527
rect 15393 17493 15427 17527
rect 15427 17493 15436 17527
rect 15384 17484 15436 17493
rect 16028 17527 16080 17536
rect 16028 17493 16037 17527
rect 16037 17493 16071 17527
rect 16071 17493 16080 17527
rect 16028 17484 16080 17493
rect 16396 17484 16448 17536
rect 20720 17552 20772 17604
rect 18512 17484 18564 17536
rect 20444 17484 20496 17536
rect 20996 17484 21048 17536
rect 21824 17484 21876 17536
rect 22560 17595 22612 17604
rect 22560 17561 22569 17595
rect 22569 17561 22603 17595
rect 22603 17561 22612 17595
rect 22560 17552 22612 17561
rect 26608 17799 26660 17808
rect 26608 17765 26617 17799
rect 26617 17765 26651 17799
rect 26651 17765 26660 17799
rect 26608 17756 26660 17765
rect 28448 17756 28500 17808
rect 24676 17688 24728 17740
rect 25780 17688 25832 17740
rect 27804 17688 27856 17740
rect 29644 17688 29696 17740
rect 30288 17731 30340 17740
rect 30288 17697 30297 17731
rect 30297 17697 30331 17731
rect 30331 17697 30340 17731
rect 30288 17688 30340 17697
rect 29092 17620 29144 17672
rect 30840 17620 30892 17672
rect 31300 17663 31352 17672
rect 31300 17629 31309 17663
rect 31309 17629 31343 17663
rect 31343 17629 31352 17663
rect 31300 17620 31352 17629
rect 37372 17620 37424 17672
rect 25136 17595 25188 17604
rect 25136 17561 25145 17595
rect 25145 17561 25179 17595
rect 25179 17561 25188 17595
rect 25136 17552 25188 17561
rect 26976 17552 27028 17604
rect 27344 17595 27396 17604
rect 27344 17561 27353 17595
rect 27353 17561 27387 17595
rect 27387 17561 27396 17595
rect 27344 17552 27396 17561
rect 29644 17552 29696 17604
rect 24400 17527 24452 17536
rect 24400 17493 24409 17527
rect 24409 17493 24443 17527
rect 24443 17493 24452 17527
rect 30932 17552 30984 17604
rect 24400 17484 24452 17493
rect 30196 17527 30248 17536
rect 30196 17493 30205 17527
rect 30205 17493 30239 17527
rect 30239 17493 30248 17527
rect 30196 17484 30248 17493
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 3976 17280 4028 17332
rect 4896 17323 4948 17332
rect 4896 17289 4905 17323
rect 4905 17289 4939 17323
rect 4939 17289 4948 17323
rect 4896 17280 4948 17289
rect 6828 17323 6880 17332
rect 6828 17289 6837 17323
rect 6837 17289 6871 17323
rect 6871 17289 6880 17323
rect 6828 17280 6880 17289
rect 7748 17280 7800 17332
rect 4344 17255 4396 17264
rect 4344 17221 4353 17255
rect 4353 17221 4387 17255
rect 4387 17221 4396 17255
rect 4344 17212 4396 17221
rect 7288 17212 7340 17264
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 12440 17280 12492 17332
rect 9588 17212 9640 17264
rect 13360 17280 13412 17332
rect 13728 17323 13780 17332
rect 13728 17289 13737 17323
rect 13737 17289 13771 17323
rect 13771 17289 13780 17323
rect 13728 17280 13780 17289
rect 14280 17280 14332 17332
rect 16212 17280 16264 17332
rect 17132 17280 17184 17332
rect 17868 17280 17920 17332
rect 22468 17280 22520 17332
rect 8392 17187 8444 17196
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 1308 17076 1360 17128
rect 3516 17076 3568 17128
rect 4620 17076 4672 17128
rect 5908 17119 5960 17128
rect 5908 17085 5917 17119
rect 5917 17085 5951 17119
rect 5951 17085 5960 17119
rect 5908 17076 5960 17085
rect 6368 17076 6420 17128
rect 6460 17119 6512 17128
rect 6460 17085 6469 17119
rect 6469 17085 6503 17119
rect 6503 17085 6512 17119
rect 6460 17076 6512 17085
rect 7564 17076 7616 17128
rect 8576 17076 8628 17128
rect 8760 17144 8812 17196
rect 9312 17144 9364 17196
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 12808 17212 12860 17264
rect 10324 17076 10376 17128
rect 11796 17187 11848 17196
rect 11796 17153 11805 17187
rect 11805 17153 11839 17187
rect 11839 17153 11848 17187
rect 11796 17144 11848 17153
rect 12256 17076 12308 17128
rect 13912 17144 13964 17196
rect 17776 17212 17828 17264
rect 18144 17212 18196 17264
rect 18512 17212 18564 17264
rect 15660 17187 15712 17196
rect 15660 17153 15669 17187
rect 15669 17153 15703 17187
rect 15703 17153 15712 17187
rect 15660 17144 15712 17153
rect 16672 17144 16724 17196
rect 17224 17187 17276 17196
rect 17224 17153 17233 17187
rect 17233 17153 17267 17187
rect 17267 17153 17276 17187
rect 17224 17144 17276 17153
rect 19800 17144 19852 17196
rect 8760 17008 8812 17060
rect 12348 17008 12400 17060
rect 15292 17076 15344 17128
rect 15844 17076 15896 17128
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 22560 17212 22612 17264
rect 20628 17144 20680 17196
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 21272 17144 21324 17196
rect 24400 17280 24452 17332
rect 23756 17212 23808 17264
rect 29092 17280 29144 17332
rect 29644 17280 29696 17332
rect 30196 17280 30248 17332
rect 30840 17323 30892 17332
rect 30840 17289 30849 17323
rect 30849 17289 30883 17323
rect 30883 17289 30892 17323
rect 30840 17280 30892 17289
rect 30932 17323 30984 17332
rect 30932 17289 30941 17323
rect 30941 17289 30975 17323
rect 30975 17289 30984 17323
rect 30932 17280 30984 17289
rect 26976 17212 27028 17264
rect 13452 17008 13504 17060
rect 17040 17008 17092 17060
rect 3332 16940 3384 16992
rect 9772 16940 9824 16992
rect 10508 16940 10560 16992
rect 10876 16983 10928 16992
rect 10876 16949 10885 16983
rect 10885 16949 10919 16983
rect 10919 16949 10928 16983
rect 10876 16940 10928 16949
rect 11612 16940 11664 16992
rect 12072 16940 12124 16992
rect 13728 16940 13780 16992
rect 15292 16940 15344 16992
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 17500 16940 17552 16992
rect 20076 17008 20128 17060
rect 21732 17076 21784 17128
rect 22560 17119 22612 17128
rect 22560 17085 22569 17119
rect 22569 17085 22603 17119
rect 22603 17085 22612 17119
rect 22560 17076 22612 17085
rect 23756 17119 23808 17128
rect 23756 17085 23765 17119
rect 23765 17085 23799 17119
rect 23799 17085 23808 17119
rect 23756 17076 23808 17085
rect 24492 17144 24544 17196
rect 24676 17187 24728 17196
rect 24676 17153 24685 17187
rect 24685 17153 24719 17187
rect 24719 17153 24728 17187
rect 24676 17144 24728 17153
rect 27804 17187 27856 17196
rect 27804 17153 27813 17187
rect 27813 17153 27847 17187
rect 27847 17153 27856 17187
rect 27804 17144 27856 17153
rect 37280 17212 37332 17264
rect 48504 17212 48556 17264
rect 31760 17144 31812 17196
rect 20168 16983 20220 16992
rect 20168 16949 20177 16983
rect 20177 16949 20211 16983
rect 20211 16949 20220 16983
rect 20168 16940 20220 16949
rect 20628 16940 20680 16992
rect 20720 16983 20772 16992
rect 20720 16949 20729 16983
rect 20729 16949 20763 16983
rect 20763 16949 20772 16983
rect 20720 16940 20772 16949
rect 22192 17008 22244 17060
rect 27620 17076 27672 17128
rect 30288 17076 30340 17128
rect 30196 17008 30248 17060
rect 21548 16940 21600 16992
rect 21732 16940 21784 16992
rect 22560 16940 22612 16992
rect 23296 16983 23348 16992
rect 23296 16949 23305 16983
rect 23305 16949 23339 16983
rect 23339 16949 23348 16983
rect 23296 16940 23348 16949
rect 25320 16940 25372 16992
rect 25964 16940 26016 16992
rect 27160 16940 27212 16992
rect 30932 17008 30984 17060
rect 47400 17008 47452 17060
rect 47124 16940 47176 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 1768 16736 1820 16788
rect 10876 16736 10928 16788
rect 11704 16736 11756 16788
rect 16856 16736 16908 16788
rect 17132 16736 17184 16788
rect 19708 16736 19760 16788
rect 19800 16736 19852 16788
rect 20996 16736 21048 16788
rect 23756 16736 23808 16788
rect 30196 16736 30248 16788
rect 2136 16668 2188 16720
rect 3516 16668 3568 16720
rect 4068 16668 4120 16720
rect 5540 16668 5592 16720
rect 2320 16600 2372 16652
rect 3332 16600 3384 16652
rect 4528 16643 4580 16652
rect 4528 16609 4537 16643
rect 4537 16609 4571 16643
rect 4571 16609 4580 16643
rect 4528 16600 4580 16609
rect 5724 16600 5776 16652
rect 6276 16600 6328 16652
rect 1308 16464 1360 16516
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 10416 16668 10468 16720
rect 11612 16600 11664 16652
rect 12256 16668 12308 16720
rect 12992 16711 13044 16720
rect 12992 16677 13001 16711
rect 13001 16677 13035 16711
rect 13035 16677 13044 16711
rect 12992 16668 13044 16677
rect 13268 16668 13320 16720
rect 13544 16668 13596 16720
rect 12348 16600 12400 16652
rect 12532 16600 12584 16652
rect 18144 16668 18196 16720
rect 21088 16668 21140 16720
rect 21456 16668 21508 16720
rect 25136 16668 25188 16720
rect 14464 16600 14516 16652
rect 16304 16600 16356 16652
rect 17224 16600 17276 16652
rect 7748 16532 7800 16584
rect 5908 16507 5960 16516
rect 5908 16473 5917 16507
rect 5917 16473 5951 16507
rect 5951 16473 5960 16507
rect 5908 16464 5960 16473
rect 7932 16464 7984 16516
rect 8208 16507 8260 16516
rect 8208 16473 8217 16507
rect 8217 16473 8251 16507
rect 8251 16473 8260 16507
rect 8208 16464 8260 16473
rect 8944 16464 8996 16516
rect 6828 16396 6880 16448
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 8116 16396 8168 16448
rect 10416 16575 10468 16584
rect 10416 16541 10425 16575
rect 10425 16541 10459 16575
rect 10459 16541 10468 16575
rect 10416 16532 10468 16541
rect 10508 16575 10560 16584
rect 10508 16541 10517 16575
rect 10517 16541 10551 16575
rect 10551 16541 10560 16575
rect 10508 16532 10560 16541
rect 12808 16464 12860 16516
rect 14648 16532 14700 16584
rect 15384 16575 15436 16584
rect 15384 16541 15393 16575
rect 15393 16541 15427 16575
rect 15427 16541 15436 16575
rect 15384 16532 15436 16541
rect 15568 16532 15620 16584
rect 13544 16464 13596 16516
rect 11244 16439 11296 16448
rect 11244 16405 11253 16439
rect 11253 16405 11287 16439
rect 11287 16405 11296 16439
rect 11244 16396 11296 16405
rect 11888 16396 11940 16448
rect 14372 16439 14424 16448
rect 14372 16405 14381 16439
rect 14381 16405 14415 16439
rect 14415 16405 14424 16439
rect 14372 16396 14424 16405
rect 15568 16396 15620 16448
rect 15936 16532 15988 16584
rect 18512 16600 18564 16652
rect 20352 16600 20404 16652
rect 20720 16600 20772 16652
rect 22560 16643 22612 16652
rect 22560 16609 22569 16643
rect 22569 16609 22603 16643
rect 22603 16609 22612 16643
rect 22560 16600 22612 16609
rect 23756 16643 23808 16652
rect 23756 16609 23765 16643
rect 23765 16609 23799 16643
rect 23799 16609 23808 16643
rect 23756 16600 23808 16609
rect 24584 16600 24636 16652
rect 25228 16600 25280 16652
rect 25780 16600 25832 16652
rect 25964 16643 26016 16652
rect 25964 16609 25973 16643
rect 25973 16609 26007 16643
rect 26007 16609 26016 16643
rect 25964 16600 26016 16609
rect 27068 16643 27120 16652
rect 27068 16609 27077 16643
rect 27077 16609 27111 16643
rect 27111 16609 27120 16643
rect 27068 16600 27120 16609
rect 27160 16643 27212 16652
rect 27160 16609 27169 16643
rect 27169 16609 27203 16643
rect 27203 16609 27212 16643
rect 27160 16600 27212 16609
rect 28724 16600 28776 16652
rect 18328 16532 18380 16584
rect 19156 16532 19208 16584
rect 19432 16575 19484 16584
rect 19432 16541 19441 16575
rect 19441 16541 19475 16575
rect 19475 16541 19484 16575
rect 19432 16532 19484 16541
rect 23296 16532 23348 16584
rect 23664 16532 23716 16584
rect 24492 16532 24544 16584
rect 25044 16532 25096 16584
rect 16396 16439 16448 16448
rect 16396 16405 16405 16439
rect 16405 16405 16439 16439
rect 16439 16405 16448 16439
rect 16396 16396 16448 16405
rect 16856 16396 16908 16448
rect 18328 16396 18380 16448
rect 18604 16396 18656 16448
rect 20996 16464 21048 16516
rect 21180 16464 21232 16516
rect 20076 16396 20128 16448
rect 20720 16396 20772 16448
rect 22376 16396 22428 16448
rect 23848 16396 23900 16448
rect 24584 16396 24636 16448
rect 24676 16439 24728 16448
rect 24676 16405 24685 16439
rect 24685 16405 24719 16439
rect 24719 16405 24728 16439
rect 24676 16396 24728 16405
rect 25320 16464 25372 16516
rect 25504 16464 25556 16516
rect 25136 16439 25188 16448
rect 25136 16405 25145 16439
rect 25145 16405 25179 16439
rect 25179 16405 25188 16439
rect 25688 16439 25740 16448
rect 25136 16396 25188 16405
rect 25688 16405 25697 16439
rect 25697 16405 25731 16439
rect 25731 16405 25740 16439
rect 25688 16396 25740 16405
rect 27620 16532 27672 16584
rect 28356 16532 28408 16584
rect 30840 16600 30892 16652
rect 28448 16464 28500 16516
rect 28264 16396 28316 16448
rect 28540 16396 28592 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 3976 16192 4028 16244
rect 6920 16192 6972 16244
rect 7012 16192 7064 16244
rect 4252 16124 4304 16176
rect 5724 16167 5776 16176
rect 5724 16133 5733 16167
rect 5733 16133 5767 16167
rect 5767 16133 5776 16167
rect 5724 16124 5776 16133
rect 5816 16124 5868 16176
rect 9772 16124 9824 16176
rect 10508 16192 10560 16244
rect 10600 16235 10652 16244
rect 10600 16201 10609 16235
rect 10609 16201 10643 16235
rect 10643 16201 10652 16235
rect 10600 16192 10652 16201
rect 11152 16192 11204 16244
rect 11520 16192 11572 16244
rect 13636 16192 13688 16244
rect 12532 16124 12584 16176
rect 14004 16124 14056 16176
rect 1308 15988 1360 16040
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 3700 16056 3752 16108
rect 7288 16056 7340 16108
rect 8484 16099 8536 16108
rect 8484 16065 8493 16099
rect 8493 16065 8527 16099
rect 8527 16065 8536 16099
rect 8484 16056 8536 16065
rect 4712 15988 4764 16040
rect 6000 15988 6052 16040
rect 6552 15988 6604 16040
rect 6644 16031 6696 16040
rect 6644 15997 6653 16031
rect 6653 15997 6687 16031
rect 6687 15997 6696 16031
rect 6644 15988 6696 15997
rect 7380 15988 7432 16040
rect 7932 16031 7984 16040
rect 7932 15997 7941 16031
rect 7941 15997 7975 16031
rect 7975 15997 7984 16031
rect 7932 15988 7984 15997
rect 6368 15920 6420 15972
rect 8484 15920 8536 15972
rect 9956 15988 10008 16040
rect 10140 15988 10192 16040
rect 10876 15988 10928 16040
rect 10968 15963 11020 15972
rect 10968 15929 10977 15963
rect 10977 15929 11011 15963
rect 11011 15929 11020 15963
rect 10968 15920 11020 15929
rect 5264 15895 5316 15904
rect 5264 15861 5273 15895
rect 5273 15861 5307 15895
rect 5307 15861 5316 15895
rect 5264 15852 5316 15861
rect 7012 15852 7064 15904
rect 11796 15852 11848 15904
rect 11980 16099 12032 16108
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 12256 16031 12308 16040
rect 12256 15997 12265 16031
rect 12265 15997 12299 16031
rect 12299 15997 12308 16031
rect 12256 15988 12308 15997
rect 12348 15988 12400 16040
rect 16488 16124 16540 16176
rect 16672 16192 16724 16244
rect 16948 16235 17000 16244
rect 16948 16201 16957 16235
rect 16957 16201 16991 16235
rect 16991 16201 17000 16235
rect 16948 16192 17000 16201
rect 17132 16235 17184 16244
rect 17132 16201 17141 16235
rect 17141 16201 17175 16235
rect 17175 16201 17184 16235
rect 17132 16192 17184 16201
rect 17500 16192 17552 16244
rect 17868 16235 17920 16244
rect 17868 16201 17877 16235
rect 17877 16201 17911 16235
rect 17911 16201 17920 16235
rect 17868 16192 17920 16201
rect 19708 16235 19760 16244
rect 19708 16201 19717 16235
rect 19717 16201 19751 16235
rect 19751 16201 19760 16235
rect 19708 16192 19760 16201
rect 21180 16192 21232 16244
rect 24952 16192 25004 16244
rect 26976 16235 27028 16244
rect 26976 16201 26985 16235
rect 26985 16201 27019 16235
rect 27019 16201 27028 16235
rect 26976 16192 27028 16201
rect 27620 16192 27672 16244
rect 28356 16192 28408 16244
rect 15016 16056 15068 16108
rect 13636 15920 13688 15972
rect 14924 15988 14976 16040
rect 15476 16031 15528 16040
rect 15476 15997 15485 16031
rect 15485 15997 15519 16031
rect 15519 15997 15528 16031
rect 15476 15988 15528 15997
rect 17592 16056 17644 16108
rect 16580 15988 16632 16040
rect 16672 15988 16724 16040
rect 17868 16056 17920 16108
rect 12440 15852 12492 15904
rect 13728 15852 13780 15904
rect 14924 15852 14976 15904
rect 16396 15852 16448 15904
rect 16580 15852 16632 15904
rect 17592 15920 17644 15972
rect 18696 16056 18748 16108
rect 18880 16099 18932 16108
rect 18880 16065 18889 16099
rect 18889 16065 18923 16099
rect 18923 16065 18932 16099
rect 18880 16056 18932 16065
rect 20444 16099 20496 16108
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 21456 16099 21508 16108
rect 21456 16065 21465 16099
rect 21465 16065 21499 16099
rect 21499 16065 21508 16099
rect 21456 16056 21508 16065
rect 23664 16099 23716 16108
rect 23664 16065 23673 16099
rect 23673 16065 23707 16099
rect 23707 16065 23716 16099
rect 23664 16056 23716 16065
rect 23848 16056 23900 16108
rect 21640 15988 21692 16040
rect 22284 16031 22336 16040
rect 22284 15997 22293 16031
rect 22293 15997 22327 16031
rect 22327 15997 22336 16031
rect 22284 15988 22336 15997
rect 24032 15988 24084 16040
rect 24492 16124 24544 16176
rect 24584 16167 24636 16176
rect 24584 16133 24593 16167
rect 24593 16133 24627 16167
rect 24627 16133 24636 16167
rect 24584 16124 24636 16133
rect 24860 16099 24912 16108
rect 24860 16065 24869 16099
rect 24869 16065 24903 16099
rect 24903 16065 24912 16099
rect 24860 16056 24912 16065
rect 27160 15988 27212 16040
rect 18604 15852 18656 15904
rect 23388 15920 23440 15972
rect 22468 15852 22520 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 1308 15512 1360 15564
rect 3884 15512 3936 15564
rect 5816 15648 5868 15700
rect 7196 15648 7248 15700
rect 7932 15648 7984 15700
rect 8576 15648 8628 15700
rect 8668 15648 8720 15700
rect 6000 15580 6052 15632
rect 5172 15512 5224 15564
rect 7012 15580 7064 15632
rect 8300 15580 8352 15632
rect 9220 15580 9272 15632
rect 6736 15512 6788 15564
rect 6920 15555 6972 15564
rect 6920 15521 6929 15555
rect 6929 15521 6963 15555
rect 6963 15521 6972 15555
rect 6920 15512 6972 15521
rect 7104 15512 7156 15564
rect 3424 15444 3476 15496
rect 2780 15376 2832 15428
rect 3792 15308 3844 15360
rect 4344 15351 4396 15360
rect 4344 15317 4353 15351
rect 4353 15317 4387 15351
rect 4387 15317 4396 15351
rect 4344 15308 4396 15317
rect 5724 15308 5776 15360
rect 6368 15351 6420 15360
rect 6368 15317 6377 15351
rect 6377 15317 6411 15351
rect 6411 15317 6420 15351
rect 6368 15308 6420 15317
rect 6644 15444 6696 15496
rect 8024 15444 8076 15496
rect 7932 15376 7984 15428
rect 8208 15512 8260 15564
rect 8484 15555 8536 15564
rect 8484 15521 8493 15555
rect 8493 15521 8527 15555
rect 8527 15521 8536 15555
rect 8484 15512 8536 15521
rect 12808 15648 12860 15700
rect 13544 15691 13596 15700
rect 13544 15657 13553 15691
rect 13553 15657 13587 15691
rect 13587 15657 13596 15691
rect 13544 15648 13596 15657
rect 14832 15648 14884 15700
rect 15476 15648 15528 15700
rect 15844 15691 15896 15700
rect 15844 15657 15853 15691
rect 15853 15657 15887 15691
rect 15887 15657 15896 15691
rect 15844 15648 15896 15657
rect 10692 15580 10744 15632
rect 20076 15648 20128 15700
rect 10876 15512 10928 15564
rect 13360 15512 13412 15564
rect 14556 15512 14608 15564
rect 9220 15419 9272 15428
rect 9220 15385 9229 15419
rect 9229 15385 9263 15419
rect 9263 15385 9272 15419
rect 9220 15376 9272 15385
rect 9864 15444 9916 15496
rect 11520 15444 11572 15496
rect 11796 15444 11848 15496
rect 13636 15444 13688 15496
rect 14832 15487 14884 15496
rect 14832 15453 14841 15487
rect 14841 15453 14875 15487
rect 14875 15453 14884 15487
rect 14832 15444 14884 15453
rect 8944 15308 8996 15360
rect 9312 15308 9364 15360
rect 9772 15351 9824 15360
rect 9772 15317 9781 15351
rect 9781 15317 9815 15351
rect 9815 15317 9824 15351
rect 9772 15308 9824 15317
rect 9864 15351 9916 15360
rect 9864 15317 9873 15351
rect 9873 15317 9907 15351
rect 9907 15317 9916 15351
rect 9864 15308 9916 15317
rect 10324 15308 10376 15360
rect 10692 15308 10744 15360
rect 10876 15351 10928 15360
rect 10876 15317 10885 15351
rect 10885 15317 10919 15351
rect 10919 15317 10928 15351
rect 10876 15308 10928 15317
rect 11152 15308 11204 15360
rect 12072 15351 12124 15360
rect 12072 15317 12081 15351
rect 12081 15317 12115 15351
rect 12115 15317 12124 15351
rect 12072 15308 12124 15317
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 14004 15308 14056 15360
rect 14372 15308 14424 15360
rect 15016 15376 15068 15428
rect 19616 15580 19668 15632
rect 21640 15648 21692 15700
rect 22928 15580 22980 15632
rect 23664 15648 23716 15700
rect 24584 15648 24636 15700
rect 29736 15580 29788 15632
rect 19432 15512 19484 15564
rect 20628 15512 20680 15564
rect 20996 15512 21048 15564
rect 17040 15487 17092 15496
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 20168 15444 20220 15496
rect 17316 15419 17368 15428
rect 17316 15385 17325 15419
rect 17325 15385 17359 15419
rect 17359 15385 17368 15419
rect 17316 15376 17368 15385
rect 17776 15376 17828 15428
rect 19156 15376 19208 15428
rect 15476 15351 15528 15360
rect 15476 15317 15485 15351
rect 15485 15317 15519 15351
rect 15519 15317 15528 15351
rect 15476 15308 15528 15317
rect 16120 15308 16172 15360
rect 16396 15308 16448 15360
rect 17408 15308 17460 15360
rect 19340 15308 19392 15360
rect 22560 15444 22612 15496
rect 21916 15308 21968 15360
rect 25780 15555 25832 15564
rect 25780 15521 25789 15555
rect 25789 15521 25823 15555
rect 25823 15521 25832 15555
rect 25780 15512 25832 15521
rect 23296 15444 23348 15496
rect 26148 15444 26200 15496
rect 37280 15444 37332 15496
rect 23940 15419 23992 15428
rect 23940 15385 23949 15419
rect 23949 15385 23983 15419
rect 23983 15385 23992 15419
rect 23940 15376 23992 15385
rect 23388 15308 23440 15360
rect 25228 15351 25280 15360
rect 25228 15317 25237 15351
rect 25237 15317 25271 15351
rect 25271 15317 25280 15351
rect 25228 15308 25280 15317
rect 25596 15351 25648 15360
rect 25596 15317 25605 15351
rect 25605 15317 25639 15351
rect 25639 15317 25648 15351
rect 25596 15308 25648 15317
rect 26148 15308 26200 15360
rect 26884 15308 26936 15360
rect 44824 15308 44876 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 3516 15147 3568 15156
rect 3516 15113 3525 15147
rect 3525 15113 3559 15147
rect 3559 15113 3568 15147
rect 3516 15104 3568 15113
rect 3792 15104 3844 15156
rect 4620 15104 4672 15156
rect 4712 15104 4764 15156
rect 7932 15104 7984 15156
rect 11244 15104 11296 15156
rect 4436 15036 4488 15088
rect 5816 15036 5868 15088
rect 2872 14968 2924 15020
rect 3516 14968 3568 15020
rect 4160 15011 4212 15020
rect 4160 14977 4169 15011
rect 4169 14977 4203 15011
rect 4203 14977 4212 15011
rect 4160 14968 4212 14977
rect 5540 14968 5592 15020
rect 6460 14968 6512 15020
rect 6736 14968 6788 15020
rect 8852 15036 8904 15088
rect 10048 15036 10100 15088
rect 10508 15036 10560 15088
rect 10600 15036 10652 15088
rect 15476 15104 15528 15156
rect 18420 15147 18472 15156
rect 18420 15113 18429 15147
rect 18429 15113 18463 15147
rect 18463 15113 18472 15147
rect 18420 15104 18472 15113
rect 22100 15104 22152 15156
rect 22560 15104 22612 15156
rect 24952 15104 25004 15156
rect 27068 15147 27120 15156
rect 27068 15113 27077 15147
rect 27077 15113 27111 15147
rect 27111 15113 27120 15147
rect 27068 15104 27120 15113
rect 1308 14900 1360 14952
rect 4804 14900 4856 14952
rect 4896 14900 4948 14952
rect 5908 14900 5960 14952
rect 8668 14968 8720 15020
rect 9312 14968 9364 15020
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14968 12032 14977
rect 9588 14900 9640 14952
rect 9680 14900 9732 14952
rect 10784 14900 10836 14952
rect 4436 14764 4488 14816
rect 6920 14764 6972 14816
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 7932 14832 7984 14884
rect 10324 14832 10376 14884
rect 10600 14832 10652 14884
rect 8208 14764 8260 14816
rect 8484 14764 8536 14816
rect 8852 14764 8904 14816
rect 9404 14764 9456 14816
rect 11796 14900 11848 14952
rect 14924 15036 14976 15088
rect 15384 15036 15436 15088
rect 16396 15036 16448 15088
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 13268 14900 13320 14952
rect 12624 14832 12676 14884
rect 13728 14832 13780 14884
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 17776 14968 17828 15020
rect 19432 14968 19484 15020
rect 20260 15036 20312 15088
rect 20720 15036 20772 15088
rect 20996 15036 21048 15088
rect 22192 15036 22244 15088
rect 14280 14900 14332 14952
rect 14924 14900 14976 14952
rect 15568 14900 15620 14952
rect 19616 14900 19668 14952
rect 20260 14900 20312 14952
rect 20628 14968 20680 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 23388 14968 23440 15020
rect 23940 14968 23992 15020
rect 11152 14764 11204 14816
rect 13820 14764 13872 14816
rect 16948 14832 17000 14884
rect 17500 14832 17552 14884
rect 16304 14807 16356 14816
rect 16304 14773 16313 14807
rect 16313 14773 16347 14807
rect 16347 14773 16356 14807
rect 16304 14764 16356 14773
rect 19248 14764 19300 14816
rect 19340 14807 19392 14816
rect 19340 14773 19349 14807
rect 19349 14773 19383 14807
rect 19383 14773 19392 14807
rect 19340 14764 19392 14773
rect 19984 14832 20036 14884
rect 21916 14832 21968 14884
rect 23388 14832 23440 14884
rect 20996 14764 21048 14816
rect 23848 14764 23900 14816
rect 25320 14764 25372 14816
rect 26608 14807 26660 14816
rect 26608 14773 26617 14807
rect 26617 14773 26651 14807
rect 26651 14773 26660 14807
rect 26608 14764 26660 14773
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 4160 14492 4212 14544
rect 5356 14492 5408 14544
rect 1308 14424 1360 14476
rect 4436 14424 4488 14476
rect 5724 14560 5776 14612
rect 6828 14492 6880 14544
rect 8208 14492 8260 14544
rect 9496 14560 9548 14612
rect 9588 14560 9640 14612
rect 13360 14560 13412 14612
rect 13728 14603 13780 14612
rect 13728 14569 13737 14603
rect 13737 14569 13771 14603
rect 13771 14569 13780 14603
rect 13728 14560 13780 14569
rect 14740 14560 14792 14612
rect 14924 14560 14976 14612
rect 35072 14560 35124 14612
rect 11796 14492 11848 14544
rect 13820 14492 13872 14544
rect 14188 14492 14240 14544
rect 14280 14492 14332 14544
rect 6460 14424 6512 14476
rect 6736 14424 6788 14476
rect 6920 14424 6972 14476
rect 7012 14424 7064 14476
rect 7748 14424 7800 14476
rect 9680 14424 9732 14476
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 10416 14424 10468 14476
rect 10600 14424 10652 14476
rect 10692 14424 10744 14476
rect 10968 14424 11020 14476
rect 13452 14424 13504 14476
rect 13728 14424 13780 14476
rect 21548 14492 21600 14544
rect 23572 14492 23624 14544
rect 25780 14492 25832 14544
rect 26884 14535 26936 14544
rect 16304 14424 16356 14476
rect 17132 14424 17184 14476
rect 17224 14424 17276 14476
rect 20076 14424 20128 14476
rect 20168 14424 20220 14476
rect 22008 14424 22060 14476
rect 23940 14424 23992 14476
rect 2596 14288 2648 14340
rect 2872 14220 2924 14272
rect 4528 14220 4580 14272
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 5172 14356 5224 14408
rect 6828 14356 6880 14408
rect 9404 14356 9456 14408
rect 10876 14356 10928 14408
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 18144 14356 18196 14408
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 20720 14356 20772 14408
rect 21824 14356 21876 14408
rect 25596 14424 25648 14476
rect 26884 14501 26893 14535
rect 26893 14501 26927 14535
rect 26927 14501 26936 14535
rect 26884 14492 26936 14501
rect 26608 14424 26660 14476
rect 6000 14288 6052 14340
rect 8484 14288 8536 14340
rect 6736 14220 6788 14272
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 8668 14220 8720 14272
rect 9312 14220 9364 14272
rect 9680 14220 9732 14272
rect 10600 14263 10652 14272
rect 10600 14229 10609 14263
rect 10609 14229 10643 14263
rect 10643 14229 10652 14263
rect 10600 14220 10652 14229
rect 11520 14288 11572 14340
rect 11152 14220 11204 14272
rect 14004 14288 14056 14340
rect 15384 14288 15436 14340
rect 12624 14220 12676 14272
rect 12900 14220 12952 14272
rect 16856 14288 16908 14340
rect 17408 14288 17460 14340
rect 17776 14288 17828 14340
rect 21916 14288 21968 14340
rect 23848 14288 23900 14340
rect 16396 14263 16448 14272
rect 16396 14229 16405 14263
rect 16405 14229 16439 14263
rect 16439 14229 16448 14263
rect 16396 14220 16448 14229
rect 16580 14220 16632 14272
rect 18512 14220 18564 14272
rect 20536 14263 20588 14272
rect 20536 14229 20545 14263
rect 20545 14229 20579 14263
rect 20579 14229 20588 14263
rect 20536 14220 20588 14229
rect 21548 14220 21600 14272
rect 22008 14220 22060 14272
rect 22836 14220 22888 14272
rect 23388 14220 23440 14272
rect 25136 14288 25188 14340
rect 26148 14331 26200 14340
rect 26148 14297 26157 14331
rect 26157 14297 26191 14331
rect 26191 14297 26200 14331
rect 26148 14288 26200 14297
rect 24584 14263 24636 14272
rect 24584 14229 24593 14263
rect 24593 14229 24627 14263
rect 24627 14229 24636 14263
rect 24584 14220 24636 14229
rect 25320 14220 25372 14272
rect 25780 14263 25832 14272
rect 25780 14229 25789 14263
rect 25789 14229 25823 14263
rect 25823 14229 25832 14263
rect 25780 14220 25832 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 3424 14059 3476 14068
rect 3424 14025 3433 14059
rect 3433 14025 3467 14059
rect 3467 14025 3476 14059
rect 3424 14016 3476 14025
rect 4712 14016 4764 14068
rect 6368 14016 6420 14068
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 2596 13948 2648 14000
rect 4620 13948 4672 14000
rect 6460 13991 6512 14000
rect 6460 13957 6469 13991
rect 6469 13957 6503 13991
rect 6503 13957 6512 13991
rect 6460 13948 6512 13957
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 7472 14016 7524 14068
rect 7748 14016 7800 14068
rect 9220 14016 9272 14068
rect 8576 13991 8628 14000
rect 8576 13957 8585 13991
rect 8585 13957 8619 13991
rect 8619 13957 8628 13991
rect 8576 13948 8628 13957
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 1308 13812 1360 13864
rect 4896 13880 4948 13932
rect 5264 13880 5316 13932
rect 10324 13948 10376 14000
rect 11152 14016 11204 14068
rect 11244 13948 11296 14000
rect 11612 13991 11664 14000
rect 11612 13957 11621 13991
rect 11621 13957 11655 13991
rect 11655 13957 11664 13991
rect 11612 13948 11664 13957
rect 11796 13948 11848 14000
rect 12256 14016 12308 14068
rect 12624 14016 12676 14068
rect 13084 14016 13136 14068
rect 12164 13948 12216 14000
rect 4712 13855 4764 13864
rect 4712 13821 4721 13855
rect 4721 13821 4755 13855
rect 4755 13821 4764 13855
rect 4712 13812 4764 13821
rect 5908 13855 5960 13864
rect 5908 13821 5917 13855
rect 5917 13821 5951 13855
rect 5951 13821 5960 13855
rect 5908 13812 5960 13821
rect 6736 13812 6788 13864
rect 5724 13744 5776 13796
rect 6092 13744 6144 13796
rect 6368 13744 6420 13796
rect 7012 13812 7064 13864
rect 8484 13812 8536 13864
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 10784 13812 10836 13864
rect 14188 14016 14240 14068
rect 14832 14059 14884 14068
rect 14832 14025 14841 14059
rect 14841 14025 14875 14059
rect 14875 14025 14884 14059
rect 14832 14016 14884 14025
rect 16580 14016 16632 14068
rect 17316 14016 17368 14068
rect 16672 13948 16724 14000
rect 13544 13923 13596 13932
rect 13544 13889 13553 13923
rect 13553 13889 13587 13923
rect 13587 13889 13596 13923
rect 13544 13880 13596 13889
rect 5264 13719 5316 13728
rect 5264 13685 5273 13719
rect 5273 13685 5307 13719
rect 5307 13685 5316 13719
rect 5264 13676 5316 13685
rect 5356 13676 5408 13728
rect 9036 13676 9088 13728
rect 12348 13744 12400 13796
rect 13084 13812 13136 13864
rect 15752 13880 15804 13932
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 16948 13880 17000 13932
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 14464 13812 14516 13864
rect 14924 13855 14976 13864
rect 14924 13821 14933 13855
rect 14933 13821 14967 13855
rect 14967 13821 14976 13855
rect 14924 13812 14976 13821
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 17868 13948 17920 14000
rect 20076 14059 20128 14068
rect 20076 14025 20085 14059
rect 20085 14025 20119 14059
rect 20119 14025 20128 14059
rect 20076 14016 20128 14025
rect 20352 14016 20404 14068
rect 20996 14016 21048 14068
rect 21180 14016 21232 14068
rect 25780 14016 25832 14068
rect 20904 13948 20956 14000
rect 21824 13991 21876 14000
rect 21824 13957 21833 13991
rect 21833 13957 21867 13991
rect 21867 13957 21876 13991
rect 21824 13948 21876 13957
rect 10692 13676 10744 13728
rect 14832 13744 14884 13796
rect 15200 13744 15252 13796
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 17776 13812 17828 13864
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 22376 13880 22428 13932
rect 22560 13923 22612 13932
rect 22560 13889 22569 13923
rect 22569 13889 22603 13923
rect 22603 13889 22612 13923
rect 24584 13948 24636 14000
rect 25136 13948 25188 14000
rect 22560 13880 22612 13889
rect 18788 13812 18840 13864
rect 20352 13812 20404 13864
rect 19248 13744 19300 13796
rect 14464 13676 14516 13728
rect 16672 13719 16724 13728
rect 16672 13685 16681 13719
rect 16681 13685 16715 13719
rect 16715 13685 16724 13719
rect 16672 13676 16724 13685
rect 17408 13719 17460 13728
rect 17408 13685 17438 13719
rect 17438 13685 17460 13719
rect 17408 13676 17460 13685
rect 20628 13744 20680 13796
rect 20996 13812 21048 13864
rect 24124 13880 24176 13932
rect 25320 13880 25372 13932
rect 22744 13744 22796 13796
rect 23756 13744 23808 13796
rect 24032 13855 24084 13864
rect 24032 13821 24041 13855
rect 24041 13821 24075 13855
rect 24075 13821 24084 13855
rect 24032 13812 24084 13821
rect 25136 13812 25188 13864
rect 22836 13676 22888 13728
rect 24584 13719 24636 13728
rect 24584 13685 24593 13719
rect 24593 13685 24627 13719
rect 24627 13685 24636 13719
rect 24584 13676 24636 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 4252 13472 4304 13524
rect 4620 13472 4672 13524
rect 7380 13472 7432 13524
rect 5448 13404 5500 13456
rect 9036 13472 9088 13524
rect 14372 13472 14424 13524
rect 15016 13472 15068 13524
rect 17408 13472 17460 13524
rect 20352 13472 20404 13524
rect 2044 13379 2096 13388
rect 2044 13345 2053 13379
rect 2053 13345 2087 13379
rect 2087 13345 2096 13379
rect 2044 13336 2096 13345
rect 5172 13336 5224 13388
rect 1768 13311 1820 13320
rect 1768 13277 1777 13311
rect 1777 13277 1811 13311
rect 1811 13277 1820 13311
rect 1768 13268 1820 13277
rect 5540 13268 5592 13320
rect 5816 13268 5868 13320
rect 4436 13243 4488 13252
rect 4436 13209 4445 13243
rect 4445 13209 4479 13243
rect 4479 13209 4488 13243
rect 4436 13200 4488 13209
rect 4528 13200 4580 13252
rect 1860 13132 1912 13184
rect 3792 13132 3844 13184
rect 4712 13132 4764 13184
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 6184 13132 6236 13184
rect 10692 13404 10744 13456
rect 11520 13447 11572 13456
rect 11520 13413 11529 13447
rect 11529 13413 11563 13447
rect 11563 13413 11572 13447
rect 11520 13404 11572 13413
rect 7472 13336 7524 13388
rect 8484 13379 8536 13388
rect 8484 13345 8493 13379
rect 8493 13345 8527 13379
rect 8527 13345 8536 13379
rect 8484 13336 8536 13345
rect 9036 13336 9088 13388
rect 9404 13379 9456 13388
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 10876 13379 10928 13388
rect 10876 13345 10885 13379
rect 10885 13345 10919 13379
rect 10919 13345 10928 13379
rect 10876 13336 10928 13345
rect 11244 13336 11296 13388
rect 11796 13404 11848 13456
rect 13728 13447 13780 13456
rect 13728 13413 13737 13447
rect 13737 13413 13771 13447
rect 13771 13413 13780 13447
rect 13728 13404 13780 13413
rect 22192 13472 22244 13524
rect 22560 13515 22612 13524
rect 22560 13481 22569 13515
rect 22569 13481 22603 13515
rect 22603 13481 22612 13515
rect 22560 13472 22612 13481
rect 23296 13472 23348 13524
rect 23940 13515 23992 13524
rect 23940 13481 23949 13515
rect 23949 13481 23983 13515
rect 23983 13481 23992 13515
rect 23940 13472 23992 13481
rect 24124 13515 24176 13524
rect 24124 13481 24133 13515
rect 24133 13481 24167 13515
rect 24167 13481 24176 13515
rect 24124 13472 24176 13481
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 15200 13336 15252 13388
rect 16396 13336 16448 13388
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 17132 13379 17184 13388
rect 17132 13345 17141 13379
rect 17141 13345 17175 13379
rect 17175 13345 17184 13379
rect 17132 13336 17184 13345
rect 17500 13336 17552 13388
rect 20076 13336 20128 13388
rect 22192 13336 22244 13388
rect 22836 13404 22888 13456
rect 32496 13472 32548 13524
rect 23480 13379 23532 13388
rect 23480 13345 23489 13379
rect 23489 13345 23523 13379
rect 23523 13345 23532 13379
rect 23480 13336 23532 13345
rect 23756 13336 23808 13388
rect 24676 13336 24728 13388
rect 14004 13268 14056 13320
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 23020 13268 23072 13320
rect 7012 13243 7064 13252
rect 7012 13209 7021 13243
rect 7021 13209 7055 13243
rect 7055 13209 7064 13243
rect 7012 13200 7064 13209
rect 7104 13200 7156 13252
rect 9680 13200 9732 13252
rect 9772 13132 9824 13184
rect 11612 13132 11664 13184
rect 12348 13200 12400 13252
rect 13728 13200 13780 13252
rect 14096 13200 14148 13252
rect 14188 13200 14240 13252
rect 14832 13200 14884 13252
rect 15292 13200 15344 13252
rect 17408 13243 17460 13252
rect 13636 13132 13688 13184
rect 13820 13132 13872 13184
rect 17408 13209 17417 13243
rect 17417 13209 17451 13243
rect 17451 13209 17460 13243
rect 17408 13200 17460 13209
rect 17868 13200 17920 13252
rect 16212 13132 16264 13184
rect 18972 13200 19024 13252
rect 22376 13200 22428 13252
rect 21272 13132 21324 13184
rect 23112 13200 23164 13252
rect 23756 13200 23808 13252
rect 23940 13200 23992 13252
rect 27528 13200 27580 13252
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 3608 12971 3660 12980
rect 3608 12937 3617 12971
rect 3617 12937 3651 12971
rect 3651 12937 3660 12971
rect 3608 12928 3660 12937
rect 4528 12928 4580 12980
rect 5632 12928 5684 12980
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 6184 12928 6236 12980
rect 6828 12928 6880 12980
rect 7104 12928 7156 12980
rect 10600 12928 10652 12980
rect 12440 12928 12492 12980
rect 14556 12928 14608 12980
rect 15292 12928 15344 12980
rect 16672 12928 16724 12980
rect 16948 12928 17000 12980
rect 18788 12928 18840 12980
rect 21180 12928 21232 12980
rect 21272 12928 21324 12980
rect 22008 12928 22060 12980
rect 2872 12860 2924 12912
rect 3700 12860 3752 12912
rect 3976 12860 4028 12912
rect 4344 12860 4396 12912
rect 4436 12860 4488 12912
rect 1216 12792 1268 12844
rect 2320 12792 2372 12844
rect 2504 12792 2556 12844
rect 3884 12792 3936 12844
rect 5080 12792 5132 12844
rect 5448 12792 5500 12844
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 5356 12724 5408 12776
rect 2504 12656 2556 12708
rect 7288 12792 7340 12844
rect 9404 12792 9456 12844
rect 7472 12724 7524 12776
rect 8300 12767 8352 12776
rect 8300 12733 8309 12767
rect 8309 12733 8343 12767
rect 8343 12733 8352 12767
rect 8300 12724 8352 12733
rect 10324 12860 10376 12912
rect 13636 12860 13688 12912
rect 13820 12860 13872 12912
rect 14280 12860 14332 12912
rect 9956 12792 10008 12844
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 10140 12724 10192 12776
rect 13084 12792 13136 12844
rect 13452 12792 13504 12844
rect 14740 12792 14792 12844
rect 15108 12792 15160 12844
rect 18420 12860 18472 12912
rect 18880 12860 18932 12912
rect 17408 12792 17460 12844
rect 18052 12792 18104 12844
rect 22284 12860 22336 12912
rect 10508 12699 10560 12708
rect 10508 12665 10517 12699
rect 10517 12665 10551 12699
rect 10551 12665 10560 12699
rect 10508 12656 10560 12665
rect 12256 12656 12308 12708
rect 2228 12588 2280 12640
rect 2964 12631 3016 12640
rect 2964 12597 2973 12631
rect 2973 12597 3007 12631
rect 3007 12597 3016 12631
rect 2964 12588 3016 12597
rect 3516 12588 3568 12640
rect 4620 12588 4672 12640
rect 5448 12588 5500 12640
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 6920 12588 6972 12640
rect 7472 12588 7524 12640
rect 8024 12588 8076 12640
rect 9312 12588 9364 12640
rect 11428 12588 11480 12640
rect 12164 12588 12216 12640
rect 12900 12588 12952 12640
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 15200 12724 15252 12776
rect 15292 12724 15344 12776
rect 15108 12656 15160 12708
rect 15476 12656 15528 12708
rect 18420 12767 18472 12776
rect 18420 12733 18429 12767
rect 18429 12733 18463 12767
rect 18463 12733 18472 12767
rect 18420 12724 18472 12733
rect 20076 12724 20128 12776
rect 21456 12724 21508 12776
rect 22468 12724 22520 12776
rect 22744 12928 22796 12980
rect 23204 12928 23256 12980
rect 23480 12928 23532 12980
rect 23572 12860 23624 12912
rect 23848 12860 23900 12912
rect 23020 12835 23072 12844
rect 23020 12801 23029 12835
rect 23029 12801 23063 12835
rect 23063 12801 23072 12835
rect 23020 12792 23072 12801
rect 23848 12724 23900 12776
rect 18328 12588 18380 12640
rect 21732 12656 21784 12708
rect 24400 12656 24452 12708
rect 20904 12588 20956 12640
rect 22008 12588 22060 12640
rect 22284 12588 22336 12640
rect 23020 12588 23072 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 3332 12384 3384 12436
rect 3792 12384 3844 12436
rect 3976 12427 4028 12436
rect 3976 12393 3985 12427
rect 3985 12393 4019 12427
rect 4019 12393 4028 12427
rect 3976 12384 4028 12393
rect 4160 12316 4212 12368
rect 1492 12180 1544 12232
rect 3424 12248 3476 12300
rect 3976 12248 4028 12300
rect 7748 12384 7800 12436
rect 10876 12384 10928 12436
rect 12532 12384 12584 12436
rect 7012 12316 7064 12368
rect 5172 12248 5224 12300
rect 6092 12248 6144 12300
rect 6184 12248 6236 12300
rect 2964 12223 3016 12232
rect 2964 12189 2973 12223
rect 2973 12189 3007 12223
rect 3007 12189 3016 12223
rect 2964 12180 3016 12189
rect 4252 12180 4304 12232
rect 7472 12248 7524 12300
rect 13728 12316 13780 12368
rect 15292 12316 15344 12368
rect 15476 12316 15528 12368
rect 18052 12427 18104 12436
rect 18052 12393 18061 12427
rect 18061 12393 18095 12427
rect 18095 12393 18104 12427
rect 18052 12384 18104 12393
rect 18880 12427 18932 12436
rect 18880 12393 18889 12427
rect 18889 12393 18923 12427
rect 18923 12393 18932 12427
rect 18880 12384 18932 12393
rect 20720 12384 20772 12436
rect 21916 12384 21968 12436
rect 19432 12316 19484 12368
rect 25596 12384 25648 12436
rect 9312 12248 9364 12300
rect 12072 12248 12124 12300
rect 12256 12291 12308 12300
rect 12256 12257 12265 12291
rect 12265 12257 12299 12291
rect 12299 12257 12308 12291
rect 12256 12248 12308 12257
rect 12348 12291 12400 12300
rect 12348 12257 12357 12291
rect 12357 12257 12391 12291
rect 12391 12257 12400 12291
rect 12348 12248 12400 12257
rect 10416 12180 10468 12232
rect 3424 12044 3476 12096
rect 5724 12112 5776 12164
rect 6644 12112 6696 12164
rect 7748 12112 7800 12164
rect 8024 12112 8076 12164
rect 8392 12112 8444 12164
rect 8576 12112 8628 12164
rect 8668 12112 8720 12164
rect 9036 12112 9088 12164
rect 9128 12155 9180 12164
rect 9128 12121 9137 12155
rect 9137 12121 9171 12155
rect 9171 12121 9180 12155
rect 9128 12112 9180 12121
rect 9680 12112 9732 12164
rect 13176 12180 13228 12232
rect 11612 12112 11664 12164
rect 15200 12248 15252 12300
rect 16672 12248 16724 12300
rect 19616 12291 19668 12300
rect 19616 12257 19625 12291
rect 19625 12257 19659 12291
rect 19659 12257 19668 12291
rect 19616 12248 19668 12257
rect 20076 12291 20128 12300
rect 20076 12257 20085 12291
rect 20085 12257 20119 12291
rect 20119 12257 20128 12291
rect 20076 12248 20128 12257
rect 20812 12248 20864 12300
rect 21916 12248 21968 12300
rect 14464 12180 14516 12232
rect 22192 12180 22244 12232
rect 13728 12112 13780 12164
rect 14740 12155 14792 12164
rect 14740 12121 14749 12155
rect 14749 12121 14783 12155
rect 14783 12121 14792 12155
rect 14740 12112 14792 12121
rect 14832 12112 14884 12164
rect 16672 12112 16724 12164
rect 4344 12044 4396 12096
rect 6276 12044 6328 12096
rect 7104 12044 7156 12096
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 11060 12044 11112 12096
rect 13176 12044 13228 12096
rect 13912 12044 13964 12096
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 14188 12044 14240 12096
rect 16580 12044 16632 12096
rect 17868 12112 17920 12164
rect 18696 12112 18748 12164
rect 18880 12112 18932 12164
rect 20352 12155 20404 12164
rect 20352 12121 20361 12155
rect 20361 12121 20395 12155
rect 20395 12121 20404 12155
rect 20352 12112 20404 12121
rect 21824 12112 21876 12164
rect 23020 12112 23072 12164
rect 24032 12087 24084 12096
rect 24032 12053 24041 12087
rect 24041 12053 24075 12087
rect 24075 12053 24084 12087
rect 24032 12044 24084 12053
rect 24400 12087 24452 12096
rect 24400 12053 24409 12087
rect 24409 12053 24443 12087
rect 24443 12053 24452 12087
rect 24400 12044 24452 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 1768 11840 1820 11892
rect 1952 11840 2004 11892
rect 3608 11840 3660 11892
rect 5448 11840 5500 11892
rect 4252 11772 4304 11824
rect 2412 11747 2464 11756
rect 2412 11713 2421 11747
rect 2421 11713 2455 11747
rect 2455 11713 2464 11747
rect 2412 11704 2464 11713
rect 4436 11704 4488 11756
rect 5264 11704 5316 11756
rect 6828 11772 6880 11824
rect 6920 11704 6972 11756
rect 7748 11772 7800 11824
rect 8208 11772 8260 11824
rect 1952 11636 2004 11688
rect 5172 11636 5224 11688
rect 5908 11636 5960 11688
rect 6092 11636 6144 11688
rect 9128 11704 9180 11756
rect 10600 11840 10652 11892
rect 9864 11772 9916 11824
rect 10508 11772 10560 11824
rect 11612 11815 11664 11824
rect 11612 11781 11621 11815
rect 11621 11781 11655 11815
rect 11655 11781 11664 11815
rect 11612 11772 11664 11781
rect 11796 11772 11848 11824
rect 8392 11636 8444 11688
rect 9864 11636 9916 11688
rect 13820 11840 13872 11892
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 17316 11883 17368 11892
rect 17316 11849 17325 11883
rect 17325 11849 17359 11883
rect 17359 11849 17368 11883
rect 17316 11840 17368 11849
rect 17868 11840 17920 11892
rect 18328 11840 18380 11892
rect 15476 11772 15528 11824
rect 17132 11772 17184 11824
rect 15936 11747 15988 11756
rect 15936 11713 15945 11747
rect 15945 11713 15979 11747
rect 15979 11713 15988 11747
rect 15936 11704 15988 11713
rect 20904 11840 20956 11892
rect 21824 11772 21876 11824
rect 8668 11568 8720 11620
rect 10232 11568 10284 11620
rect 15016 11636 15068 11688
rect 17040 11636 17092 11688
rect 13176 11568 13228 11620
rect 14556 11568 14608 11620
rect 17592 11679 17644 11688
rect 17592 11645 17601 11679
rect 17601 11645 17635 11679
rect 17635 11645 17644 11679
rect 17592 11636 17644 11645
rect 18604 11679 18656 11688
rect 18604 11645 18613 11679
rect 18613 11645 18647 11679
rect 18647 11645 18656 11679
rect 18604 11636 18656 11645
rect 18696 11679 18748 11688
rect 18696 11645 18705 11679
rect 18705 11645 18739 11679
rect 18739 11645 18748 11679
rect 18696 11636 18748 11645
rect 19708 11679 19760 11688
rect 19708 11645 19717 11679
rect 19717 11645 19751 11679
rect 19751 11645 19760 11679
rect 19708 11636 19760 11645
rect 24032 11840 24084 11892
rect 22744 11772 22796 11824
rect 23112 11772 23164 11824
rect 22192 11636 22244 11688
rect 19616 11568 19668 11620
rect 23664 11636 23716 11688
rect 24400 11611 24452 11620
rect 5264 11500 5316 11552
rect 5724 11500 5776 11552
rect 8300 11500 8352 11552
rect 9404 11500 9456 11552
rect 9496 11500 9548 11552
rect 10324 11500 10376 11552
rect 11980 11543 12032 11552
rect 11980 11509 11989 11543
rect 11989 11509 12023 11543
rect 12023 11509 12032 11543
rect 11980 11500 12032 11509
rect 12072 11500 12124 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 18604 11500 18656 11552
rect 21456 11543 21508 11552
rect 21456 11509 21465 11543
rect 21465 11509 21499 11543
rect 21499 11509 21508 11543
rect 21456 11500 21508 11509
rect 21824 11500 21876 11552
rect 23112 11500 23164 11552
rect 24400 11577 24409 11611
rect 24409 11577 24443 11611
rect 24443 11577 24452 11611
rect 24400 11568 24452 11577
rect 23756 11500 23808 11552
rect 25136 11500 25188 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 3700 11296 3752 11348
rect 5724 11296 5776 11348
rect 10600 11296 10652 11348
rect 11244 11296 11296 11348
rect 11612 11296 11664 11348
rect 12348 11296 12400 11348
rect 13360 11296 13412 11348
rect 13452 11296 13504 11348
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 1584 11024 1636 11076
rect 3700 11092 3752 11144
rect 6828 11160 6880 11212
rect 8668 11228 8720 11280
rect 9404 11228 9456 11280
rect 7840 11160 7892 11212
rect 8484 11203 8536 11212
rect 8484 11169 8493 11203
rect 8493 11169 8527 11203
rect 8527 11169 8536 11203
rect 8484 11160 8536 11169
rect 9220 11160 9272 11212
rect 10876 11228 10928 11280
rect 14832 11296 14884 11348
rect 15108 11296 15160 11348
rect 18972 11296 19024 11348
rect 22836 11296 22888 11348
rect 31760 11296 31812 11348
rect 10784 11203 10836 11212
rect 10784 11169 10793 11203
rect 10793 11169 10827 11203
rect 10827 11169 10836 11203
rect 10784 11160 10836 11169
rect 13360 11160 13412 11212
rect 15016 11160 15068 11212
rect 18696 11160 18748 11212
rect 21824 11160 21876 11212
rect 27528 11160 27580 11212
rect 6644 11092 6696 11144
rect 1952 10956 2004 11008
rect 4988 11024 5040 11076
rect 5172 11024 5224 11076
rect 7196 11024 7248 11076
rect 8852 11092 8904 11144
rect 9772 11092 9824 11144
rect 9864 11092 9916 11144
rect 14464 11092 14516 11144
rect 16856 11092 16908 11144
rect 18880 11092 18932 11144
rect 8300 11024 8352 11076
rect 7104 10956 7156 11008
rect 9220 10956 9272 11008
rect 9404 11024 9456 11076
rect 12256 11024 12308 11076
rect 13820 10999 13872 11008
rect 13820 10965 13829 10999
rect 13829 10965 13863 10999
rect 13863 10965 13872 10999
rect 13820 10956 13872 10965
rect 14096 10956 14148 11008
rect 15016 11067 15068 11076
rect 15016 11033 15025 11067
rect 15025 11033 15059 11067
rect 15059 11033 15068 11067
rect 15016 11024 15068 11033
rect 15476 11024 15528 11076
rect 16488 11024 16540 11076
rect 15384 10956 15436 11008
rect 16580 10956 16632 11008
rect 17868 11024 17920 11076
rect 19708 11024 19760 11076
rect 21180 11067 21232 11076
rect 21180 11033 21189 11067
rect 21189 11033 21223 11067
rect 21223 11033 21232 11067
rect 21180 11024 21232 11033
rect 21824 11024 21876 11076
rect 27620 11024 27672 11076
rect 31300 11024 31352 11076
rect 47860 11024 47912 11076
rect 18420 10956 18472 11008
rect 21364 10956 21416 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 4436 10752 4488 10804
rect 4804 10727 4856 10736
rect 4804 10693 4813 10727
rect 4813 10693 4847 10727
rect 4847 10693 4856 10727
rect 4804 10684 4856 10693
rect 4896 10684 4948 10736
rect 1124 10480 1176 10532
rect 3700 10591 3752 10600
rect 3700 10557 3709 10591
rect 3709 10557 3743 10591
rect 3743 10557 3752 10591
rect 3700 10548 3752 10557
rect 4252 10548 4304 10600
rect 5356 10659 5408 10668
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 5356 10616 5408 10625
rect 8852 10616 8904 10668
rect 9956 10795 10008 10804
rect 9956 10761 9965 10795
rect 9965 10761 9999 10795
rect 9999 10761 10008 10795
rect 9956 10752 10008 10761
rect 11152 10752 11204 10804
rect 11888 10752 11940 10804
rect 9496 10727 9548 10736
rect 9496 10693 9505 10727
rect 9505 10693 9539 10727
rect 9539 10693 9548 10727
rect 9496 10684 9548 10693
rect 14740 10752 14792 10804
rect 16948 10752 17000 10804
rect 17040 10752 17092 10804
rect 12900 10684 12952 10736
rect 15752 10684 15804 10736
rect 13636 10616 13688 10668
rect 14832 10616 14884 10668
rect 4896 10480 4948 10532
rect 6736 10548 6788 10600
rect 1952 10412 2004 10464
rect 2412 10412 2464 10464
rect 7104 10480 7156 10532
rect 6736 10412 6788 10464
rect 8116 10548 8168 10600
rect 8208 10548 8260 10600
rect 10232 10548 10284 10600
rect 10968 10591 11020 10600
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 11244 10548 11296 10600
rect 10416 10480 10468 10532
rect 11888 10480 11940 10532
rect 11980 10480 12032 10532
rect 15200 10548 15252 10600
rect 14648 10480 14700 10532
rect 16120 10591 16172 10600
rect 16120 10557 16129 10591
rect 16129 10557 16163 10591
rect 16163 10557 16172 10591
rect 16120 10548 16172 10557
rect 16304 10548 16356 10600
rect 17868 10684 17920 10736
rect 17500 10659 17552 10668
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 21456 10752 21508 10804
rect 20260 10684 20312 10736
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 22836 10548 22888 10600
rect 7840 10412 7892 10464
rect 9864 10412 9916 10464
rect 11520 10412 11572 10464
rect 11796 10412 11848 10464
rect 15660 10412 15712 10464
rect 21364 10480 21416 10532
rect 20536 10412 20588 10464
rect 21824 10455 21876 10464
rect 21824 10421 21833 10455
rect 21833 10421 21867 10455
rect 21867 10421 21876 10455
rect 21824 10412 21876 10421
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 1216 10208 1268 10260
rect 2872 10208 2924 10260
rect 7748 10208 7800 10260
rect 8760 10208 8812 10260
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 10784 10208 10836 10260
rect 11060 10208 11112 10260
rect 11520 10208 11572 10260
rect 11980 10208 12032 10260
rect 12072 10208 12124 10260
rect 13636 10208 13688 10260
rect 3332 10140 3384 10192
rect 4160 10140 4212 10192
rect 4896 10140 4948 10192
rect 5908 10140 5960 10192
rect 6644 10140 6696 10192
rect 8116 10140 8168 10192
rect 10968 10140 11020 10192
rect 15844 10208 15896 10260
rect 16580 10251 16632 10260
rect 16580 10217 16589 10251
rect 16589 10217 16623 10251
rect 16623 10217 16632 10251
rect 16580 10208 16632 10217
rect 18880 10251 18932 10260
rect 18880 10217 18889 10251
rect 18889 10217 18923 10251
rect 18923 10217 18932 10251
rect 18880 10208 18932 10217
rect 20168 10208 20220 10260
rect 20260 10208 20312 10260
rect 21824 10208 21876 10260
rect 1400 10072 1452 10124
rect 2688 10004 2740 10056
rect 5632 10072 5684 10124
rect 6828 10115 6880 10124
rect 6828 10081 6837 10115
rect 6837 10081 6871 10115
rect 6871 10081 6880 10115
rect 6828 10072 6880 10081
rect 7840 10072 7892 10124
rect 8300 10072 8352 10124
rect 11888 10072 11940 10124
rect 11980 10072 12032 10124
rect 13820 10140 13872 10192
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 15200 10072 15252 10124
rect 16212 10072 16264 10124
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 4344 10004 4396 10056
rect 8852 10004 8904 10056
rect 9312 10004 9364 10056
rect 9496 10004 9548 10056
rect 11060 10004 11112 10056
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 14464 10004 14516 10056
rect 16856 10004 16908 10056
rect 19708 10072 19760 10124
rect 21824 10004 21876 10056
rect 23572 10004 23624 10056
rect 4160 9936 4212 9988
rect 6368 9936 6420 9988
rect 3700 9868 3752 9920
rect 5356 9911 5408 9920
rect 5356 9877 5365 9911
rect 5365 9877 5399 9911
rect 5399 9877 5408 9911
rect 5356 9868 5408 9877
rect 11428 9936 11480 9988
rect 11796 9936 11848 9988
rect 8484 9868 8536 9920
rect 8576 9868 8628 9920
rect 10784 9868 10836 9920
rect 11980 9936 12032 9988
rect 15476 9936 15528 9988
rect 17040 9936 17092 9988
rect 12164 9868 12216 9920
rect 15016 9868 15068 9920
rect 16580 9868 16632 9920
rect 17868 9936 17920 9988
rect 19248 9936 19300 9988
rect 20168 9936 20220 9988
rect 23388 9936 23440 9988
rect 21180 9911 21232 9920
rect 21180 9877 21189 9911
rect 21189 9877 21223 9911
rect 21223 9877 21232 9911
rect 21180 9868 21232 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 6644 9664 6696 9716
rect 6736 9664 6788 9716
rect 13636 9664 13688 9716
rect 13820 9707 13872 9716
rect 13820 9673 13829 9707
rect 13829 9673 13863 9707
rect 13863 9673 13872 9707
rect 13820 9664 13872 9673
rect 1492 9639 1544 9648
rect 1492 9605 1501 9639
rect 1501 9605 1535 9639
rect 1535 9605 1544 9639
rect 1492 9596 1544 9605
rect 1768 9596 1820 9648
rect 2596 9596 2648 9648
rect 3608 9596 3660 9648
rect 5448 9596 5500 9648
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 3332 9528 3384 9580
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 1492 9460 1544 9512
rect 8392 9596 8444 9648
rect 10600 9596 10652 9648
rect 11888 9596 11940 9648
rect 16212 9707 16264 9716
rect 16212 9673 16221 9707
rect 16221 9673 16255 9707
rect 16255 9673 16264 9707
rect 16212 9664 16264 9673
rect 16396 9596 16448 9648
rect 18420 9664 18472 9716
rect 18880 9664 18932 9716
rect 18512 9596 18564 9648
rect 24584 9596 24636 9648
rect 6644 9528 6696 9580
rect 7748 9528 7800 9580
rect 9496 9528 9548 9580
rect 9680 9528 9732 9580
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 7840 9460 7892 9512
rect 10232 9460 10284 9512
rect 10968 9503 11020 9512
rect 10968 9469 10977 9503
rect 10977 9469 11011 9503
rect 11011 9469 11020 9503
rect 10968 9460 11020 9469
rect 11244 9460 11296 9512
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 14740 9460 14792 9469
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 17500 9460 17552 9512
rect 23756 9528 23808 9580
rect 28448 9528 28500 9580
rect 21180 9460 21232 9512
rect 23388 9460 23440 9512
rect 3608 9435 3660 9444
rect 3608 9401 3617 9435
rect 3617 9401 3651 9435
rect 3651 9401 3660 9435
rect 3608 9392 3660 9401
rect 940 9324 992 9376
rect 6644 9392 6696 9444
rect 9496 9392 9548 9444
rect 10784 9392 10836 9444
rect 13360 9392 13412 9444
rect 5632 9324 5684 9376
rect 6000 9324 6052 9376
rect 8484 9324 8536 9376
rect 10324 9367 10376 9376
rect 10324 9333 10333 9367
rect 10333 9333 10367 9367
rect 10367 9333 10376 9367
rect 10324 9324 10376 9333
rect 12164 9324 12216 9376
rect 12532 9324 12584 9376
rect 12716 9324 12768 9376
rect 13728 9324 13780 9376
rect 18512 9392 18564 9444
rect 14188 9324 14240 9376
rect 16028 9324 16080 9376
rect 16120 9324 16172 9376
rect 19064 9435 19116 9444
rect 19064 9401 19073 9435
rect 19073 9401 19107 9435
rect 19107 9401 19116 9435
rect 19064 9392 19116 9401
rect 31300 9596 31352 9648
rect 20168 9324 20220 9376
rect 28448 9367 28500 9376
rect 28448 9333 28457 9367
rect 28457 9333 28491 9367
rect 28491 9333 28500 9367
rect 28448 9324 28500 9333
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 3424 9120 3476 9172
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 2964 9052 3016 9104
rect 3884 9052 3936 9104
rect 4528 8984 4580 9036
rect 4988 9120 5040 9172
rect 6644 9120 6696 9172
rect 7472 9120 7524 9172
rect 9680 9120 9732 9172
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 11060 9120 11112 9172
rect 11612 9120 11664 9172
rect 12532 9120 12584 9172
rect 14188 9120 14240 9172
rect 15936 9120 15988 9172
rect 17592 9120 17644 9172
rect 28448 9120 28500 9172
rect 36360 9120 36412 9172
rect 2872 8916 2924 8968
rect 3332 8959 3384 8968
rect 3332 8925 3341 8959
rect 3341 8925 3375 8959
rect 3375 8925 3384 8959
rect 3332 8916 3384 8925
rect 8944 9052 8996 9104
rect 6184 9027 6236 9036
rect 6184 8993 6193 9027
rect 6193 8993 6227 9027
rect 6227 8993 6236 9027
rect 6184 8984 6236 8993
rect 6828 8984 6880 9036
rect 3424 8848 3476 8900
rect 5540 8891 5592 8900
rect 5540 8857 5549 8891
rect 5549 8857 5583 8891
rect 5583 8857 5592 8891
rect 5540 8848 5592 8857
rect 7748 8916 7800 8968
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8484 9027 8536 9036
rect 8484 8993 8493 9027
rect 8493 8993 8527 9027
rect 8527 8993 8536 9027
rect 8484 8984 8536 8993
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 15016 9052 15068 9104
rect 15384 9095 15436 9104
rect 15384 9061 15393 9095
rect 15393 9061 15427 9095
rect 15427 9061 15436 9095
rect 15384 9052 15436 9061
rect 15844 9052 15896 9104
rect 10876 8984 10928 9036
rect 12256 8984 12308 9036
rect 13728 8984 13780 9036
rect 15752 8984 15804 9036
rect 16856 8984 16908 9036
rect 9128 8848 9180 8900
rect 10968 8848 11020 8900
rect 12808 8848 12860 8900
rect 5172 8780 5224 8832
rect 7012 8780 7064 8832
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 9496 8780 9548 8832
rect 9680 8780 9732 8832
rect 10692 8780 10744 8832
rect 12440 8780 12492 8832
rect 16212 8848 16264 8900
rect 17224 8780 17276 8832
rect 18512 8780 18564 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 2872 8576 2924 8628
rect 3700 8576 3752 8628
rect 3792 8576 3844 8628
rect 3516 8508 3568 8560
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 5908 8576 5960 8628
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 6644 8619 6696 8628
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 7748 8576 7800 8628
rect 8116 8576 8168 8628
rect 10048 8576 10100 8628
rect 10416 8576 10468 8628
rect 10508 8619 10560 8628
rect 10508 8585 10517 8619
rect 10517 8585 10551 8619
rect 10551 8585 10560 8619
rect 10508 8576 10560 8585
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 12164 8619 12216 8628
rect 12164 8585 12173 8619
rect 12173 8585 12207 8619
rect 12207 8585 12216 8619
rect 12164 8576 12216 8585
rect 12256 8576 12308 8628
rect 14832 8576 14884 8628
rect 6920 8508 6972 8560
rect 7564 8508 7616 8560
rect 10692 8508 10744 8560
rect 1676 8440 1728 8492
rect 2136 8440 2188 8492
rect 3332 8440 3384 8492
rect 4252 8440 4304 8492
rect 5172 8440 5224 8492
rect 3516 8372 3568 8424
rect 1032 8304 1084 8356
rect 8116 8372 8168 8424
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 11060 8440 11112 8492
rect 12624 8483 12676 8492
rect 12624 8449 12633 8483
rect 12633 8449 12667 8483
rect 12667 8449 12676 8483
rect 12624 8440 12676 8449
rect 16304 8576 16356 8628
rect 17224 8576 17276 8628
rect 32404 8576 32456 8628
rect 15844 8508 15896 8560
rect 16120 8508 16172 8560
rect 18420 8508 18472 8560
rect 20444 8440 20496 8492
rect 9496 8372 9548 8424
rect 10416 8372 10468 8424
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 12072 8372 12124 8424
rect 12348 8372 12400 8424
rect 12808 8372 12860 8424
rect 16120 8372 16172 8424
rect 20352 8372 20404 8424
rect 2964 8236 3016 8288
rect 7380 8236 7432 8288
rect 32864 8304 32916 8356
rect 8392 8236 8444 8288
rect 12440 8236 12492 8288
rect 16672 8236 16724 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 1492 8032 1544 8084
rect 3332 8075 3384 8084
rect 3332 8041 3341 8075
rect 3341 8041 3375 8075
rect 3375 8041 3384 8075
rect 3332 8032 3384 8041
rect 3516 8075 3568 8084
rect 3516 8041 3525 8075
rect 3525 8041 3559 8075
rect 3559 8041 3568 8075
rect 3516 8032 3568 8041
rect 3976 8032 4028 8084
rect 4160 8032 4212 8084
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 8300 8032 8352 8084
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 7196 7964 7248 8016
rect 2596 7896 2648 7948
rect 11704 8032 11756 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 17500 8032 17552 8084
rect 11336 7964 11388 8016
rect 2872 7828 2924 7880
rect 5356 7760 5408 7812
rect 10232 7939 10284 7948
rect 10232 7905 10241 7939
rect 10241 7905 10275 7939
rect 10275 7905 10284 7939
rect 10232 7896 10284 7905
rect 5632 7828 5684 7880
rect 15200 8007 15252 8016
rect 15200 7973 15209 8007
rect 15209 7973 15243 8007
rect 15243 7973 15252 8007
rect 15200 7964 15252 7973
rect 7564 7760 7616 7812
rect 12072 7828 12124 7880
rect 19248 7896 19300 7948
rect 12440 7760 12492 7812
rect 13636 7760 13688 7812
rect 12808 7692 12860 7744
rect 13360 7735 13412 7744
rect 13360 7701 13369 7735
rect 13369 7701 13403 7735
rect 13403 7701 13412 7735
rect 13360 7692 13412 7701
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 22836 7692 22888 7744
rect 23388 7692 23440 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 1952 7488 2004 7540
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 2044 7352 2096 7404
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 10968 7488 11020 7540
rect 13360 7488 13412 7540
rect 23940 7531 23992 7540
rect 23940 7497 23949 7531
rect 23949 7497 23983 7531
rect 23983 7497 23992 7531
rect 23940 7488 23992 7497
rect 27620 7488 27672 7540
rect 2964 7420 3016 7472
rect 8576 7420 8628 7472
rect 9220 7420 9272 7472
rect 2596 7352 2648 7404
rect 3608 7352 3660 7404
rect 3700 7395 3752 7404
rect 3700 7361 3709 7395
rect 3709 7361 3743 7395
rect 3743 7361 3752 7395
rect 3700 7352 3752 7361
rect 7656 7352 7708 7404
rect 5264 7284 5316 7336
rect 10324 7284 10376 7336
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 23572 7352 23624 7404
rect 22468 7327 22520 7336
rect 22468 7293 22477 7327
rect 22477 7293 22511 7327
rect 22511 7293 22520 7327
rect 22468 7284 22520 7293
rect 1308 7216 1360 7268
rect 3700 7216 3752 7268
rect 15660 7216 15712 7268
rect 2964 7148 3016 7200
rect 5724 7148 5776 7200
rect 14004 7148 14056 7200
rect 17500 7148 17552 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 3424 6987 3476 6996
rect 3424 6953 3433 6987
rect 3433 6953 3467 6987
rect 3467 6953 3476 6987
rect 3424 6944 3476 6953
rect 23940 6944 23992 6996
rect 2780 6876 2832 6928
rect 1308 6808 1360 6860
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 2596 6740 2648 6792
rect 3976 6851 4028 6860
rect 3976 6817 3985 6851
rect 3985 6817 4019 6851
rect 4019 6817 4028 6851
rect 3976 6808 4028 6817
rect 10508 6808 10560 6860
rect 19340 6808 19392 6860
rect 20720 6808 20772 6860
rect 23756 6851 23808 6860
rect 3608 6740 3660 6792
rect 21732 6740 21784 6792
rect 23756 6817 23765 6851
rect 23765 6817 23799 6851
rect 23799 6817 23808 6851
rect 23756 6808 23808 6817
rect 7288 6672 7340 6724
rect 2320 6604 2372 6656
rect 9772 6604 9824 6656
rect 23388 6647 23440 6656
rect 23388 6613 23397 6647
rect 23397 6613 23431 6647
rect 23431 6613 23440 6647
rect 23388 6604 23440 6613
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 4436 6400 4488 6452
rect 22836 6443 22888 6452
rect 22836 6409 22845 6443
rect 22845 6409 22879 6443
rect 22879 6409 22888 6443
rect 22836 6400 22888 6409
rect 1768 6332 1820 6384
rect 3976 6332 4028 6384
rect 2872 6264 2924 6316
rect 1308 6196 1360 6248
rect 11428 6196 11480 6248
rect 22744 6060 22796 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 1308 5856 1360 5908
rect 22468 5856 22520 5908
rect 7748 5788 7800 5840
rect 12624 5788 12676 5840
rect 21732 5831 21784 5840
rect 21732 5797 21741 5831
rect 21741 5797 21775 5831
rect 21775 5797 21784 5831
rect 21732 5788 21784 5797
rect 6552 5720 6604 5772
rect 14004 5720 14056 5772
rect 16856 5720 16908 5772
rect 1308 5652 1360 5704
rect 12624 5652 12676 5704
rect 17040 5516 17092 5568
rect 18512 5652 18564 5704
rect 20904 5695 20956 5704
rect 20904 5661 20913 5695
rect 20913 5661 20947 5695
rect 20947 5661 20956 5695
rect 22744 5720 22796 5772
rect 28724 5720 28776 5772
rect 28908 5720 28960 5772
rect 20904 5652 20956 5661
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 22192 5584 22244 5636
rect 23388 5584 23440 5636
rect 25504 5584 25556 5636
rect 21364 5559 21416 5568
rect 21364 5525 21373 5559
rect 21373 5525 21407 5559
rect 21407 5525 21416 5559
rect 21364 5516 21416 5525
rect 27160 5627 27212 5636
rect 27160 5593 27169 5627
rect 27169 5593 27203 5627
rect 27203 5593 27212 5627
rect 27160 5584 27212 5593
rect 27620 5516 27672 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 27160 5312 27212 5364
rect 28540 5244 28592 5296
rect 1308 5176 1360 5228
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 17500 5219 17552 5228
rect 17500 5185 17509 5219
rect 17509 5185 17543 5219
rect 17543 5185 17552 5219
rect 17500 5176 17552 5185
rect 9036 5108 9088 5160
rect 15476 5108 15528 5160
rect 21364 5176 21416 5228
rect 22192 5219 22244 5228
rect 22192 5185 22210 5219
rect 22210 5185 22244 5219
rect 22192 5176 22244 5185
rect 17684 5151 17736 5160
rect 17684 5117 17693 5151
rect 17693 5117 17727 5151
rect 17727 5117 17736 5151
rect 17684 5108 17736 5117
rect 28816 5151 28868 5160
rect 28816 5117 28825 5151
rect 28825 5117 28859 5151
rect 28859 5117 28868 5151
rect 28816 5108 28868 5117
rect 41420 5108 41472 5160
rect 33508 5040 33560 5092
rect 1860 4972 1912 5024
rect 17868 4972 17920 5024
rect 20536 4972 20588 5024
rect 25964 4972 26016 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 7564 4768 7616 4820
rect 17408 4768 17460 4820
rect 1308 4632 1360 4684
rect 10784 4632 10836 4684
rect 2872 4564 2924 4616
rect 20904 4768 20956 4820
rect 28816 4768 28868 4820
rect 27804 4632 27856 4684
rect 17684 4428 17736 4480
rect 25964 4539 26016 4548
rect 25964 4505 25973 4539
rect 25973 4505 26007 4539
rect 26007 4505 26016 4539
rect 25964 4496 26016 4505
rect 26424 4496 26476 4548
rect 27528 4496 27580 4548
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 1308 4224 1360 4276
rect 1400 4088 1452 4140
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 4160 4088 4212 4140
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 9680 3952 9732 4004
rect 3332 3884 3384 3936
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 10600 3680 10652 3732
rect 12072 3723 12124 3732
rect 12072 3689 12081 3723
rect 12081 3689 12115 3723
rect 12115 3689 12124 3723
rect 12072 3680 12124 3689
rect 13452 3612 13504 3664
rect 28908 3612 28960 3664
rect 44088 3612 44140 3664
rect 1308 3476 1360 3528
rect 27528 3544 27580 3596
rect 46756 3544 46808 3596
rect 2504 3476 2556 3528
rect 2872 3476 2924 3528
rect 4068 3476 4120 3528
rect 12072 3476 12124 3528
rect 27620 3476 27672 3528
rect 49424 3476 49476 3528
rect 20720 3408 20772 3460
rect 38752 3408 38804 3460
rect 11612 3383 11664 3392
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 9772 3136 9824 3188
rect 10416 3068 10468 3120
rect 12624 3111 12676 3120
rect 12624 3077 12633 3111
rect 12633 3077 12667 3111
rect 12667 3077 12676 3111
rect 12624 3068 12676 3077
rect 15476 3068 15528 3120
rect 17684 3068 17736 3120
rect 1308 2932 1360 2984
rect 2780 3000 2832 3052
rect 3332 3000 3384 3052
rect 2412 2932 2464 2984
rect 7840 3000 7892 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17868 3000 17920 3052
rect 20536 3043 20588 3052
rect 20536 3009 20545 3043
rect 20545 3009 20579 3043
rect 20579 3009 20588 3043
rect 20536 3000 20588 3009
rect 17408 2932 17460 2984
rect 8300 2796 8352 2848
rect 12440 2864 12492 2916
rect 17500 2796 17552 2848
rect 20076 2796 20128 2848
rect 22008 2796 22060 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 7748 2592 7800 2644
rect 25504 2635 25556 2644
rect 25504 2601 25513 2635
rect 25513 2601 25547 2635
rect 25547 2601 25556 2635
rect 25504 2592 25556 2601
rect 27804 2592 27856 2644
rect 28724 2592 28776 2644
rect 33508 2635 33560 2644
rect 33508 2601 33517 2635
rect 33517 2601 33551 2635
rect 33551 2601 33560 2635
rect 33508 2592 33560 2601
rect 2780 2524 2832 2576
rect 1216 2456 1268 2508
rect 4068 2456 4120 2508
rect 11612 2524 11664 2576
rect 6736 2456 6788 2508
rect 9404 2456 9456 2508
rect 12072 2456 12124 2508
rect 14740 2456 14792 2508
rect 17408 2456 17460 2508
rect 20168 2456 20220 2508
rect 22744 2456 22796 2508
rect 36360 2499 36412 2508
rect 36360 2465 36369 2499
rect 36369 2465 36403 2499
rect 36403 2465 36412 2499
rect 36360 2456 36412 2465
rect 1308 2320 1360 2372
rect 8300 2388 8352 2440
rect 9772 2388 9824 2440
rect 12440 2388 12492 2440
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 22008 2388 22060 2440
rect 25412 2388 25464 2440
rect 28356 2431 28408 2440
rect 28356 2397 28365 2431
rect 28365 2397 28399 2431
rect 28399 2397 28408 2431
rect 28356 2388 28408 2397
rect 30748 2388 30800 2440
rect 33416 2388 33468 2440
rect 36084 2431 36136 2440
rect 36084 2397 36093 2431
rect 36093 2397 36127 2431
rect 36127 2397 36136 2431
rect 36084 2388 36136 2397
rect 4896 2252 4948 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
<< metal2 >>
rect 2226 26200 2282 27000
rect 2870 26200 2926 27000
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26330 4858 27000
rect 4802 26302 5120 26330
rect 4802 26200 4858 26302
rect 1492 24336 1544 24342
rect 1492 24278 1544 24284
rect 1216 23588 1268 23594
rect 1216 23530 1268 23536
rect 1032 22772 1084 22778
rect 1032 22714 1084 22720
rect 1044 22094 1072 22714
rect 1124 22568 1176 22574
rect 1124 22510 1176 22516
rect 952 22066 1072 22094
rect 952 9382 980 22066
rect 1136 18086 1164 22510
rect 1124 18080 1176 18086
rect 1124 18022 1176 18028
rect 1228 17898 1256 23530
rect 1308 22092 1360 22098
rect 1504 22094 1532 24278
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 1768 23520 1820 23526
rect 2148 23497 2176 23666
rect 1768 23462 1820 23468
rect 2134 23488 2190 23497
rect 1504 22066 1624 22094
rect 1308 22034 1360 22040
rect 1320 20777 1348 22034
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1044 17870 1256 17898
rect 940 9376 992 9382
rect 940 9318 992 9324
rect 1044 8362 1072 17870
rect 1124 17740 1176 17746
rect 1124 17682 1176 17688
rect 1136 10538 1164 17682
rect 1216 17604 1268 17610
rect 1216 17546 1268 17552
rect 1228 17105 1256 17546
rect 1308 17128 1360 17134
rect 1214 17096 1270 17105
rect 1308 17070 1360 17076
rect 1214 17031 1270 17040
rect 1320 16697 1348 17070
rect 1306 16688 1362 16697
rect 1306 16623 1362 16632
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15881 1348 15982
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15473 1348 15506
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1306 15056 1362 15065
rect 1306 14991 1362 15000
rect 1320 14958 1348 14991
rect 1308 14952 1360 14958
rect 1308 14894 1360 14900
rect 1306 14648 1362 14657
rect 1306 14583 1362 14592
rect 1320 14482 1348 14583
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 1306 14240 1362 14249
rect 1306 14175 1362 14184
rect 1320 13870 1348 14175
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 1214 13424 1270 13433
rect 1214 13359 1270 13368
rect 1228 12850 1256 13359
rect 1216 12844 1268 12850
rect 1216 12786 1268 12792
rect 1124 10532 1176 10538
rect 1124 10474 1176 10480
rect 1228 10266 1256 12786
rect 1492 12232 1544 12238
rect 1306 12200 1362 12209
rect 1362 12180 1492 12186
rect 1362 12174 1544 12180
rect 1362 12158 1532 12174
rect 1306 12135 1362 12144
rect 1398 11792 1454 11801
rect 1398 11727 1454 11736
rect 1216 10260 1268 10266
rect 1216 10202 1268 10208
rect 1412 10130 1440 11727
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1504 9654 1532 12158
rect 1596 11082 1624 22066
rect 1674 21856 1730 21865
rect 1674 21791 1730 21800
rect 1688 11234 1716 21791
rect 1780 20466 1808 23462
rect 2134 23423 2190 23432
rect 1860 23316 1912 23322
rect 1860 23258 1912 23264
rect 1872 22642 1900 23258
rect 1952 22704 2004 22710
rect 1952 22646 2004 22652
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 1964 22030 1992 22646
rect 2134 22400 2190 22409
rect 2134 22335 2190 22344
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 2044 21480 2096 21486
rect 2044 21422 2096 21428
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1872 17814 1900 20878
rect 2056 19961 2084 21422
rect 2148 21010 2176 22335
rect 2240 22166 2268 26200
rect 2778 24440 2834 24449
rect 2778 24375 2834 24384
rect 2412 24200 2464 24206
rect 2412 24142 2464 24148
rect 2228 22160 2280 22166
rect 2228 22102 2280 22108
rect 2136 21004 2188 21010
rect 2136 20946 2188 20952
rect 2042 19952 2098 19961
rect 2042 19887 2098 19896
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 2056 17513 2084 18158
rect 2226 17776 2282 17785
rect 2226 17711 2282 17720
rect 2042 17504 2098 17513
rect 2042 17439 2098 17448
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1780 16794 1808 17138
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 2136 16720 2188 16726
rect 2136 16662 2188 16668
rect 1766 13968 1822 13977
rect 1766 13903 1768 13912
rect 1820 13903 1822 13912
rect 1768 13874 1820 13880
rect 1780 13818 1808 13874
rect 2042 13832 2098 13841
rect 1780 13790 1992 13818
rect 1768 13320 1820 13326
rect 1766 13288 1768 13297
rect 1820 13288 1822 13297
rect 1766 13223 1822 13232
rect 1780 11898 1808 13223
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1688 11206 1808 11234
rect 1780 11150 1808 11206
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1032 8356 1084 8362
rect 1032 8298 1084 8304
rect 1504 8090 1532 9454
rect 1596 9042 1624 9687
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1688 8498 1716 10911
rect 1780 9654 1808 11086
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1872 9042 1900 13126
rect 1964 11898 1992 13790
rect 2042 13767 2098 13776
rect 2056 13394 2084 13767
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2042 12608 2098 12617
rect 2042 12543 2098 12552
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 11014 1992 11630
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1964 10470 1992 10950
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1766 8936 1822 8945
rect 1766 8871 1822 8880
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 1320 7274 1348 7647
rect 1308 7268 1360 7274
rect 1308 7210 1360 7216
rect 1308 6860 1360 6866
rect 1308 6802 1360 6808
rect 1320 6497 1348 6802
rect 1780 6798 1808 8871
rect 1964 7546 1992 10406
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 2056 7410 2084 12543
rect 2148 8498 2176 16662
rect 2240 12730 2268 17711
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 2332 12850 2360 16594
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2240 12702 2360 12730
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2240 9586 2268 12582
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2226 7848 2282 7857
rect 2226 7783 2282 7792
rect 2240 7546 2268 7783
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1306 6488 1362 6497
rect 1306 6423 1362 6432
rect 1780 6390 1808 6734
rect 2332 6662 2360 12702
rect 2424 11762 2452 24142
rect 2792 24138 2820 24375
rect 2780 24132 2832 24138
rect 2780 24074 2832 24080
rect 2688 23724 2740 23730
rect 2688 23666 2740 23672
rect 2596 22432 2648 22438
rect 2596 22374 2648 22380
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2516 12850 2544 21490
rect 2608 14346 2636 22374
rect 2596 14340 2648 14346
rect 2596 14282 2648 14288
rect 2596 14000 2648 14006
rect 2596 13942 2648 13948
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 1768 6384 1820 6390
rect 1768 6326 1820 6332
rect 1308 6248 1360 6254
rect 1308 6190 1360 6196
rect 1320 6089 1348 6190
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 1320 5914 1348 6015
rect 1308 5908 1360 5914
rect 1308 5850 1360 5856
rect 1308 5704 1360 5710
rect 1306 5672 1308 5681
rect 1360 5672 1362 5681
rect 1306 5607 1362 5616
rect 1306 5264 1362 5273
rect 1306 5199 1308 5208
rect 1360 5199 1362 5208
rect 1308 5170 1360 5176
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1306 4856 1362 4865
rect 1306 4791 1362 4800
rect 1320 4690 1348 4791
rect 1308 4684 1360 4690
rect 1308 4626 1360 4632
rect 1320 4282 1348 4626
rect 1308 4276 1360 4282
rect 1308 4218 1360 4224
rect 1872 4146 1900 4966
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1320 3233 1348 3470
rect 1306 3224 1362 3233
rect 1306 3159 1362 3168
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 1320 2825 1348 2926
rect 1306 2816 1362 2825
rect 1306 2751 1362 2760
rect 1216 2508 1268 2514
rect 1216 2450 1268 2456
rect 1228 2417 1256 2450
rect 1214 2408 1270 2417
rect 1214 2343 1270 2352
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 1320 2009 1348 2314
rect 1306 2000 1362 2009
rect 1306 1935 1362 1944
rect 1412 800 1440 4082
rect 2424 2990 2452 10406
rect 2516 3534 2544 12650
rect 2608 9654 2636 13942
rect 2700 10062 2728 23666
rect 2884 23186 2912 26200
rect 3054 24848 3110 24857
rect 3054 24783 3110 24792
rect 3068 24682 3096 24783
rect 3056 24676 3108 24682
rect 3056 24618 3108 24624
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2872 23180 2924 23186
rect 2872 23122 2924 23128
rect 3436 23118 3464 24550
rect 3528 24274 3556 26200
rect 3790 25664 3846 25673
rect 3790 25599 3846 25608
rect 3698 25256 3754 25265
rect 3698 25191 3754 25200
rect 3712 25090 3740 25191
rect 3700 25084 3752 25090
rect 3700 25026 3752 25032
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3516 24064 3568 24070
rect 3516 24006 3568 24012
rect 3700 24064 3752 24070
rect 3700 24006 3752 24012
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3528 23050 3556 24006
rect 3712 23866 3740 24006
rect 3700 23860 3752 23866
rect 3700 23802 3752 23808
rect 3698 23216 3754 23225
rect 3698 23151 3754 23160
rect 3608 23112 3660 23118
rect 3606 23080 3608 23089
rect 3660 23080 3662 23089
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 3516 23044 3568 23050
rect 3606 23015 3662 23024
rect 3516 22986 3568 22992
rect 2792 22234 2820 22986
rect 3528 22658 3556 22986
rect 3344 22630 3556 22658
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 2780 22228 2832 22234
rect 2780 22170 2832 22176
rect 2778 21176 2834 21185
rect 2884 21162 2912 22510
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2964 22228 3016 22234
rect 2964 22170 3016 22176
rect 2976 21593 3004 22170
rect 2962 21584 3018 21593
rect 2962 21519 3018 21528
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2834 21134 2912 21162
rect 2778 21111 2834 21120
rect 3344 21078 3372 22630
rect 3516 22568 3568 22574
rect 3516 22510 3568 22516
rect 3332 21072 3384 21078
rect 3332 21014 3384 21020
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2792 19553 2820 20810
rect 2872 20392 2924 20398
rect 2872 20334 2924 20340
rect 2778 19544 2834 19553
rect 2884 19530 2912 20334
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3344 20058 3372 21014
rect 3528 20992 3556 22510
rect 3608 21888 3660 21894
rect 3608 21830 3660 21836
rect 3620 21457 3648 21830
rect 3606 21448 3662 21457
rect 3606 21383 3662 21392
rect 3528 20964 3648 20992
rect 3516 20868 3568 20874
rect 3516 20810 3568 20816
rect 3424 20460 3476 20466
rect 3424 20402 3476 20408
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 2884 19502 3004 19530
rect 2778 19479 2834 19488
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2792 17921 2820 18634
rect 2884 18329 2912 19314
rect 2976 19281 3004 19502
rect 2962 19272 3018 19281
rect 2962 19207 3018 19216
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3344 18737 3372 19858
rect 3330 18728 3386 18737
rect 3056 18692 3108 18698
rect 3330 18663 3386 18672
rect 3056 18634 3108 18640
rect 2870 18320 2926 18329
rect 2870 18255 2926 18264
rect 3068 18068 3096 18634
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 2884 18040 3096 18068
rect 2778 17912 2834 17921
rect 2778 17847 2834 17856
rect 2780 15428 2832 15434
rect 2780 15370 2832 15376
rect 2792 10713 2820 15370
rect 2884 15026 2912 18040
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3344 16998 3372 18566
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 3344 16658 3372 16934
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3436 16266 3464 20402
rect 3528 17134 3556 20810
rect 3620 19553 3648 20964
rect 3712 19718 3740 23151
rect 3804 22250 3832 25599
rect 4066 24032 4122 24041
rect 4066 23967 4122 23976
rect 3884 23724 3936 23730
rect 3884 23666 3936 23672
rect 3896 23633 3924 23666
rect 3882 23624 3938 23633
rect 3882 23559 3938 23568
rect 4080 22386 4108 23967
rect 4172 23798 4200 26200
rect 4802 24712 4858 24721
rect 4802 24647 4858 24656
rect 4252 24200 4304 24206
rect 4250 24168 4252 24177
rect 4304 24168 4306 24177
rect 4250 24103 4306 24112
rect 4436 24132 4488 24138
rect 4436 24074 4488 24080
rect 4160 23792 4212 23798
rect 4160 23734 4212 23740
rect 4344 23180 4396 23186
rect 4344 23122 4396 23128
rect 4252 23112 4304 23118
rect 4252 23054 4304 23060
rect 4160 22976 4212 22982
rect 4160 22918 4212 22924
rect 4172 22545 4200 22918
rect 4264 22642 4292 23054
rect 4252 22636 4304 22642
rect 4252 22578 4304 22584
rect 4158 22536 4214 22545
rect 4158 22471 4214 22480
rect 4080 22358 4200 22386
rect 3804 22222 3924 22250
rect 3792 22160 3844 22166
rect 3792 22102 3844 22108
rect 3700 19712 3752 19718
rect 3700 19654 3752 19660
rect 3606 19544 3662 19553
rect 3606 19479 3662 19488
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3514 16824 3570 16833
rect 3514 16759 3570 16768
rect 3528 16726 3556 16759
rect 3516 16720 3568 16726
rect 3516 16662 3568 16668
rect 3344 16238 3464 16266
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2884 13410 2912 14214
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2884 13382 3004 13410
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2778 10704 2834 10713
rect 2778 10639 2834 10648
rect 2778 10568 2834 10577
rect 2778 10503 2834 10512
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2792 9466 2820 10503
rect 2884 10266 2912 12854
rect 2976 12646 3004 13382
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 3344 12442 3372 16238
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3436 14074 3464 15438
rect 3528 15162 3556 16050
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3422 13016 3478 13025
rect 3422 12951 3478 12960
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 2962 12336 3018 12345
rect 2962 12271 3018 12280
rect 3330 12336 3386 12345
rect 3436 12306 3464 12951
rect 3528 12866 3556 14962
rect 3620 12986 3648 19314
rect 3804 18222 3832 22102
rect 3896 20534 3924 22222
rect 4172 22094 4200 22358
rect 4172 22066 4292 22094
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3988 21729 4016 21966
rect 3974 21720 4030 21729
rect 3974 21655 4030 21664
rect 4264 21162 4292 22066
rect 4356 21622 4384 23122
rect 4448 22094 4476 24074
rect 4816 23730 4844 24647
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4528 22976 4580 22982
rect 4526 22944 4528 22953
rect 4580 22944 4582 22953
rect 4526 22879 4582 22888
rect 4448 22066 4568 22094
rect 4344 21616 4396 21622
rect 4344 21558 4396 21564
rect 4264 21134 4384 21162
rect 4250 21040 4306 21049
rect 4160 21004 4212 21010
rect 4250 20975 4252 20984
rect 4160 20946 4212 20952
rect 4304 20975 4306 20984
rect 4252 20946 4304 20952
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 4066 20904 4122 20913
rect 3884 20528 3936 20534
rect 3884 20470 3936 20476
rect 3884 20392 3936 20398
rect 3882 20360 3884 20369
rect 3936 20360 3938 20369
rect 3882 20295 3938 20304
rect 3884 19780 3936 19786
rect 3884 19722 3936 19728
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3790 17776 3846 17785
rect 3790 17711 3846 17720
rect 3804 17678 3832 17711
rect 3792 17672 3844 17678
rect 3792 17614 3844 17620
rect 3896 17490 3924 19722
rect 3988 18057 4016 20878
rect 4066 20839 4122 20848
rect 4080 19854 4108 20839
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 4172 19446 4200 20946
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 4160 19440 4212 19446
rect 4160 19382 4212 19388
rect 4066 19136 4122 19145
rect 4066 19071 4122 19080
rect 4080 18698 4108 19071
rect 4068 18692 4120 18698
rect 4068 18634 4120 18640
rect 3974 18048 4030 18057
rect 3974 17983 4030 17992
rect 4160 17672 4212 17678
rect 4066 17640 4122 17649
rect 4160 17614 4212 17620
rect 4066 17575 4068 17584
rect 4120 17575 4122 17584
rect 4068 17546 4120 17552
rect 3896 17462 4016 17490
rect 3988 17338 4016 17462
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 4066 17096 4122 17105
rect 4066 17031 4122 17040
rect 4080 16726 4108 17031
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3988 16250 4016 16526
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3712 12918 3740 16050
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3792 15360 3844 15366
rect 3790 15328 3792 15337
rect 3844 15328 3846 15337
rect 3790 15263 3846 15272
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3804 13190 3832 15098
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3700 12912 3752 12918
rect 3528 12838 3648 12866
rect 3700 12854 3752 12860
rect 3896 12850 3924 15506
rect 4172 15026 4200 17614
rect 4264 16182 4292 20470
rect 4356 17270 4384 21134
rect 4434 18864 4490 18873
rect 4434 18799 4490 18808
rect 4448 18766 4476 18799
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4344 17264 4396 17270
rect 4344 17206 4396 17212
rect 4434 17232 4490 17241
rect 4434 17167 4490 17176
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3330 12271 3386 12280
rect 3424 12300 3476 12306
rect 2976 12238 3004 12271
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 3344 10198 3372 12271
rect 3424 12242 3476 12248
rect 3528 12186 3556 12582
rect 3620 12288 3648 12838
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3620 12260 3740 12288
rect 3436 12158 3556 12186
rect 3606 12200 3662 12209
rect 3436 12102 3464 12158
rect 3606 12135 3662 12144
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11354 3464 12038
rect 3620 11898 3648 12135
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3712 11354 3740 12260
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3514 11248 3570 11257
rect 3514 11183 3570 11192
rect 3698 11248 3754 11257
rect 3698 11183 3754 11192
rect 3332 10192 3384 10198
rect 2870 10160 2926 10169
rect 3332 10134 3384 10140
rect 3422 10160 3478 10169
rect 2870 10095 2926 10104
rect 3422 10095 3478 10104
rect 2608 9438 2820 9466
rect 2608 7954 2636 9438
rect 2778 9344 2834 9353
rect 2778 9279 2834 9288
rect 2792 8242 2820 9279
rect 2884 8974 2912 10095
rect 3436 10062 3464 10095
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8634 2912 8910
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2870 8528 2926 8537
rect 2870 8463 2926 8472
rect 2700 8214 2820 8242
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 2700 7426 2728 8214
rect 2778 8120 2834 8129
rect 2778 8055 2834 8064
rect 2608 7410 2728 7426
rect 2596 7404 2728 7410
rect 2648 7398 2728 7404
rect 2596 7346 2648 7352
rect 2792 7154 2820 8055
rect 2884 7886 2912 8463
rect 2976 8294 3004 9046
rect 3344 8974 3372 9522
rect 3436 9178 3464 9998
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3332 8968 3384 8974
rect 3330 8936 3332 8945
rect 3384 8936 3386 8945
rect 3330 8871 3386 8880
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 3344 8090 3372 8434
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2870 7304 2926 7313
rect 2870 7239 2926 7248
rect 2700 7126 2820 7154
rect 2596 6792 2648 6798
rect 2700 6746 2728 7126
rect 2780 6928 2832 6934
rect 2780 6870 2832 6876
rect 2792 6746 2820 6870
rect 2648 6740 2820 6746
rect 2596 6734 2820 6740
rect 2608 6718 2820 6734
rect 2884 6322 2912 7239
rect 2976 7206 3004 7414
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3436 7002 3464 8842
rect 3528 8566 3556 11183
rect 3712 11150 3740 11183
rect 3700 11144 3752 11150
rect 3620 11092 3700 11098
rect 3620 11086 3752 11092
rect 3620 11070 3740 11086
rect 3620 9654 3648 11070
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3712 10441 3740 10542
rect 3698 10432 3754 10441
rect 3698 10367 3754 10376
rect 3698 10160 3754 10169
rect 3698 10095 3754 10104
rect 3712 9926 3740 10095
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3608 9648 3660 9654
rect 3608 9590 3660 9596
rect 3606 9480 3662 9489
rect 3606 9415 3608 9424
rect 3660 9415 3662 9424
rect 3608 9386 3660 9392
rect 3712 8634 3740 9862
rect 3804 8634 3832 12378
rect 3896 9110 3924 12786
rect 3988 12442 4016 12854
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4172 12374 4200 14486
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4264 12764 4292 13466
rect 4356 12918 4384 15302
rect 4448 15094 4476 17167
rect 4540 16658 4568 22066
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4632 22001 4660 22034
rect 4618 21992 4674 22001
rect 4618 21927 4674 21936
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4632 17678 4660 18702
rect 4724 18680 4752 23122
rect 4986 22808 5042 22817
rect 4986 22743 5042 22752
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 4816 22234 4844 22578
rect 4804 22228 4856 22234
rect 4804 22170 4856 22176
rect 4896 21412 4948 21418
rect 4896 21354 4948 21360
rect 4804 19780 4856 19786
rect 4804 19722 4856 19728
rect 4816 19174 4844 19722
rect 4908 19514 4936 21354
rect 5000 20466 5028 22743
rect 5092 22574 5120 26302
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26330 7434 27000
rect 8022 26330 8078 27000
rect 6932 26302 7434 26330
rect 5460 23662 5488 26200
rect 5724 23860 5776 23866
rect 5724 23802 5776 23808
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5736 21622 5764 23802
rect 6104 23186 6132 26200
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6564 23526 6592 23666
rect 6552 23520 6604 23526
rect 6550 23488 6552 23497
rect 6604 23488 6606 23497
rect 6550 23423 6606 23432
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6000 22500 6052 22506
rect 6000 22442 6052 22448
rect 5724 21616 5776 21622
rect 5724 21558 5776 21564
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4804 18692 4856 18698
rect 4724 18652 4804 18680
rect 4804 18634 4856 18640
rect 4802 17912 4858 17921
rect 4802 17847 4858 17856
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4816 17610 4844 17847
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4632 15162 4660 17070
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4724 15162 4752 15982
rect 4908 15745 4936 17274
rect 4894 15736 4950 15745
rect 4894 15671 4950 15680
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4436 15088 4488 15094
rect 4436 15030 4488 15036
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4448 14482 4476 14758
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4448 13258 4476 14418
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4540 13988 4568 14214
rect 4724 14074 4752 14214
rect 4816 14113 4844 14894
rect 4802 14104 4858 14113
rect 4712 14068 4764 14074
rect 4802 14039 4858 14048
rect 4712 14010 4764 14016
rect 4620 14000 4672 14006
rect 4540 13960 4620 13988
rect 4620 13942 4672 13948
rect 4712 13864 4764 13870
rect 4632 13824 4712 13852
rect 4632 13530 4660 13824
rect 4816 13852 4844 14039
rect 4908 13938 4936 14894
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 4764 13824 4844 13852
rect 4712 13806 4764 13812
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4908 13410 4936 13874
rect 4816 13382 4936 13410
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 4528 13252 4580 13258
rect 4580 13212 4660 13240
rect 4528 13194 4580 13200
rect 4448 12918 4476 13194
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4264 12736 4476 12764
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4250 12336 4306 12345
rect 3976 12300 4028 12306
rect 4250 12271 4306 12280
rect 3976 12242 4028 12248
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3528 8090 3556 8366
rect 3988 8090 4016 12242
rect 4264 12238 4292 12271
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4264 11830 4292 12174
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4158 11384 4214 11393
rect 4158 11319 4214 11328
rect 4172 10198 4200 11319
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 4160 9988 4212 9994
rect 4160 9930 4212 9936
rect 4172 8090 4200 9930
rect 4264 9586 4292 10542
rect 4356 10062 4384 12038
rect 4448 11762 4476 12736
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4448 10810 4476 11698
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4434 10704 4490 10713
rect 4434 10639 4490 10648
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4250 8528 4306 8537
rect 4250 8463 4252 8472
rect 4304 8463 4306 8472
rect 4252 8434 4304 8440
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4264 8022 4292 8434
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3620 6905 3648 7346
rect 3712 7274 3740 7346
rect 3700 7268 3752 7274
rect 3700 7210 3752 7216
rect 3606 6896 3662 6905
rect 3606 6831 3662 6840
rect 3976 6860 4028 6866
rect 3620 6798 3648 6831
rect 3976 6802 4028 6808
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3988 6390 4016 6802
rect 4448 6458 4476 10639
rect 4540 9042 4568 12922
rect 4632 12646 4660 13212
rect 4712 13184 4764 13190
rect 4710 13152 4712 13161
rect 4764 13152 4766 13161
rect 4710 13087 4766 13096
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4618 11112 4674 11121
rect 4618 11047 4674 11056
rect 4632 9178 4660 11047
rect 4816 10742 4844 13382
rect 5000 13138 5028 19450
rect 4908 13110 5028 13138
rect 4908 10742 4936 13110
rect 5092 13002 5120 21422
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 5184 15570 5212 21286
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 5276 20058 5304 20742
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5276 19786 5304 19994
rect 5460 19922 5488 20878
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 5276 19417 5304 19722
rect 5262 19408 5318 19417
rect 5262 19343 5264 19352
rect 5316 19343 5318 19352
rect 5448 19346 5500 19352
rect 5264 19314 5316 19320
rect 5448 19288 5500 19294
rect 5356 19236 5408 19242
rect 5356 19178 5408 19184
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5184 13394 5212 14350
rect 5276 13938 5304 15846
rect 5368 14550 5396 19178
rect 5460 18698 5488 19288
rect 5448 18692 5500 18698
rect 5448 18634 5500 18640
rect 5460 17610 5488 18634
rect 5448 17604 5500 17610
rect 5448 17546 5500 17552
rect 5460 16504 5488 17546
rect 5552 16726 5580 21490
rect 5644 21321 5672 21490
rect 5630 21312 5686 21321
rect 5630 21247 5686 21256
rect 5632 20868 5684 20874
rect 5632 20810 5684 20816
rect 5644 20618 5672 20810
rect 5736 20777 5764 21558
rect 5908 20800 5960 20806
rect 5722 20768 5778 20777
rect 5908 20742 5960 20748
rect 5722 20703 5778 20712
rect 5644 20590 5764 20618
rect 5736 20534 5764 20590
rect 5724 20528 5776 20534
rect 5724 20470 5776 20476
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5816 20392 5868 20398
rect 5816 20334 5868 20340
rect 5632 20324 5684 20330
rect 5632 20266 5684 20272
rect 5644 18426 5672 20266
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5630 18320 5686 18329
rect 5630 18255 5632 18264
rect 5684 18255 5686 18264
rect 5632 18226 5684 18232
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 5630 16688 5686 16697
rect 5736 16658 5764 20334
rect 5828 17490 5856 20334
rect 5920 19310 5948 20742
rect 6012 19514 6040 22442
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 6104 20466 6132 21830
rect 6182 21584 6238 21593
rect 6182 21519 6238 21528
rect 6196 21350 6224 21519
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6196 20874 6224 21286
rect 6184 20868 6236 20874
rect 6184 20810 6236 20816
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 6090 20360 6146 20369
rect 6090 20295 6146 20304
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 5920 18358 5948 19246
rect 6104 18465 6132 20295
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6090 18456 6146 18465
rect 6090 18391 6146 18400
rect 5908 18352 5960 18358
rect 5908 18294 5960 18300
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 5908 18216 5960 18222
rect 5906 18184 5908 18193
rect 5960 18184 5962 18193
rect 5906 18119 5962 18128
rect 5828 17462 5948 17490
rect 5920 17134 5948 17462
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5630 16623 5686 16632
rect 5724 16652 5776 16658
rect 5460 16476 5580 16504
rect 5552 15026 5580 16476
rect 5644 16164 5672 16623
rect 5724 16594 5776 16600
rect 5908 16516 5960 16522
rect 5908 16458 5960 16464
rect 5724 16176 5776 16182
rect 5644 16136 5724 16164
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5000 12974 5120 13002
rect 5000 11082 5028 12974
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4908 10198 4936 10474
rect 4896 10192 4948 10198
rect 4896 10134 4948 10140
rect 5000 9178 5028 11018
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2884 3641 2912 4558
rect 4158 4448 4214 4457
rect 4158 4383 4214 4392
rect 4172 4146 4200 4383
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4066 4040 4122 4049
rect 4066 3975 4122 3984
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2870 3632 2926 3641
rect 2870 3567 2926 3576
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2792 2582 2820 2994
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 2884 1601 2912 3470
rect 3344 3058 3372 3878
rect 4080 3534 4108 3975
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 5092 2774 5120 12786
rect 5184 12306 5212 13330
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5276 11762 5304 13670
rect 5368 12782 5396 13670
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5460 12850 5488 13398
rect 5552 13326 5580 14962
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5644 12986 5672 16136
rect 5724 16118 5776 16124
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5828 15706 5856 16118
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5736 15065 5764 15302
rect 5816 15088 5868 15094
rect 5722 15056 5778 15065
rect 5816 15030 5868 15036
rect 5722 14991 5778 15000
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5736 13802 5764 14554
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5736 12986 5764 13738
rect 5828 13326 5856 15030
rect 5920 14958 5948 16458
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 6012 15638 6040 15982
rect 6000 15632 6052 15638
rect 6000 15574 6052 15580
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 6012 14346 6040 15574
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5460 11898 5488 12582
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5184 11082 5212 11630
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5354 11520 5410 11529
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5184 8634 5212 8774
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5184 8498 5212 8570
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5276 7342 5304 11494
rect 5354 11455 5410 11464
rect 5368 10674 5396 11455
rect 5446 11112 5502 11121
rect 5446 11047 5502 11056
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 7818 5396 9862
rect 5460 9654 5488 11047
rect 5644 10130 5672 12786
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5736 11558 5764 12106
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5736 11354 5764 11494
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5828 10690 5856 13262
rect 5920 13190 5948 13806
rect 6104 13802 6132 18226
rect 6196 17814 6224 18566
rect 6288 18154 6316 22918
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 6380 19334 6408 22374
rect 6656 22137 6684 24142
rect 6748 22710 6776 26200
rect 6932 24290 6960 26302
rect 7378 26200 7434 26302
rect 7852 26302 8078 26330
rect 7564 25084 7616 25090
rect 7564 25026 7616 25032
rect 7288 24676 7340 24682
rect 7288 24618 7340 24624
rect 6840 24274 6960 24290
rect 6828 24268 6960 24274
rect 6880 24262 6960 24268
rect 6828 24210 6880 24216
rect 7104 23860 7156 23866
rect 7104 23802 7156 23808
rect 7116 23633 7144 23802
rect 7102 23624 7158 23633
rect 7102 23559 7158 23568
rect 7196 23112 7248 23118
rect 7196 23054 7248 23060
rect 6736 22704 6788 22710
rect 6736 22646 6788 22652
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6642 22128 6698 22137
rect 6642 22063 6698 22072
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6472 20369 6500 21966
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6552 21480 6604 21486
rect 6552 21422 6604 21428
rect 6458 20360 6514 20369
rect 6458 20295 6514 20304
rect 6380 19306 6500 19334
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6380 18630 6408 19110
rect 6368 18624 6420 18630
rect 6368 18566 6420 18572
rect 6472 18193 6500 19306
rect 6458 18184 6514 18193
rect 6276 18148 6328 18154
rect 6458 18119 6514 18128
rect 6276 18090 6328 18096
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 6182 17504 6238 17513
rect 6182 17439 6238 17448
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6196 13682 6224 17439
rect 6368 17128 6420 17134
rect 6368 17070 6420 17076
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6012 13654 6224 13682
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5920 11694 5948 13126
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5736 10662 5856 10690
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5538 9616 5594 9625
rect 5538 9551 5594 9560
rect 5552 8906 5580 9551
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5644 7886 5672 9318
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5736 7206 5764 10662
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 5920 8634 5948 10134
rect 6012 9382 6040 13654
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6196 12986 6224 13126
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6196 12306 6224 12922
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6104 11694 6132 12242
rect 6288 12102 6316 16594
rect 6380 15978 6408 17070
rect 6472 16561 6500 17070
rect 6458 16552 6514 16561
rect 6458 16487 6514 16496
rect 6368 15972 6420 15978
rect 6368 15914 6420 15920
rect 6472 15473 6500 16487
rect 6564 16046 6592 21422
rect 6748 21078 6776 21558
rect 6736 21072 6788 21078
rect 6736 21014 6788 21020
rect 6734 19952 6790 19961
rect 6734 19887 6790 19896
rect 6748 19786 6776 19887
rect 6736 19780 6788 19786
rect 6736 19722 6788 19728
rect 6644 19236 6696 19242
rect 6644 19178 6696 19184
rect 6656 18290 6684 19178
rect 6734 18320 6790 18329
rect 6644 18284 6696 18290
rect 6734 18255 6736 18264
rect 6644 18226 6696 18232
rect 6788 18255 6790 18264
rect 6736 18226 6788 18232
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6458 15464 6514 15473
rect 6458 15399 6514 15408
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6380 14074 6408 15302
rect 6564 15042 6592 15982
rect 6656 15502 6684 15982
rect 6748 15570 6776 18022
rect 6840 17338 6868 22578
rect 7012 22568 7064 22574
rect 7012 22510 7064 22516
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6932 20777 6960 21966
rect 7024 21010 7052 22510
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7116 21146 7144 22374
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 7104 20868 7156 20874
rect 7104 20810 7156 20816
rect 6918 20768 6974 20777
rect 6918 20703 6974 20712
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6932 19378 6960 19654
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6564 15026 6776 15042
rect 6460 15020 6512 15026
rect 6564 15020 6788 15026
rect 6564 15014 6736 15020
rect 6460 14962 6512 14968
rect 6736 14962 6788 14968
rect 6472 14521 6500 14962
rect 6458 14512 6514 14521
rect 6748 14482 6776 14962
rect 6840 14550 6868 16390
rect 6932 16250 6960 18362
rect 7024 18290 7052 20538
rect 7116 20534 7144 20810
rect 7208 20777 7236 23054
rect 7194 20768 7250 20777
rect 7194 20703 7250 20712
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 7024 16250 7052 18090
rect 7116 17678 7144 20198
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7208 17814 7236 18634
rect 7300 18222 7328 24618
rect 7380 23656 7432 23662
rect 7380 23598 7432 23604
rect 7392 22098 7420 23598
rect 7380 22092 7432 22098
rect 7380 22034 7432 22040
rect 7576 21842 7604 25026
rect 7748 23724 7800 23730
rect 7748 23666 7800 23672
rect 7656 22092 7708 22098
rect 7656 22034 7708 22040
rect 7484 21814 7604 21842
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7392 21321 7420 21490
rect 7378 21312 7434 21321
rect 7378 21247 7434 21256
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7392 20466 7420 20946
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7286 17912 7342 17921
rect 7286 17847 7342 17856
rect 7196 17808 7248 17814
rect 7196 17750 7248 17756
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 7194 17640 7250 17649
rect 7194 17575 7196 17584
rect 7248 17575 7250 17584
rect 7196 17546 7248 17552
rect 7300 17354 7328 17847
rect 7392 17542 7420 20198
rect 7484 19938 7512 21814
rect 7668 21706 7696 22034
rect 7576 21678 7696 21706
rect 7576 21622 7604 21678
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7576 20058 7604 21558
rect 7656 21072 7708 21078
rect 7656 21014 7708 21020
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7484 19910 7604 19938
rect 7472 19780 7524 19786
rect 7472 19722 7524 19728
rect 7484 19417 7512 19722
rect 7576 19446 7604 19910
rect 7564 19440 7616 19446
rect 7470 19408 7526 19417
rect 7564 19382 7616 19388
rect 7470 19343 7526 19352
rect 7484 18680 7512 19343
rect 7564 18692 7616 18698
rect 7484 18652 7564 18680
rect 7564 18634 7616 18640
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7116 17326 7328 17354
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 7024 15638 7052 15846
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6932 14822 6960 15506
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 7024 14482 7052 15574
rect 7116 15570 7144 17326
rect 7288 17264 7340 17270
rect 7208 17224 7288 17252
rect 7208 15706 7236 17224
rect 7288 17206 7340 17212
rect 7392 16153 7420 17478
rect 7378 16144 7434 16153
rect 7288 16108 7340 16114
rect 7378 16079 7434 16088
rect 7288 16050 7340 16056
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7300 14906 7328 16050
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7392 15337 7420 15982
rect 7378 15328 7434 15337
rect 7378 15263 7434 15272
rect 7208 14878 7328 14906
rect 6458 14447 6460 14456
rect 6512 14447 6514 14456
rect 6736 14476 6788 14482
rect 6460 14418 6512 14424
rect 6736 14418 6788 14424
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 6828 14408 6880 14414
rect 6458 14376 6514 14385
rect 6828 14350 6880 14356
rect 6458 14311 6514 14320
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6472 14006 6500 14311
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6550 14104 6606 14113
rect 6550 14039 6552 14048
rect 6604 14039 6606 14048
rect 6552 14010 6604 14016
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6182 11928 6238 11937
rect 6182 11863 6238 11872
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6196 9042 6224 11863
rect 6380 9994 6408 13738
rect 6472 12434 6500 13942
rect 6748 13870 6776 14214
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6840 12986 6868 14350
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6932 12646 6960 14418
rect 7024 13870 7052 14418
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7024 13258 7052 13806
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6472 12406 6592 12434
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6366 9616 6422 9625
rect 6366 9551 6422 9560
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6380 8634 6408 9551
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 6564 5778 6592 12406
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6656 11150 6684 12106
rect 6840 11830 6868 12582
rect 7024 12374 7052 13194
rect 7116 12986 7144 13194
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7012 12368 7064 12374
rect 7208 12356 7236 14878
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 14074 7328 14758
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7392 13530 7420 15263
rect 7484 14074 7512 18294
rect 7564 17808 7616 17814
rect 7564 17750 7616 17756
rect 7576 17134 7604 17750
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7300 12753 7328 12786
rect 7484 12782 7512 13330
rect 7472 12776 7524 12782
rect 7286 12744 7342 12753
rect 7472 12718 7524 12724
rect 7286 12679 7342 12688
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7208 12328 7328 12356
rect 7012 12310 7064 12316
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6734 11656 6790 11665
rect 6734 11591 6790 11600
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6656 10198 6684 11086
rect 6748 10606 6776 11591
rect 6932 11529 6960 11698
rect 6918 11520 6974 11529
rect 6918 11455 6974 11464
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6656 9722 6684 10134
rect 6748 9722 6776 10406
rect 6840 10130 6868 11154
rect 7116 11014 7144 12038
rect 7194 11112 7250 11121
rect 7194 11047 7196 11056
rect 7248 11047 7250 11056
rect 7196 11018 7248 11024
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7010 10704 7066 10713
rect 7010 10639 7066 10648
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6918 10024 6974 10033
rect 6918 9959 6974 9968
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6656 9450 6684 9522
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6656 9178 6684 9386
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6840 9042 6868 9454
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6642 8664 6698 8673
rect 6642 8599 6644 8608
rect 6696 8599 6698 8608
rect 6644 8570 6696 8576
rect 6932 8566 6960 9959
rect 7024 8838 7052 10639
rect 7116 10538 7144 10950
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 7208 8022 7236 11018
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7300 6730 7328 12328
rect 7378 12336 7434 12345
rect 7484 12306 7512 12582
rect 7562 12472 7618 12481
rect 7562 12407 7618 12416
rect 7378 12271 7434 12280
rect 7472 12300 7524 12306
rect 7392 10441 7420 12271
rect 7472 12242 7524 12248
rect 7378 10432 7434 10441
rect 7378 10367 7434 10376
rect 7392 8294 7420 10367
rect 7576 10146 7604 12407
rect 7484 10118 7604 10146
rect 7484 9178 7512 10118
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7576 8090 7604 8502
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 7576 4826 7604 7754
rect 7668 7410 7696 21014
rect 7760 17338 7788 23666
rect 7852 23186 7880 26302
rect 8022 26200 8078 26302
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26330 10654 27000
rect 10598 26302 10732 26330
rect 10598 26200 10654 26302
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8484 23792 8536 23798
rect 8484 23734 8536 23740
rect 7932 23724 7984 23730
rect 7932 23666 7984 23672
rect 7944 23497 7972 23666
rect 7930 23488 7986 23497
rect 7930 23423 7986 23432
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7932 22704 7984 22710
rect 7932 22646 7984 22652
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7852 17814 7880 22578
rect 7944 22098 7972 22646
rect 8300 22636 8352 22642
rect 8300 22578 8352 22584
rect 7932 22092 7984 22098
rect 7932 22034 7984 22040
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8024 21616 8076 21622
rect 8022 21584 8024 21593
rect 8076 21584 8078 21593
rect 8022 21519 8078 21528
rect 8206 21584 8262 21593
rect 8206 21519 8262 21528
rect 8220 20942 8248 21519
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 8036 20058 8064 20198
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8312 19281 8340 22578
rect 8392 22092 8444 22098
rect 8496 22094 8524 23734
rect 8588 22420 8616 24142
rect 8680 22574 8708 26200
rect 9324 24290 9352 26200
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9692 24313 9720 24346
rect 9232 24274 9352 24290
rect 9220 24268 9352 24274
rect 9272 24262 9352 24268
rect 9678 24304 9734 24313
rect 9678 24239 9734 24248
rect 9220 24210 9272 24216
rect 8758 24168 8814 24177
rect 8758 24103 8814 24112
rect 8772 24070 8800 24103
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8588 22392 8708 22420
rect 8496 22066 8616 22094
rect 8392 22034 8444 22040
rect 8404 21622 8432 22034
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8392 21616 8444 21622
rect 8392 21558 8444 21564
rect 8404 20602 8432 21558
rect 8496 21486 8524 21830
rect 8484 21480 8536 21486
rect 8484 21422 8536 21428
rect 8588 20942 8616 22066
rect 8576 20936 8628 20942
rect 8576 20878 8628 20884
rect 8392 20596 8444 20602
rect 8392 20538 8444 20544
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8298 19272 8354 19281
rect 8404 19242 8432 20198
rect 8576 20052 8628 20058
rect 8576 19994 8628 20000
rect 8588 19961 8616 19994
rect 8574 19952 8630 19961
rect 8574 19887 8630 19896
rect 8680 19530 8708 22392
rect 8772 20534 8800 24006
rect 9968 23798 9996 26200
rect 10140 25696 10192 25702
rect 10140 25638 10192 25644
rect 10048 25560 10100 25566
rect 10048 25502 10100 25508
rect 9956 23792 10008 23798
rect 9956 23734 10008 23740
rect 9588 23520 9640 23526
rect 9588 23462 9640 23468
rect 9600 23168 9628 23462
rect 9508 23140 9720 23168
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 8852 23044 8904 23050
rect 8852 22986 8904 22992
rect 8864 21010 8892 22986
rect 8956 21350 8984 23054
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 9404 22976 9456 22982
rect 9508 22964 9536 23140
rect 9692 23050 9720 23140
rect 9588 23044 9640 23050
rect 9588 22986 9640 22992
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9456 22936 9536 22964
rect 9404 22918 9456 22924
rect 9048 22098 9076 22918
rect 9496 22160 9548 22166
rect 9496 22102 9548 22108
rect 9036 22092 9088 22098
rect 9036 22034 9088 22040
rect 9508 22001 9536 22102
rect 9310 21992 9366 22001
rect 9310 21927 9366 21936
rect 9494 21992 9550 22001
rect 9494 21927 9550 21936
rect 9324 21894 9352 21927
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8852 21004 8904 21010
rect 8852 20946 8904 20952
rect 8760 20528 8812 20534
rect 8760 20470 8812 20476
rect 8496 19502 8708 19530
rect 8298 19207 8354 19216
rect 8392 19236 8444 19242
rect 8392 19178 8444 19184
rect 8496 18986 8524 19502
rect 8772 19417 8800 20470
rect 8956 20398 8984 21286
rect 9036 20936 9088 20942
rect 9036 20878 9088 20884
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8956 19922 8984 20334
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 8758 19408 8814 19417
rect 8668 19372 8720 19378
rect 8758 19343 8814 19352
rect 8668 19314 8720 19320
rect 8574 19136 8630 19145
rect 8574 19071 8630 19080
rect 8312 18958 8524 18986
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 7944 18154 7972 18226
rect 7932 18148 7984 18154
rect 7932 18090 7984 18096
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7944 17626 7972 18090
rect 8022 17912 8078 17921
rect 8022 17847 8078 17856
rect 7852 17598 7972 17626
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7852 16538 7880 17598
rect 8036 17542 8064 17847
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8114 16824 8170 16833
rect 8114 16759 8170 16768
rect 7760 14482 7788 16526
rect 7852 16522 7972 16538
rect 7852 16516 7984 16522
rect 7852 16510 7932 16516
rect 7932 16458 7984 16464
rect 8128 16454 8156 16759
rect 8206 16552 8262 16561
rect 8312 16538 8340 18958
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8404 17882 8432 18226
rect 8496 18204 8524 18770
rect 8588 18698 8616 19071
rect 8576 18692 8628 18698
rect 8576 18634 8628 18640
rect 8576 18216 8628 18222
rect 8496 18176 8576 18204
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8404 16697 8432 17138
rect 8390 16688 8446 16697
rect 8390 16623 8446 16632
rect 8312 16510 8432 16538
rect 8206 16487 8208 16496
rect 8260 16487 8262 16496
rect 8208 16458 8260 16464
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 7852 14929 7880 16390
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7930 16144 7986 16153
rect 7930 16079 7986 16088
rect 7944 16046 7972 16079
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7944 15434 7972 15642
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8024 15496 8076 15502
rect 8220 15450 8248 15506
rect 8076 15444 8248 15450
rect 8024 15438 8248 15444
rect 7932 15428 7984 15434
rect 8036 15422 8248 15438
rect 7932 15370 7984 15376
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 7838 14920 7894 14929
rect 7944 14890 7972 15098
rect 8312 15042 8340 15574
rect 8220 15014 8340 15042
rect 7838 14855 7894 14864
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 8220 14822 8248 15014
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 8220 14278 8248 14486
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7760 12442 7788 14010
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7760 11830 7788 12106
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7852 11218 7880 14214
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8036 12170 8064 12582
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 8220 11098 8248 11766
rect 8312 11558 8340 12718
rect 8404 12170 8432 16510
rect 8496 16114 8524 18176
rect 8576 18158 8628 18164
rect 8576 17128 8628 17134
rect 8574 17096 8576 17105
rect 8628 17096 8630 17105
rect 8574 17031 8630 17040
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8496 15570 8524 15914
rect 8680 15706 8708 19314
rect 8944 18692 8996 18698
rect 8944 18634 8996 18640
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8772 17202 8800 18566
rect 8956 18426 8984 18634
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 8944 17876 8996 17882
rect 8944 17818 8996 17824
rect 8956 17678 8984 17818
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8942 17096 8998 17105
rect 8760 17060 8812 17066
rect 8942 17031 8998 17040
rect 8760 17002 8812 17008
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8588 15586 8616 15642
rect 8772 15586 8800 17002
rect 8850 16688 8906 16697
rect 8850 16623 8906 16632
rect 8484 15564 8536 15570
rect 8588 15558 8800 15586
rect 8484 15506 8536 15512
rect 8482 15464 8538 15473
rect 8482 15399 8538 15408
rect 8666 15464 8722 15473
rect 8666 15399 8722 15408
rect 8496 14822 8524 15399
rect 8574 15056 8630 15065
rect 8680 15026 8708 15399
rect 8864 15314 8892 16623
rect 8956 16522 8984 17031
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 8772 15286 8892 15314
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8574 14991 8630 15000
rect 8668 15020 8720 15026
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8482 14376 8538 14385
rect 8482 14311 8484 14320
rect 8536 14311 8538 14320
rect 8484 14282 8536 14288
rect 8588 14006 8616 14991
rect 8668 14962 8720 14968
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8496 13394 8524 13806
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 8392 11688 8444 11694
rect 8496 11676 8524 13330
rect 8680 12170 8708 14214
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8444 11648 8524 11676
rect 8392 11630 8444 11636
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8588 11370 8616 12106
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8404 11342 8616 11370
rect 8220 11082 8340 11098
rect 8220 11076 8352 11082
rect 8220 11070 8300 11076
rect 8300 11018 8352 11024
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7760 9586 7788 10202
rect 7852 10130 7880 10406
rect 8128 10198 8156 10542
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7852 9518 7880 10066
rect 8220 10010 8248 10542
rect 8312 10130 8340 11018
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8220 9982 8340 10010
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8312 9636 8340 9982
rect 8404 9654 8432 11342
rect 8680 11286 8708 11562
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8496 9926 8524 11154
rect 8772 10266 8800 15286
rect 8852 15088 8904 15094
rect 8852 15030 8904 15036
rect 8864 14929 8892 15030
rect 8850 14920 8906 14929
rect 8850 14855 8906 14864
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8864 11150 8892 14758
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8864 10062 8892 10610
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8220 9608 8340 9636
rect 8392 9648 8444 9654
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7746 9072 7802 9081
rect 7746 9007 7802 9016
rect 7760 8974 7788 9007
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8634 7788 8910
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 4908 2746 5120 2774
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 4080 800 4108 2450
rect 4908 2310 4936 2746
rect 7760 2650 7788 5782
rect 7852 3058 7880 9454
rect 8220 8974 8248 9608
rect 8392 9590 8444 9596
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8128 8430 8156 8570
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8312 8090 8340 8774
rect 8404 8294 8432 9590
rect 8496 9382 8524 9862
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8496 9042 8524 9318
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8588 7478 8616 9862
rect 8666 9616 8722 9625
rect 8666 9551 8722 9560
rect 8680 8498 8708 9551
rect 8956 9110 8984 15302
rect 9048 13734 9076 20878
rect 9220 20800 9272 20806
rect 9220 20742 9272 20748
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9140 18766 9168 20402
rect 9232 20233 9260 20742
rect 9324 20641 9352 21626
rect 9600 21622 9628 22986
rect 10060 22642 10088 25502
rect 10152 24206 10180 25638
rect 10232 25220 10284 25226
rect 10232 25162 10284 25168
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 10060 22438 10088 22578
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 9864 22092 9916 22098
rect 10244 22094 10272 25162
rect 10704 22710 10732 26302
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26200 12586 27000
rect 13174 26330 13230 27000
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 10784 25492 10836 25498
rect 10784 25434 10836 25440
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10796 22098 10824 25434
rect 11256 22098 11284 26200
rect 11794 24032 11850 24041
rect 11794 23967 11850 23976
rect 11440 23854 11652 23882
rect 11440 23730 11468 23854
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 11520 23724 11572 23730
rect 11520 23666 11572 23672
rect 11532 23526 11560 23666
rect 11624 23526 11652 23854
rect 11520 23520 11572 23526
rect 11520 23462 11572 23468
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11428 23180 11480 23186
rect 11428 23122 11480 23128
rect 11440 22964 11468 23122
rect 11704 22976 11756 22982
rect 11440 22936 11704 22964
rect 11704 22918 11756 22924
rect 11808 22778 11836 23967
rect 11900 22778 11928 26200
rect 12164 25764 12216 25770
rect 12164 25706 12216 25712
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 12084 23633 12112 24006
rect 12070 23624 12126 23633
rect 12070 23559 12126 23568
rect 12176 23508 12204 25706
rect 12256 25356 12308 25362
rect 12256 25298 12308 25304
rect 12268 24614 12296 25298
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12268 23866 12296 24550
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12452 24070 12480 24142
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12544 23798 12572 26200
rect 12808 25628 12860 25634
rect 12808 25570 12860 25576
rect 12820 24206 12848 25570
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12808 24200 12860 24206
rect 12808 24142 12860 24148
rect 12532 23792 12584 23798
rect 12346 23760 12402 23769
rect 12256 23724 12308 23730
rect 12532 23734 12584 23740
rect 12346 23695 12402 23704
rect 12256 23666 12308 23672
rect 12084 23480 12204 23508
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11796 22636 11848 22642
rect 11796 22578 11848 22584
rect 11808 22166 11836 22578
rect 11796 22160 11848 22166
rect 11796 22102 11848 22108
rect 11980 22160 12032 22166
rect 11980 22102 12032 22108
rect 9864 22034 9916 22040
rect 10152 22066 10272 22094
rect 10784 22092 10836 22098
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9588 21616 9640 21622
rect 9588 21558 9640 21564
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 9508 21434 9536 21490
rect 9508 21406 9628 21434
rect 9600 21350 9628 21406
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9310 20632 9366 20641
rect 9310 20567 9366 20576
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9218 20224 9274 20233
rect 9218 20159 9274 20168
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9048 13394 9076 13466
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 9140 12170 9168 17614
rect 9232 17082 9260 20159
rect 9508 19786 9536 20538
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 9404 18964 9456 18970
rect 9404 18906 9456 18912
rect 9312 18828 9364 18834
rect 9312 18770 9364 18776
rect 9324 18193 9352 18770
rect 9310 18184 9366 18193
rect 9310 18119 9366 18128
rect 9324 17202 9352 18119
rect 9416 17610 9444 18906
rect 9508 18222 9536 19178
rect 9600 18358 9628 21286
rect 9692 20777 9720 21830
rect 9678 20768 9734 20777
rect 9678 20703 9734 20712
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9588 18352 9640 18358
rect 9588 18294 9640 18300
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9586 17776 9642 17785
rect 9692 17746 9720 20198
rect 9784 18970 9812 21830
rect 9876 20058 9904 22034
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9784 17814 9812 18770
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9876 18465 9904 18566
rect 9862 18456 9918 18465
rect 9862 18391 9918 18400
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9586 17711 9642 17720
rect 9680 17740 9732 17746
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9232 17054 9352 17082
rect 9220 15632 9272 15638
rect 9218 15600 9220 15609
rect 9272 15600 9274 15609
rect 9218 15535 9274 15544
rect 9232 15434 9260 15535
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9324 15366 9352 17054
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9324 14278 9352 14962
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9416 14414 9444 14758
rect 9508 14618 9536 17614
rect 9600 17270 9628 17711
rect 9680 17682 9732 17688
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9784 16998 9812 17750
rect 9876 17202 9904 18022
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9876 16561 9904 17138
rect 9862 16552 9918 16561
rect 9862 16487 9918 16496
rect 9772 16176 9824 16182
rect 9772 16118 9824 16124
rect 9784 15366 9812 16118
rect 9968 16046 9996 18770
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10060 17746 10088 18702
rect 10152 18086 10180 22066
rect 10784 22034 10836 22040
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10324 21480 10376 21486
rect 10520 21457 10548 21966
rect 10966 21856 11022 21865
rect 10966 21791 11022 21800
rect 10980 21690 11008 21791
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 11992 21554 12020 22102
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 10600 21480 10652 21486
rect 10324 21422 10376 21428
rect 10506 21448 10562 21457
rect 10336 21146 10364 21422
rect 10600 21422 10652 21428
rect 10506 21383 10562 21392
rect 10324 21140 10376 21146
rect 10324 21082 10376 21088
rect 10612 20874 10640 21422
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 10600 20868 10652 20874
rect 10600 20810 10652 20816
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10980 19718 11008 20334
rect 11072 19854 11100 21286
rect 11532 21010 11560 21286
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11426 20904 11482 20913
rect 11336 20868 11388 20874
rect 11426 20839 11482 20848
rect 11336 20810 11388 20816
rect 11348 20777 11376 20810
rect 11440 20806 11468 20839
rect 11428 20800 11480 20806
rect 11334 20768 11390 20777
rect 11428 20742 11480 20748
rect 11334 20703 11390 20712
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 11164 19786 11192 20198
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10874 19544 10930 19553
rect 10324 19508 10376 19514
rect 10874 19479 10876 19488
rect 10324 19450 10376 19456
rect 10928 19479 10930 19488
rect 10876 19450 10928 19456
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10244 18426 10272 18770
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10138 17912 10194 17921
rect 10138 17847 10140 17856
rect 10192 17847 10194 17856
rect 10140 17818 10192 17824
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9876 15366 9904 15438
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9600 14618 9628 14894
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9692 14482 9720 14894
rect 9784 14793 9812 15302
rect 9770 14784 9826 14793
rect 9770 14719 9826 14728
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 9048 5166 9076 12106
rect 9140 11762 9168 12106
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9140 10266 9168 11698
rect 9232 11218 9260 14010
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9324 12646 9352 13806
rect 9402 13424 9458 13433
rect 9402 13359 9404 13368
rect 9456 13359 9458 13368
rect 9404 13330 9456 13336
rect 9692 13258 9720 14214
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9324 12306 9352 12582
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9416 11642 9444 12786
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9324 11614 9444 11642
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9140 7546 9168 8842
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9232 7478 9260 10950
rect 9324 10062 9352 11614
rect 9404 11552 9456 11558
rect 9496 11552 9548 11558
rect 9404 11494 9456 11500
rect 9494 11520 9496 11529
rect 9548 11520 9550 11529
rect 9416 11286 9444 11494
rect 9494 11455 9550 11464
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9416 9042 9444 11018
rect 9508 10742 9536 11455
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9508 9586 9536 9998
rect 9692 9738 9720 12106
rect 9784 11150 9812 13126
rect 9876 11830 9904 15302
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 10060 14482 10088 15030
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10152 12866 10180 15982
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 10060 12838 10180 12866
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9876 11150 9904 11630
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9876 10470 9904 11086
rect 9968 10810 9996 12786
rect 10060 12782 10088 12838
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10046 11112 10102 11121
rect 10046 11047 10102 11056
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9692 9710 9812 9738
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9508 9450 9536 9522
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9508 8838 9536 9386
rect 9692 9178 9720 9522
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9508 8430 9536 8774
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 9692 4010 9720 8774
rect 9784 6662 9812 9710
rect 10060 8634 10088 11047
rect 10152 9178 10180 12718
rect 10244 11626 10272 18226
rect 10336 17882 10364 19450
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10598 19272 10654 19281
rect 10598 19207 10654 19216
rect 10506 18592 10562 18601
rect 10506 18527 10562 18536
rect 10414 18456 10470 18465
rect 10414 18391 10470 18400
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10336 15366 10364 17070
rect 10428 16726 10456 18391
rect 10520 18358 10548 18527
rect 10508 18352 10560 18358
rect 10508 18294 10560 18300
rect 10612 17921 10640 19207
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10704 18154 10732 18634
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 10598 17912 10654 17921
rect 10598 17847 10654 17856
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10416 16720 10468 16726
rect 10416 16662 10468 16668
rect 10428 16590 10456 16662
rect 10520 16590 10548 16934
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10612 16402 10640 17847
rect 10520 16374 10640 16402
rect 10520 16250 10548 16374
rect 10598 16280 10654 16289
rect 10508 16244 10560 16250
rect 10598 16215 10600 16224
rect 10508 16186 10560 16192
rect 10652 16215 10654 16224
rect 10600 16186 10652 16192
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10520 15094 10548 16186
rect 10612 15094 10640 16186
rect 10690 15872 10746 15881
rect 10690 15807 10746 15816
rect 10704 15638 10732 15807
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10692 15360 10744 15366
rect 10796 15337 10824 19314
rect 10980 19310 11008 19654
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11072 18873 11100 19110
rect 11058 18864 11114 18873
rect 10968 18828 11020 18834
rect 11164 18834 11192 19722
rect 11058 18799 11114 18808
rect 11152 18828 11204 18834
rect 10968 18770 11020 18776
rect 11152 18770 11204 18776
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10888 16794 10916 16934
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10980 16153 11008 18770
rect 11256 16538 11284 20198
rect 11348 20058 11376 20538
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11428 19440 11480 19446
rect 11426 19408 11428 19417
rect 11480 19408 11482 19417
rect 11426 19343 11482 19352
rect 11532 19258 11560 20946
rect 11440 19230 11560 19258
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11348 18630 11376 18702
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11072 16510 11284 16538
rect 10966 16144 11022 16153
rect 10966 16079 11022 16088
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10966 16008 11022 16017
rect 10888 15570 10916 15982
rect 10966 15943 10968 15952
rect 11020 15943 11022 15952
rect 10968 15914 11020 15920
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10876 15360 10928 15366
rect 10692 15302 10744 15308
rect 10782 15328 10838 15337
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 10600 15088 10652 15094
rect 10600 15030 10652 15036
rect 10324 14884 10376 14890
rect 10600 14884 10652 14890
rect 10376 14844 10548 14872
rect 10324 14826 10376 14832
rect 10322 14784 10378 14793
rect 10322 14719 10378 14728
rect 10336 14006 10364 14719
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 10336 12918 10364 13942
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10322 12608 10378 12617
rect 10322 12543 10378 12552
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 10336 11558 10364 12543
rect 10428 12238 10456 14418
rect 10520 12714 10548 14844
rect 10600 14826 10652 14832
rect 10612 14482 10640 14826
rect 10704 14482 10732 15302
rect 10876 15302 10928 15308
rect 10782 15263 10838 15272
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10612 12986 10640 14214
rect 10796 13870 10824 14894
rect 10888 14414 10916 15302
rect 11072 15042 11100 16510
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11164 15366 11192 16186
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11256 15162 11284 16390
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11072 15014 11284 15042
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10704 13462 10732 13670
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10690 12880 10746 12889
rect 10690 12815 10692 12824
rect 10744 12815 10746 12824
rect 10692 12786 10744 12792
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11898 10640 12038
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10520 11506 10548 11766
rect 10520 11478 10732 11506
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10244 9518 10272 10542
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10244 7954 10272 9454
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10336 7342 10364 9318
rect 10428 8634 10456 10474
rect 10612 9654 10640 11290
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10704 8922 10732 11478
rect 10796 11370 10824 13806
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10888 12442 10916 13330
rect 10980 12617 11008 14418
rect 11164 14278 11192 14758
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 10966 12608 11022 12617
rect 10966 12543 11022 12552
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10796 11342 11008 11370
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10796 10266 10824 11154
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10796 9450 10824 9862
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10888 9042 10916 11222
rect 10980 10606 11008 11342
rect 10968 10600 11020 10606
rect 11072 10577 11100 12038
rect 11164 10962 11192 14010
rect 11256 14006 11284 15014
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11256 11354 11284 13330
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11348 11064 11376 18226
rect 11440 13274 11468 19230
rect 11518 19000 11574 19009
rect 11518 18935 11574 18944
rect 11532 18737 11560 18935
rect 11518 18728 11574 18737
rect 11624 18714 11652 21490
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11808 21078 11836 21286
rect 11796 21072 11848 21078
rect 11796 21014 11848 21020
rect 12084 20942 12112 23480
rect 12268 23050 12296 23666
rect 12256 23044 12308 23050
rect 12256 22986 12308 22992
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12268 21554 12296 21830
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12254 21312 12310 21321
rect 12360 21298 12388 23695
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12452 22438 12480 23122
rect 12636 23089 12664 24142
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12622 23080 12678 23089
rect 12622 23015 12678 23024
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12452 21554 12480 22374
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12310 21270 12388 21298
rect 12254 21247 12310 21256
rect 11704 20936 11756 20942
rect 11704 20878 11756 20884
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 11716 19242 11744 20878
rect 11794 20632 11850 20641
rect 11794 20567 11850 20576
rect 11808 20534 11836 20567
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 11794 19816 11850 19825
rect 11794 19751 11850 19760
rect 11808 19718 11836 19751
rect 11900 19718 11928 19994
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 12164 19508 12216 19514
rect 12360 19496 12388 21270
rect 12452 20534 12480 21490
rect 12544 21010 12572 22714
rect 12636 21894 12664 22918
rect 12728 22817 12756 23462
rect 12820 22982 12848 23666
rect 13188 23526 13216 24210
rect 13176 23520 13228 23526
rect 13176 23462 13228 23468
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12900 23248 12952 23254
rect 12900 23190 12952 23196
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12714 22808 12770 22817
rect 12714 22743 12770 22752
rect 12820 22710 12848 22918
rect 12808 22704 12860 22710
rect 12808 22646 12860 22652
rect 12912 22556 12940 23190
rect 12820 22528 12940 22556
rect 12820 22030 12848 22528
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13372 22098 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15750 26200 15806 27000
rect 16394 26330 16450 27000
rect 16132 26302 16450 26330
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 13464 23254 13492 25230
rect 13832 24138 13860 26200
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13452 23248 13504 23254
rect 13452 23190 13504 23196
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 13464 21570 13492 22374
rect 13372 21542 13492 21570
rect 13372 21486 13400 21542
rect 13360 21480 13412 21486
rect 13556 21434 13584 23666
rect 13728 23588 13780 23594
rect 13728 23530 13780 23536
rect 13740 23361 13768 23530
rect 13726 23352 13782 23361
rect 13726 23287 13782 23296
rect 13636 23180 13688 23186
rect 13636 23122 13688 23128
rect 13648 22778 13676 23122
rect 13912 23112 13964 23118
rect 13910 23080 13912 23089
rect 13964 23080 13966 23089
rect 13910 23015 13966 23024
rect 13636 22772 13688 22778
rect 13636 22714 13688 22720
rect 13360 21422 13412 21428
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12452 19990 12480 20470
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12544 20233 12572 20334
rect 12716 20256 12768 20262
rect 12530 20224 12586 20233
rect 12716 20198 12768 20204
rect 12530 20159 12586 20168
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12164 19450 12216 19456
rect 12268 19468 12388 19496
rect 12438 19544 12494 19553
rect 12438 19479 12494 19488
rect 11888 19440 11940 19446
rect 12176 19394 12204 19450
rect 11940 19388 12204 19394
rect 11888 19382 12204 19388
rect 11900 19366 12204 19382
rect 11704 19236 11756 19242
rect 11704 19178 11756 19184
rect 11888 18760 11940 18766
rect 11624 18686 11836 18714
rect 11888 18702 11940 18708
rect 11518 18663 11574 18672
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11518 17640 11574 17649
rect 11518 17575 11574 17584
rect 11532 16969 11560 17575
rect 11624 16998 11652 18566
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11808 17626 11836 18686
rect 11900 18426 11928 18702
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 11900 18057 11928 18090
rect 11886 18048 11942 18057
rect 11886 17983 11942 17992
rect 11888 17808 11940 17814
rect 11886 17776 11888 17785
rect 11940 17776 11942 17785
rect 11886 17711 11942 17720
rect 11992 17678 12020 19366
rect 12268 19334 12296 19468
rect 12176 19306 12296 19334
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12084 18086 12112 18566
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 11980 17672 12032 17678
rect 11716 17218 11744 17614
rect 11808 17598 11928 17626
rect 11980 17614 12032 17620
rect 11716 17202 11836 17218
rect 11716 17196 11848 17202
rect 11716 17190 11796 17196
rect 11796 17138 11848 17144
rect 11612 16992 11664 16998
rect 11518 16960 11574 16969
rect 11612 16934 11664 16940
rect 11518 16895 11574 16904
rect 11532 16250 11560 16895
rect 11624 16658 11652 16934
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11532 14498 11560 15438
rect 11624 14906 11652 16594
rect 11716 15026 11744 16730
rect 11808 16697 11836 17138
rect 11794 16688 11850 16697
rect 11794 16623 11850 16632
rect 11900 16454 11928 17598
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11992 16114 12020 17614
rect 12084 16998 12112 18022
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11808 15502 11836 15846
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 12070 15464 12126 15473
rect 12070 15399 12126 15408
rect 12084 15366 12112 15399
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11978 15056 12034 15065
rect 11704 15020 11756 15026
rect 11978 14991 11980 15000
rect 11704 14962 11756 14968
rect 12032 14991 12034 15000
rect 11980 14962 12032 14968
rect 11796 14952 11848 14958
rect 11624 14878 11744 14906
rect 11796 14894 11848 14900
rect 11532 14470 11652 14498
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11532 13462 11560 14282
rect 11624 14006 11652 14470
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11440 13246 11560 13274
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 11529 11468 12582
rect 11426 11520 11482 11529
rect 11426 11455 11482 11464
rect 11532 11121 11560 13246
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11624 12170 11652 13126
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11624 11830 11652 12106
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11518 11112 11574 11121
rect 11348 11036 11468 11064
rect 11518 11047 11574 11056
rect 11164 10934 11376 10962
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 10968 10542 11020 10548
rect 11058 10568 11114 10577
rect 11058 10503 11114 10512
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 10980 9518 11008 10134
rect 11072 10062 11100 10202
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10704 8894 10824 8922
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 6748 800 6776 2450
rect 8312 2446 8340 2790
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9416 800 9444 2450
rect 9784 2446 9812 3130
rect 10428 3126 10456 8366
rect 10520 6866 10548 8570
rect 10704 8566 10732 8774
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10612 3738 10640 8366
rect 10796 4690 10824 8894
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10980 7546 11008 8842
rect 11072 8498 11100 9114
rect 11164 8634 11192 10746
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11256 10062 11284 10542
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11256 9518 11284 9998
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11348 8022 11376 10934
rect 11440 9994 11468 11036
rect 11518 10568 11574 10577
rect 11518 10503 11574 10512
rect 11532 10470 11560 10503
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11426 9888 11482 9897
rect 11426 9823 11482 9832
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11440 6254 11468 9823
rect 11532 8634 11560 10202
rect 11624 9178 11652 11290
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11716 8090 11744 14878
rect 11808 14550 11836 14894
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11886 14512 11942 14521
rect 11886 14447 11942 14456
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11808 13462 11836 13942
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11808 10470 11836 11766
rect 11900 10810 11928 14447
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11992 13394 12020 14350
rect 12176 14090 12204 19306
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12268 17610 12296 18906
rect 12360 17882 12388 19246
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 12268 16726 12296 17070
rect 12360 17066 12388 17818
rect 12452 17338 12480 19479
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12530 17504 12586 17513
rect 12530 17439 12586 17448
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12348 17060 12400 17066
rect 12348 17002 12400 17008
rect 12544 16969 12572 17439
rect 12530 16960 12586 16969
rect 12530 16895 12586 16904
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12360 16046 12388 16594
rect 12544 16182 12572 16594
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12268 15201 12296 15982
rect 12254 15192 12310 15201
rect 12254 15127 12310 15136
rect 12176 14074 12296 14090
rect 12176 14068 12308 14074
rect 12176 14062 12256 14068
rect 12256 14010 12308 14016
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 12176 12646 12204 13942
rect 12360 13802 12388 15982
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12256 12708 12308 12714
rect 12256 12650 12308 12656
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12268 12306 12296 12650
rect 12360 12306 12388 13194
rect 12452 12986 12480 15846
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12438 12744 12494 12753
rect 12438 12679 12494 12688
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12084 11558 12112 12242
rect 12268 11937 12296 12242
rect 12254 11928 12310 11937
rect 12254 11863 12310 11872
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11992 11393 12020 11494
rect 11978 11384 12034 11393
rect 11978 11319 12034 11328
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 12084 10690 12112 11494
rect 12360 11354 12388 12242
rect 12452 11914 12480 12679
rect 12544 12442 12572 15302
rect 12636 14890 12664 18022
rect 12728 17728 12756 20198
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 19922 13400 21422
rect 13464 21406 13584 21434
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13268 19780 13320 19786
rect 13268 19722 13320 19728
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13188 19310 13216 19654
rect 13280 19378 13308 19722
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 13188 19174 13216 19246
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13372 18766 13400 19654
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 13188 18601 13216 18634
rect 13174 18592 13230 18601
rect 13174 18527 13230 18536
rect 13188 18222 13216 18527
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 12820 17864 12848 18090
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12820 17836 12940 17864
rect 12912 17746 12940 17836
rect 13268 17808 13320 17814
rect 13266 17776 13268 17785
rect 13320 17776 13322 17785
rect 12900 17740 12952 17746
rect 12728 17700 12848 17728
rect 12820 17354 12848 17700
rect 13266 17711 13322 17720
rect 12900 17682 12952 17688
rect 12728 17326 12848 17354
rect 13360 17332 13412 17338
rect 12728 15586 12756 17326
rect 13360 17274 13412 17280
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12820 16833 12848 17206
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12806 16824 12862 16833
rect 12950 16827 13258 16836
rect 13372 16833 13400 17274
rect 13464 17218 13492 21406
rect 13544 21344 13596 21350
rect 13648 21298 13676 22714
rect 14096 21956 14148 21962
rect 14096 21898 14148 21904
rect 14108 21486 14136 21898
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 13596 21292 13676 21298
rect 13544 21286 13676 21292
rect 13556 21270 13676 21286
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13556 18698 13584 20470
rect 13544 18692 13596 18698
rect 13544 18634 13596 18640
rect 13648 18601 13676 21270
rect 13910 21176 13966 21185
rect 13910 21111 13966 21120
rect 13924 20806 13952 21111
rect 14096 20868 14148 20874
rect 14096 20810 14148 20816
rect 13912 20800 13964 20806
rect 13910 20768 13912 20777
rect 13964 20768 13966 20777
rect 13910 20703 13966 20712
rect 13818 20496 13874 20505
rect 13818 20431 13874 20440
rect 13832 20058 13860 20431
rect 14004 20392 14056 20398
rect 14004 20334 14056 20340
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13634 18592 13690 18601
rect 13634 18527 13690 18536
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13556 17610 13584 18022
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13464 17190 13584 17218
rect 13452 17060 13504 17066
rect 13452 17002 13504 17008
rect 12806 16759 12862 16768
rect 13358 16824 13414 16833
rect 13358 16759 13414 16768
rect 12992 16720 13044 16726
rect 12990 16688 12992 16697
rect 13268 16720 13320 16726
rect 13044 16688 13046 16697
rect 13268 16662 13320 16668
rect 12990 16623 13046 16632
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12820 15706 12848 16458
rect 13280 15994 13308 16662
rect 13280 15966 13400 15994
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13372 15745 13400 15966
rect 13358 15736 13414 15745
rect 12808 15700 12860 15706
rect 13358 15671 13414 15680
rect 12808 15642 12860 15648
rect 13464 15586 13492 17002
rect 13556 16726 13584 17190
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13556 15706 13584 16458
rect 13648 16250 13676 17682
rect 13740 17338 13768 18362
rect 14016 18358 14044 20334
rect 14108 19700 14136 20810
rect 14200 20058 14228 24142
rect 14292 24070 14320 24686
rect 14476 24342 14504 26200
rect 15016 25016 15068 25022
rect 15016 24958 15068 24964
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14740 24676 14792 24682
rect 14740 24618 14792 24624
rect 14464 24336 14516 24342
rect 14464 24278 14516 24284
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14280 24064 14332 24070
rect 14476 24041 14504 24142
rect 14280 24006 14332 24012
rect 14462 24032 14518 24041
rect 14462 23967 14518 23976
rect 14476 23497 14504 23967
rect 14462 23488 14518 23497
rect 14462 23423 14518 23432
rect 14370 23352 14426 23361
rect 14370 23287 14426 23296
rect 14384 23118 14412 23287
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14568 22778 14596 22918
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14752 22166 14780 24618
rect 14740 22160 14792 22166
rect 14740 22102 14792 22108
rect 14370 21992 14426 22001
rect 14370 21927 14372 21936
rect 14424 21927 14426 21936
rect 14372 21898 14424 21904
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14660 21078 14688 21490
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14648 21072 14700 21078
rect 14648 21014 14700 21020
rect 14752 20398 14780 21286
rect 14844 20641 14872 24890
rect 14922 24304 14978 24313
rect 14922 24239 14978 24248
rect 14936 23633 14964 24239
rect 14922 23624 14978 23633
rect 14922 23559 14978 23568
rect 15028 22642 15056 24958
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 15120 22098 15148 26200
rect 15660 25152 15712 25158
rect 15660 25094 15712 25100
rect 15476 25084 15528 25090
rect 15476 25026 15528 25032
rect 15200 24880 15252 24886
rect 15200 24822 15252 24828
rect 15108 22092 15160 22098
rect 15108 22034 15160 22040
rect 15212 22030 15240 24822
rect 15384 24132 15436 24138
rect 15384 24074 15436 24080
rect 15200 22024 15252 22030
rect 14922 21992 14978 22001
rect 15200 21966 15252 21972
rect 14922 21927 14924 21936
rect 14976 21927 14978 21936
rect 14924 21898 14976 21904
rect 14936 21457 14964 21898
rect 15108 21616 15160 21622
rect 15108 21558 15160 21564
rect 14922 21448 14978 21457
rect 14922 21383 14978 21392
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14936 21010 14964 21286
rect 14924 21004 14976 21010
rect 14924 20946 14976 20952
rect 14924 20800 14976 20806
rect 14924 20742 14976 20748
rect 14830 20632 14886 20641
rect 14830 20567 14886 20576
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14188 19712 14240 19718
rect 14108 19672 14188 19700
rect 14188 19654 14240 19660
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 14004 17604 14056 17610
rect 14004 17546 14056 17552
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13728 16992 13780 16998
rect 13726 16960 13728 16969
rect 13780 16960 13782 16969
rect 13726 16895 13782 16904
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 12728 15558 12848 15586
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 14074 12664 14214
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12452 11886 12572 11914
rect 12438 11792 12494 11801
rect 12438 11727 12494 11736
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12346 11112 12402 11121
rect 12256 11076 12308 11082
rect 12346 11047 12402 11056
rect 12256 11018 12308 11024
rect 12268 10849 12296 11018
rect 12254 10840 12310 10849
rect 12254 10775 12310 10784
rect 11992 10662 12112 10690
rect 11992 10538 12020 10662
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11900 10418 11928 10474
rect 11808 9994 11836 10406
rect 11900 10390 12112 10418
rect 12084 10266 12112 10390
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11992 10130 12020 10202
rect 12268 10146 12296 10775
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 12084 10118 12296 10146
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11900 9874 11928 10066
rect 11980 9988 12032 9994
rect 12084 9976 12112 10118
rect 12032 9948 12112 9976
rect 11980 9930 12032 9936
rect 12164 9920 12216 9926
rect 11900 9868 12164 9874
rect 11900 9862 12216 9868
rect 11900 9846 12204 9862
rect 11900 9654 11928 9846
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 12070 9480 12126 9489
rect 12070 9415 12126 9424
rect 12084 8430 12112 9415
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12176 8634 12204 9318
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12268 8634 12296 8978
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12360 8430 12388 11047
rect 12452 8838 12480 11727
rect 12544 9466 12572 11886
rect 12544 9438 12756 9466
rect 12728 9382 12756 9438
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12544 9178 12572 9318
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12820 8906 12848 15558
rect 13360 15564 13412 15570
rect 13464 15558 13584 15586
rect 13360 15506 13412 15512
rect 13372 15450 13400 15506
rect 13372 15422 13492 15450
rect 13266 15192 13322 15201
rect 13266 15127 13322 15136
rect 13280 14958 13308 15127
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13372 14618 13400 14962
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13464 14482 13492 15422
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 12898 14376 12954 14385
rect 13556 14362 13584 15558
rect 13648 15502 13676 15914
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13740 15008 13768 15846
rect 12898 14311 12954 14320
rect 13372 14334 13584 14362
rect 13648 14980 13768 15008
rect 12912 14278 12940 14311
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13096 13870 13124 14010
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 12900 12640 12952 12646
rect 13096 12628 13124 12786
rect 12952 12600 13124 12628
rect 12900 12582 12952 12588
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13372 12434 13400 14334
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13096 12406 13400 12434
rect 13096 11801 13124 12406
rect 13176 12232 13228 12238
rect 13228 12180 13400 12186
rect 13176 12174 13400 12180
rect 13188 12158 13400 12174
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13082 11792 13138 11801
rect 13082 11727 13138 11736
rect 13188 11626 13216 12038
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13372 11354 13400 12158
rect 13464 11354 13492 12786
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 12898 10840 12954 10849
rect 12898 10775 12954 10784
rect 12912 10742 12940 10775
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13372 9450 13400 11154
rect 13556 10130 13584 13874
rect 13648 13190 13676 14980
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14618 13768 14826
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13832 14550 13860 14758
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13740 13462 13768 14418
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13636 12912 13688 12918
rect 13740 12900 13768 13194
rect 13832 13190 13860 13806
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13688 12872 13768 12900
rect 13820 12912 13872 12918
rect 13636 12854 13688 12860
rect 13820 12854 13872 12860
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13740 12170 13768 12310
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13832 11898 13860 12854
rect 13924 12102 13952 17138
rect 14016 16182 14044 17546
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 14016 15366 14044 16118
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 14016 14346 14044 15302
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14016 13326 14044 14282
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 14016 13161 14044 13262
rect 14108 13258 14136 19314
rect 14200 19174 14228 19654
rect 14476 19446 14504 19790
rect 14568 19514 14596 19790
rect 14844 19514 14872 20567
rect 14556 19508 14608 19514
rect 14832 19508 14884 19514
rect 14556 19450 14608 19456
rect 14752 19468 14832 19496
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14384 18970 14412 19110
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14476 18902 14504 19110
rect 14464 18896 14516 18902
rect 14464 18838 14516 18844
rect 14476 18737 14504 18838
rect 14462 18728 14518 18737
rect 14462 18663 14518 18672
rect 14568 18358 14596 19450
rect 14648 19304 14700 19310
rect 14752 19292 14780 19468
rect 14832 19450 14884 19456
rect 14936 19394 14964 20742
rect 15120 20618 15148 21558
rect 15212 21146 15240 21966
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15028 20590 15332 20618
rect 15028 19718 15056 20590
rect 15304 20534 15332 20590
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15108 20324 15160 20330
rect 15108 20266 15160 20272
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 14936 19366 15056 19394
rect 14700 19264 14780 19292
rect 14924 19304 14976 19310
rect 14922 19272 14924 19281
rect 14976 19272 14978 19281
rect 14648 19246 14700 19252
rect 14922 19207 14978 19216
rect 14832 18964 14884 18970
rect 15028 18952 15056 19366
rect 15120 19310 15148 20266
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 14832 18906 14884 18912
rect 14936 18924 15056 18952
rect 14844 18766 14872 18906
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14556 18352 14608 18358
rect 14556 18294 14608 18300
rect 14738 18048 14794 18057
rect 14738 17983 14794 17992
rect 14462 17640 14518 17649
rect 14462 17575 14518 17584
rect 14476 17542 14504 17575
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14292 17338 14320 17478
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14370 16552 14426 16561
rect 14370 16487 14426 16496
rect 14384 16454 14412 16487
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14292 14550 14320 14894
rect 14188 14544 14240 14550
rect 14188 14486 14240 14492
rect 14280 14544 14332 14550
rect 14280 14486 14332 14492
rect 14200 14074 14228 14486
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14292 13326 14320 14486
rect 14384 13530 14412 15302
rect 14476 13870 14504 16594
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14002 13152 14058 13161
rect 14002 13087 14058 13096
rect 13912 12096 13964 12102
rect 14016 12084 14044 13087
rect 14200 12782 14228 13194
rect 14292 12918 14320 13262
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14200 12102 14228 12718
rect 14476 12434 14504 13670
rect 14568 12986 14596 15506
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14476 12406 14596 12434
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14096 12096 14148 12102
rect 14016 12056 14096 12084
rect 13912 12038 13964 12044
rect 14096 12038 14148 12044
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 14108 11014 14136 12038
rect 14476 11150 14504 12174
rect 14568 11626 14596 12406
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 13832 10849 13860 10950
rect 13818 10840 13874 10849
rect 13818 10775 13874 10784
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13648 10266 13676 10610
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13832 10198 13860 10775
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13832 9722 13860 10134
rect 14476 10062 14504 11086
rect 14660 10538 14688 16526
rect 14752 14618 14780 17983
rect 14936 16046 14964 18924
rect 15014 18864 15070 18873
rect 15014 18799 15070 18808
rect 15108 18828 15160 18834
rect 15028 18154 15056 18799
rect 15212 18816 15240 20334
rect 15396 19281 15424 24074
rect 15488 23118 15516 25026
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15488 21010 15516 22918
rect 15566 21448 15622 21457
rect 15566 21383 15568 21392
rect 15620 21383 15622 21392
rect 15568 21354 15620 21360
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15568 20528 15620 20534
rect 15568 20470 15620 20476
rect 15580 20262 15608 20470
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15488 19922 15516 20198
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15672 19378 15700 25094
rect 15764 23798 15792 26200
rect 15844 25424 15896 25430
rect 15844 25366 15896 25372
rect 15752 23792 15804 23798
rect 15752 23734 15804 23740
rect 15750 21584 15806 21593
rect 15856 21570 15884 25366
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15948 23866 15976 24550
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 16026 23760 16082 23769
rect 16026 23695 16082 23704
rect 16040 21690 16068 23695
rect 16132 22710 16160 26302
rect 16394 26200 16450 26302
rect 17038 26330 17094 27000
rect 17682 26330 17738 27000
rect 17038 26302 17356 26330
rect 17038 26200 17094 26302
rect 16210 25256 16266 25265
rect 16210 25191 16266 25200
rect 16224 24274 16252 25191
rect 16212 24268 16264 24274
rect 16212 24210 16264 24216
rect 17224 24132 17276 24138
rect 17224 24074 17276 24080
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 17040 24064 17092 24070
rect 17040 24006 17092 24012
rect 16960 23730 16988 24006
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 16868 23202 16896 23666
rect 17052 23662 17080 24006
rect 17236 23866 17264 24074
rect 17132 23860 17184 23866
rect 17132 23802 17184 23808
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 16868 23174 16988 23202
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 16764 22704 16816 22710
rect 16764 22646 16816 22652
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 15936 21616 15988 21622
rect 15806 21542 15884 21570
rect 15750 21519 15806 21528
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15382 19272 15438 19281
rect 15382 19207 15438 19216
rect 15566 19272 15622 19281
rect 15566 19207 15622 19216
rect 15160 18788 15240 18816
rect 15108 18770 15160 18776
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 15198 18456 15254 18465
rect 15198 18391 15254 18400
rect 15212 18290 15240 18391
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15016 18148 15068 18154
rect 15016 18090 15068 18096
rect 15120 17542 15148 18158
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15028 16114 15056 17478
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14844 15502 14872 15642
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14936 15094 14964 15846
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 14924 15088 14976 15094
rect 14924 15030 14976 15036
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14936 14618 14964 14894
rect 14740 14612 14792 14618
rect 14924 14612 14976 14618
rect 14792 14572 14872 14600
rect 14740 14554 14792 14560
rect 14844 14074 14872 14572
rect 14924 14554 14976 14560
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14936 13870 14964 14554
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14832 13796 14884 13802
rect 14832 13738 14884 13744
rect 14844 13258 14872 13738
rect 15028 13530 15056 15370
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14752 12170 14780 12786
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14832 12164 14884 12170
rect 14832 12106 14884 12112
rect 14752 10810 14780 12106
rect 14844 11354 14872 12106
rect 15028 11694 15056 13466
rect 15120 12850 15148 17478
rect 15212 13802 15240 17818
rect 15304 17134 15332 18566
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15304 15858 15332 16934
rect 15396 16590 15424 17478
rect 15580 16590 15608 19207
rect 15672 18068 15700 19314
rect 15764 19009 15792 20742
rect 15750 19000 15806 19009
rect 15750 18935 15806 18944
rect 15856 18578 15884 21542
rect 15934 21584 15936 21593
rect 15988 21584 15990 21593
rect 15934 21519 15990 21528
rect 16132 20602 16160 22170
rect 16408 21010 16436 22170
rect 16776 21894 16804 22646
rect 16868 22574 16896 23054
rect 16960 22681 16988 23174
rect 17052 23050 17080 23598
rect 17040 23044 17092 23050
rect 17040 22986 17092 22992
rect 16946 22672 17002 22681
rect 16946 22607 17002 22616
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16764 21888 16816 21894
rect 16764 21830 16816 21836
rect 16578 21312 16634 21321
rect 16578 21247 16634 21256
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16592 20942 16620 21247
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16040 19174 16068 20402
rect 16592 20330 16620 20538
rect 16580 20324 16632 20330
rect 16580 20266 16632 20272
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16132 19786 16160 20198
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16118 19544 16174 19553
rect 16118 19479 16174 19488
rect 16132 19174 16160 19479
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 15856 18550 15976 18578
rect 15752 18080 15804 18086
rect 15672 18040 15752 18068
rect 15752 18022 15804 18028
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15382 15872 15438 15881
rect 15304 15830 15382 15858
rect 15382 15807 15438 15816
rect 15396 15094 15424 15807
rect 15488 15706 15516 15982
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15488 15162 15516 15302
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15396 14346 15424 15030
rect 15580 14958 15608 16390
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15566 14784 15622 14793
rect 15566 14719 15622 14728
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15212 12782 15240 13330
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15304 13161 15332 13194
rect 15290 13152 15346 13161
rect 15290 13087 15346 13096
rect 15304 12986 15332 13087
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 15120 11354 15148 12650
rect 15198 12608 15254 12617
rect 15198 12543 15254 12552
rect 15212 12306 15240 12543
rect 15304 12374 15332 12718
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15488 12374 15516 12650
rect 15292 12368 15344 12374
rect 15292 12310 15344 12316
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15580 11898 15608 14719
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15028 11082 15056 11154
rect 15488 11082 15516 11766
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 8090 12480 8230
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 12084 3738 12112 7822
rect 12452 7818 12480 8026
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12636 5846 12664 8434
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12820 7750 12848 8366
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 13648 7818 13676 9658
rect 14476 9518 14504 9998
rect 14464 9512 14516 9518
rect 14740 9512 14792 9518
rect 14464 9454 14516 9460
rect 14738 9480 14740 9489
rect 14792 9480 14794 9489
rect 14738 9415 14794 9424
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 13740 9042 13768 9318
rect 14200 9178 14228 9318
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 14844 8634 14872 10610
rect 15028 9926 15056 11018
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15212 10130 15240 10542
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 15028 9110 15056 9862
rect 15396 9110 15424 10950
rect 15488 10305 15516 11018
rect 15672 10470 15700 17138
rect 15764 13938 15792 18022
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 15856 15706 15884 17070
rect 15948 16590 15976 18550
rect 16040 18358 16068 18634
rect 16028 18352 16080 18358
rect 16028 18294 16080 18300
rect 16040 17542 16068 18294
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 16132 15366 16160 19110
rect 16212 18828 16264 18834
rect 16316 18816 16344 19246
rect 16264 18788 16344 18816
rect 16212 18770 16264 18776
rect 16212 17808 16264 17814
rect 16212 17750 16264 17756
rect 16224 17338 16252 17750
rect 16316 17746 16344 18788
rect 16408 18630 16436 19654
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 16500 18902 16528 19178
rect 16580 19168 16632 19174
rect 16578 19136 16580 19145
rect 16632 19136 16634 19145
rect 16578 19071 16634 19080
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 16592 18714 16620 19071
rect 16684 18834 16712 20742
rect 16776 20602 16804 21830
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 16764 20324 16816 20330
rect 16764 20266 16816 20272
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 16500 18686 16620 18714
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16394 18320 16450 18329
rect 16394 18255 16450 18264
rect 16408 18086 16436 18255
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16408 17882 16436 18022
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16304 17740 16356 17746
rect 16500 17728 16528 18686
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16304 17682 16356 17688
rect 16408 17700 16528 17728
rect 16408 17626 16436 17700
rect 16316 17598 16436 17626
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16316 17218 16344 17598
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16224 17190 16344 17218
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16224 14385 16252 17190
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16316 14822 16344 16594
rect 16408 16454 16436 17478
rect 16592 16697 16620 18226
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16684 17202 16712 17818
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16578 16688 16634 16697
rect 16578 16623 16634 16632
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16408 15910 16436 16390
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16488 16176 16540 16182
rect 16684 16130 16712 16186
rect 16488 16118 16540 16124
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16408 15094 16436 15302
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16316 14482 16344 14758
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 15842 14376 15898 14385
rect 15842 14311 15898 14320
rect 16210 14376 16266 14385
rect 16210 14311 16266 14320
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15474 10296 15530 10305
rect 15474 10231 15530 10240
rect 15488 9994 15516 10231
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15016 9104 15068 9110
rect 15016 9046 15068 9052
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15764 9042 15792 10678
rect 15856 10266 15884 14311
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15948 12434 15976 13874
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16224 13190 16252 13806
rect 16408 13394 16436 14214
rect 16500 13394 16528 16118
rect 16592 16102 16712 16130
rect 16592 16046 16620 16102
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16580 15904 16632 15910
rect 16578 15872 16580 15881
rect 16632 15872 16634 15881
rect 16578 15807 16634 15816
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16592 14074 16620 14214
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16684 14006 16712 15982
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16672 13728 16724 13734
rect 16672 13670 16724 13676
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16684 12986 16712 13670
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 15948 12406 16068 12434
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15948 9178 15976 11698
rect 16040 9382 16068 12406
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16684 12170 16712 12242
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16486 11112 16542 11121
rect 16486 11047 16488 11056
rect 16540 11047 16542 11056
rect 16488 11018 16540 11024
rect 16592 11014 16620 12038
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16132 9382 16160 10542
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16224 9722 16252 10066
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 15856 8566 15884 9046
rect 16132 8922 16160 9318
rect 16132 8906 16252 8922
rect 16132 8900 16264 8906
rect 16132 8894 16212 8900
rect 16212 8842 16264 8848
rect 16316 8634 16344 10542
rect 16592 10305 16620 10950
rect 16578 10296 16634 10305
rect 16578 10231 16580 10240
rect 16632 10231 16634 10240
rect 16580 10202 16632 10208
rect 16592 9926 16620 10202
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16592 9674 16620 9862
rect 16408 9654 16620 9674
rect 16396 9648 16620 9654
rect 16448 9646 16620 9648
rect 16776 9602 16804 20266
rect 16868 19310 16896 22510
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16960 20602 16988 20742
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 16946 20088 17002 20097
rect 16946 20023 17002 20032
rect 16960 19922 16988 20023
rect 17052 19990 17080 20742
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16868 19009 16896 19110
rect 16854 19000 16910 19009
rect 16854 18935 16910 18944
rect 16868 18057 16896 18935
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 16948 18624 17000 18630
rect 17052 18601 17080 18702
rect 16948 18566 17000 18572
rect 17038 18592 17094 18601
rect 16960 18222 16988 18566
rect 17038 18527 17094 18536
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16854 18048 16910 18057
rect 16854 17983 16910 17992
rect 16960 17746 16988 18158
rect 17144 17921 17172 23802
rect 17222 22672 17278 22681
rect 17222 22607 17278 22616
rect 17236 21865 17264 22607
rect 17222 21856 17278 21865
rect 17222 21791 17278 21800
rect 17328 21486 17356 26302
rect 17420 26302 17738 26330
rect 17420 23186 17448 26302
rect 17682 26200 17738 26302
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26200 20958 27000
rect 21546 26200 21602 27000
rect 22190 26200 22246 27000
rect 22834 26200 22890 27000
rect 23478 26200 23534 27000
rect 24122 26200 24178 27000
rect 24766 26200 24822 27000
rect 25410 26330 25466 27000
rect 24964 26302 25466 26330
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23798 18368 26200
rect 18984 25265 19012 26200
rect 18970 25256 19026 25265
rect 18970 25191 19026 25200
rect 18418 24440 18474 24449
rect 18418 24375 18474 24384
rect 18432 24041 18460 24375
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18418 24032 18474 24041
rect 18418 23967 18474 23976
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 18708 23730 18736 24210
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19156 24200 19208 24206
rect 19156 24142 19208 24148
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18800 23866 18828 24074
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 18696 23724 18748 23730
rect 18696 23666 18748 23672
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17500 21956 17552 21962
rect 17500 21898 17552 21904
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17236 20074 17264 21354
rect 17408 20936 17460 20942
rect 17406 20904 17408 20913
rect 17460 20904 17462 20913
rect 17406 20839 17462 20848
rect 17512 20330 17540 21898
rect 17592 21616 17644 21622
rect 17592 21558 17644 21564
rect 17604 20806 17632 21558
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17500 20324 17552 20330
rect 17500 20266 17552 20272
rect 17236 20046 17356 20074
rect 17604 20058 17632 20402
rect 17224 19984 17276 19990
rect 17222 19952 17224 19961
rect 17276 19952 17278 19961
rect 17222 19887 17278 19896
rect 17328 19496 17356 20046
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17696 19922 17724 20742
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 17788 19802 17816 23462
rect 17880 23322 17908 23598
rect 18708 23526 18736 23666
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18800 22778 18828 23802
rect 19076 23798 19104 24142
rect 18880 23792 18932 23798
rect 18880 23734 18932 23740
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 18892 23254 18920 23734
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 19076 23050 19104 23734
rect 19064 23044 19116 23050
rect 19064 22986 19116 22992
rect 19076 22778 19104 22986
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18156 21962 18184 22510
rect 18144 21956 18196 21962
rect 18196 21916 18368 21944
rect 18144 21898 18196 21904
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18340 20602 18368 21916
rect 18418 21176 18474 21185
rect 18418 21111 18474 21120
rect 18432 20806 18460 21111
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 18328 20596 18380 20602
rect 18328 20538 18380 20544
rect 18340 20262 18368 20538
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 17696 19774 17816 19802
rect 18328 19780 18380 19786
rect 17236 19468 17356 19496
rect 17408 19508 17460 19514
rect 17130 17912 17186 17921
rect 17130 17847 17186 17856
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 17236 17490 17264 19468
rect 17460 19468 17540 19496
rect 17408 19450 17460 19456
rect 17512 19378 17540 19468
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 17500 19372 17552 19378
rect 17500 19314 17552 19320
rect 16960 17462 17264 17490
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16868 16794 16896 16934
rect 16960 16833 16988 17462
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 16946 16824 17002 16833
rect 16856 16788 16908 16794
rect 16946 16759 17002 16768
rect 16856 16730 16908 16736
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16946 16416 17002 16425
rect 16868 14346 16896 16390
rect 16946 16351 17002 16360
rect 16960 16250 16988 16351
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17052 15502 17080 17002
rect 17144 16794 17172 17274
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17236 16658 17264 17138
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17130 16280 17186 16289
rect 17130 16215 17132 16224
rect 17184 16215 17186 16224
rect 17132 16186 17184 16192
rect 17328 15586 17356 19314
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17408 19168 17460 19174
rect 17406 19136 17408 19145
rect 17460 19136 17462 19145
rect 17406 19071 17462 19080
rect 17604 18630 17632 19246
rect 17696 19145 17724 19774
rect 18328 19722 18380 19728
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17774 19544 17830 19553
rect 17950 19547 18258 19556
rect 17830 19488 18000 19496
rect 17774 19479 18000 19488
rect 17788 19468 18000 19479
rect 17972 19428 18000 19468
rect 18052 19440 18104 19446
rect 17972 19400 18052 19428
rect 18052 19382 18104 19388
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17682 19136 17738 19145
rect 17682 19071 17738 19080
rect 18064 18766 18092 19246
rect 18156 19174 18184 19314
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18340 18902 18368 19722
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17590 18320 17646 18329
rect 17590 18255 17646 18264
rect 18326 18320 18382 18329
rect 18326 18255 18382 18264
rect 17604 18222 17632 18255
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17592 18216 17644 18222
rect 17592 18158 17644 18164
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17236 15558 17356 15586
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16948 14884 17000 14890
rect 16948 14826 17000 14832
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16960 14090 16988 14826
rect 17052 14498 17080 15438
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17144 14929 17172 14962
rect 17130 14920 17186 14929
rect 17130 14855 17186 14864
rect 17052 14482 17172 14498
rect 17236 14482 17264 15558
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17052 14476 17184 14482
rect 17052 14470 17132 14476
rect 17132 14418 17184 14424
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 16960 14062 17080 14090
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16960 12986 16988 13874
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17052 12434 17080 14062
rect 17144 13870 17172 14418
rect 17328 14074 17356 15370
rect 17420 15366 17448 17070
rect 17512 16998 17540 18158
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17498 16416 17554 16425
rect 17498 16351 17554 16360
rect 17512 16250 17540 16351
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17604 16114 17632 17750
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17592 15972 17644 15978
rect 17592 15914 17644 15920
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17498 15328 17554 15337
rect 17420 14346 17448 15302
rect 17498 15263 17554 15272
rect 17512 14890 17540 15263
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17604 14226 17632 15914
rect 17420 14198 17632 14226
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17144 13394 17172 13806
rect 17420 13734 17448 14198
rect 17696 13818 17724 18022
rect 17774 17776 17830 17785
rect 17774 17711 17830 17720
rect 17788 17270 17816 17711
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17774 16688 17830 16697
rect 17774 16623 17830 16632
rect 17788 16096 17816 16623
rect 17880 16250 17908 17274
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 18156 16726 18184 17206
rect 18340 17105 18368 18255
rect 18326 17096 18382 17105
rect 18326 17031 18382 17040
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18340 16454 18368 16526
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17868 16108 17920 16114
rect 17788 16068 17868 16096
rect 17868 16050 17920 16056
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17788 15026 17816 15370
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18432 15162 18460 19654
rect 18524 19446 18552 22578
rect 19076 22574 19104 22714
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 18696 22432 18748 22438
rect 18696 22374 18748 22380
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18616 20942 18644 21286
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 18616 20602 18644 20878
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18512 19440 18564 19446
rect 18512 19382 18564 19388
rect 18602 19000 18658 19009
rect 18602 18935 18658 18944
rect 18616 18766 18644 18935
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18524 17270 18552 17478
rect 18512 17264 18564 17270
rect 18512 17206 18564 17212
rect 18616 16697 18644 18566
rect 18602 16688 18658 16697
rect 18512 16652 18564 16658
rect 18602 16623 18658 16632
rect 18512 16594 18564 16600
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17788 14346 17816 14962
rect 18144 14408 18196 14414
rect 18064 14368 18144 14396
rect 17776 14340 17828 14346
rect 18064 14328 18092 14368
rect 18144 14350 18196 14356
rect 17828 14300 18092 14328
rect 17776 14282 17828 14288
rect 17880 14006 17908 14300
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17776 13864 17828 13870
rect 17696 13812 17776 13818
rect 17696 13806 17828 13812
rect 17696 13790 17816 13806
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17420 13530 17448 13670
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17420 12850 17448 13194
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17052 12406 17172 12434
rect 17144 11830 17172 12406
rect 17314 11928 17370 11937
rect 17314 11863 17316 11872
rect 17368 11863 17370 11872
rect 17316 11834 17368 11840
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16868 10062 16896 11086
rect 16960 10810 16988 11494
rect 17052 10810 17080 11630
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16396 9590 16448 9596
rect 16684 9574 16804 9602
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 16120 8560 16172 8566
rect 16120 8502 16172 8508
rect 16132 8430 16160 8502
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16684 8294 16712 9574
rect 16868 9518 16896 9998
rect 17052 9994 17080 10746
rect 17512 10674 17540 13330
rect 17880 13258 17908 13942
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18432 12918 18460 15098
rect 18524 14278 18552 16594
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18616 15910 18644 16390
rect 18708 16114 18736 22374
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 18984 21622 19012 21898
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 18800 19922 18828 20334
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18788 19440 18840 19446
rect 18788 19382 18840 19388
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18800 14793 18828 19382
rect 18892 19174 18920 20878
rect 18984 19990 19012 21422
rect 19076 20602 19104 21422
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 18972 19984 19024 19990
rect 18972 19926 19024 19932
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 19076 19514 19104 19790
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18892 18601 18920 18702
rect 18878 18592 18934 18601
rect 18878 18527 18934 18536
rect 18878 17912 18934 17921
rect 18878 17847 18934 17856
rect 18892 16114 18920 17847
rect 18984 17746 19012 19450
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18972 17740 19024 17746
rect 18972 17682 19024 17688
rect 18970 16688 19026 16697
rect 18970 16623 19026 16632
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18786 14784 18842 14793
rect 18786 14719 18842 14728
rect 18984 14634 19012 16623
rect 18708 14606 19012 14634
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18064 12442 18092 12786
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18602 12744 18658 12753
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17880 11898 17908 12106
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18340 11898 18368 12582
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17040 9988 17092 9994
rect 17040 9930 17092 9936
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 17500 9512 17552 9518
rect 17604 9489 17632 11630
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17880 10742 17908 11018
rect 18432 11014 18460 12718
rect 18602 12679 18658 12688
rect 18616 11694 18644 12679
rect 18708 12170 18736 14606
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18800 12986 18828 13806
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18892 12442 18920 12854
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18892 12170 18920 12378
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18616 11558 18644 11630
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18708 11218 18736 11630
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18892 11150 18920 12106
rect 18984 11354 19012 13194
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17880 9994 17908 10678
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 18892 9722 18920 10202
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18880 9716 18932 9722
rect 18880 9658 18932 9664
rect 17500 9454 17552 9460
rect 17590 9480 17646 9489
rect 16868 9042 16896 9454
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13372 7546 13400 7686
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12084 3534 12112 3674
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 11624 2582 11652 3334
rect 12636 3126 12664 5646
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13464 3670 13492 7686
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 5778 14044 7142
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 15212 4146 15240 7958
rect 15660 7268 15712 7274
rect 15660 7210 15712 7216
rect 15672 5234 15700 7210
rect 16868 5778 16896 8978
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17236 8634 17264 8774
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17512 8090 17540 9454
rect 17590 9415 17646 9424
rect 17604 9178 17632 9415
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18432 8566 18460 9658
rect 18512 9648 18564 9654
rect 18512 9590 18564 9596
rect 18524 9450 18552 9590
rect 19076 9450 19104 19314
rect 19168 16590 19196 24142
rect 19524 23656 19576 23662
rect 19524 23598 19576 23604
rect 19340 23248 19392 23254
rect 19340 23190 19392 23196
rect 19352 22982 19380 23190
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 19260 22137 19288 22374
rect 19246 22128 19302 22137
rect 19444 22098 19472 22578
rect 19246 22063 19302 22072
rect 19432 22092 19484 22098
rect 19536 22094 19564 23598
rect 19628 23322 19656 26200
rect 19800 24200 19852 24206
rect 19800 24142 19852 24148
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19536 22066 19656 22094
rect 19432 22034 19484 22040
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 19260 19514 19288 19926
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19352 19394 19380 21830
rect 19444 21350 19472 22034
rect 19524 22024 19576 22030
rect 19522 21992 19524 22001
rect 19576 21992 19578 22001
rect 19522 21927 19578 21936
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19444 20942 19472 21286
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19444 20602 19472 20878
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19522 20088 19578 20097
rect 19522 20023 19578 20032
rect 19536 19786 19564 20023
rect 19432 19780 19484 19786
rect 19432 19722 19484 19728
rect 19524 19780 19576 19786
rect 19524 19722 19576 19728
rect 19260 19366 19380 19394
rect 19260 18737 19288 19366
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19246 18728 19302 18737
rect 19246 18663 19302 18672
rect 19352 18426 19380 18838
rect 19444 18465 19472 19722
rect 19522 19272 19578 19281
rect 19522 19207 19578 19216
rect 19536 18737 19564 19207
rect 19522 18728 19578 18737
rect 19522 18663 19578 18672
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19430 18456 19486 18465
rect 19340 18420 19392 18426
rect 19430 18391 19486 18400
rect 19340 18362 19392 18368
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19352 17678 19380 18158
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19156 16584 19208 16590
rect 19156 16526 19208 16532
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19338 16144 19394 16153
rect 19338 16079 19394 16088
rect 19156 15428 19208 15434
rect 19156 15370 19208 15376
rect 19168 12617 19196 15370
rect 19352 15366 19380 16079
rect 19444 15570 19472 16526
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19340 15360 19392 15366
rect 19536 15337 19564 18566
rect 19628 17746 19656 22066
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19720 21010 19748 21286
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19812 20058 19840 24142
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 20088 23186 20116 23462
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19892 22228 19944 22234
rect 19892 22170 19944 22176
rect 19904 21690 19932 22170
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 19800 20052 19852 20058
rect 19800 19994 19852 20000
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19720 19310 19748 19790
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19720 18834 19748 19246
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19812 18358 19840 18566
rect 19708 18352 19760 18358
rect 19708 18294 19760 18300
rect 19800 18352 19852 18358
rect 19800 18294 19852 18300
rect 19720 18086 19748 18294
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19614 17232 19670 17241
rect 19614 17167 19670 17176
rect 19800 17196 19852 17202
rect 19628 15638 19656 17167
rect 19800 17138 19852 17144
rect 19812 16794 19840 17138
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19720 16250 19748 16730
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19616 15632 19668 15638
rect 19616 15574 19668 15580
rect 19340 15302 19392 15308
rect 19522 15328 19578 15337
rect 19522 15263 19578 15272
rect 19536 15144 19564 15263
rect 19352 15116 19564 15144
rect 19352 15042 19380 15116
rect 19260 15014 19380 15042
rect 19432 15020 19484 15026
rect 19260 14822 19288 15014
rect 19432 14962 19484 14968
rect 19338 14920 19394 14929
rect 19338 14855 19394 14864
rect 19352 14822 19380 14855
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19248 13796 19300 13802
rect 19248 13738 19300 13744
rect 19154 12608 19210 12617
rect 19154 12543 19210 12552
rect 19260 12434 19288 13738
rect 19168 12406 19288 12434
rect 19168 11257 19196 12406
rect 19154 11248 19210 11257
rect 19154 11183 19210 11192
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 18512 9444 18564 9450
rect 18512 9386 18564 9392
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 18524 8838 18552 9386
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 12084 800 12112 2450
rect 12452 2446 12480 2858
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 14752 800 14780 2450
rect 15028 2446 15056 3878
rect 15488 3126 15516 5102
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 17052 3058 17080 5510
rect 17420 4826 17448 5578
rect 17512 5234 17540 7142
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18524 5710 18552 8774
rect 19260 7954 19288 9930
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19352 6866 19380 14758
rect 19444 12374 19472 14962
rect 19616 14952 19668 14958
rect 19616 14894 19668 14900
rect 19628 14414 19656 14894
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19904 13977 19932 19654
rect 19996 14890 20024 23054
rect 20088 22710 20116 23122
rect 20076 22704 20128 22710
rect 20076 22646 20128 22652
rect 20076 22568 20128 22574
rect 20076 22510 20128 22516
rect 20088 22234 20116 22510
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 20166 21992 20222 22001
rect 20272 21962 20300 26200
rect 20718 24848 20774 24857
rect 20718 24783 20774 24792
rect 20534 24440 20590 24449
rect 20534 24375 20590 24384
rect 20352 24064 20404 24070
rect 20352 24006 20404 24012
rect 20364 22030 20392 24006
rect 20444 23520 20496 23526
rect 20444 23462 20496 23468
rect 20456 22574 20484 23462
rect 20444 22568 20496 22574
rect 20444 22510 20496 22516
rect 20548 22250 20576 24375
rect 20628 22976 20680 22982
rect 20628 22918 20680 22924
rect 20640 22273 20668 22918
rect 20456 22222 20576 22250
rect 20626 22264 20682 22273
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20166 21927 20222 21936
rect 20260 21956 20312 21962
rect 20180 21321 20208 21927
rect 20260 21898 20312 21904
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20166 21312 20222 21321
rect 20166 21247 20222 21256
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 20088 18222 20116 18634
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 20076 17060 20128 17066
rect 20076 17002 20128 17008
rect 20088 16969 20116 17002
rect 20168 16992 20220 16998
rect 20074 16960 20130 16969
rect 20168 16934 20220 16940
rect 20074 16895 20130 16904
rect 20180 16833 20208 16934
rect 20166 16824 20222 16833
rect 20166 16759 20222 16768
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20088 15706 20116 16390
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 20272 15586 20300 21354
rect 20456 19786 20484 22222
rect 20626 22199 20682 22208
rect 20732 22148 20760 24783
rect 20916 24274 20944 26200
rect 21178 24712 21234 24721
rect 21178 24647 21234 24656
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 21192 23798 21220 24647
rect 21560 24274 21588 26200
rect 21638 24304 21694 24313
rect 21548 24268 21600 24274
rect 21638 24239 21694 24248
rect 21548 24210 21600 24216
rect 21180 23792 21232 23798
rect 21180 23734 21232 23740
rect 20904 23724 20956 23730
rect 20904 23666 20956 23672
rect 20640 22120 20760 22148
rect 20640 22094 20668 22120
rect 20548 22066 20668 22094
rect 20444 19780 20496 19786
rect 20444 19722 20496 19728
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20364 16658 20392 17682
rect 20548 17649 20576 22066
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20640 19310 20668 20334
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20720 18896 20772 18902
rect 20720 18838 20772 18844
rect 20732 18426 20760 18838
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20824 18222 20852 18566
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20534 17640 20590 17649
rect 20732 17610 20760 18090
rect 20534 17575 20590 17584
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20456 16114 20484 17478
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20640 16998 20668 17138
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20732 16658 20760 16934
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20180 15558 20300 15586
rect 20628 15564 20680 15570
rect 20180 15502 20208 15558
rect 20628 15506 20680 15512
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20260 15088 20312 15094
rect 20260 15030 20312 15036
rect 20272 14958 20300 15030
rect 20640 15026 20668 15506
rect 20732 15094 20760 16390
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20088 14074 20116 14418
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 19890 13968 19946 13977
rect 19890 13903 19946 13912
rect 20076 13388 20128 13394
rect 20076 13330 20128 13336
rect 20088 12782 20116 13330
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 19614 12336 19670 12345
rect 20088 12306 20116 12718
rect 19614 12271 19616 12280
rect 19668 12271 19670 12280
rect 20076 12300 20128 12306
rect 19616 12242 19668 12248
rect 20076 12242 20128 12248
rect 19628 11626 19656 12242
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19720 11082 19748 11630
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19720 10606 19748 11018
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19720 10130 19748 10542
rect 20180 10266 20208 14418
rect 20720 14408 20772 14414
rect 20718 14376 20720 14385
rect 20772 14376 20774 14385
rect 20718 14311 20774 14320
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20364 13870 20392 14010
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20364 12170 20392 13466
rect 20352 12164 20404 12170
rect 20352 12106 20404 12112
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20272 10266 20300 10678
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 20168 9988 20220 9994
rect 20272 9976 20300 10202
rect 20220 9948 20300 9976
rect 20168 9930 20220 9936
rect 20180 9382 20208 9930
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20364 8430 20392 12106
rect 20456 8498 20484 13874
rect 20548 10470 20576 14214
rect 20628 13796 20680 13802
rect 20628 13738 20680 13744
rect 20640 12424 20668 13738
rect 20720 12436 20772 12442
rect 20640 12396 20720 12424
rect 20720 12378 20772 12384
rect 20824 12306 20852 18158
rect 20916 14006 20944 23666
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 21364 23044 21416 23050
rect 21364 22986 21416 22992
rect 21088 22976 21140 22982
rect 21088 22918 21140 22924
rect 21100 20806 21128 22918
rect 21376 22710 21404 22986
rect 21468 22778 21496 23258
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21364 22704 21416 22710
rect 21364 22646 21416 22652
rect 21376 21690 21404 22646
rect 21364 21684 21416 21690
rect 21416 21644 21496 21672
rect 21364 21626 21416 21632
rect 21364 21072 21416 21078
rect 21364 21014 21416 21020
rect 21088 20800 21140 20806
rect 21088 20742 21140 20748
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21192 19922 21220 20742
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 21284 19334 21312 19994
rect 21192 19306 21312 19334
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 21008 18426 21036 19110
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 21088 18352 21140 18358
rect 21088 18294 21140 18300
rect 21100 18057 21128 18294
rect 21086 18048 21142 18057
rect 21086 17983 21142 17992
rect 21192 17882 21220 19306
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 21284 17592 21312 17818
rect 21376 17728 21404 21014
rect 21468 21010 21496 21644
rect 21456 21004 21508 21010
rect 21456 20946 21508 20952
rect 21468 20534 21496 20946
rect 21456 20528 21508 20534
rect 21456 20470 21508 20476
rect 21468 19802 21496 20470
rect 21468 19786 21588 19802
rect 21468 19780 21600 19786
rect 21468 19774 21548 19780
rect 21548 19722 21600 19728
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21468 18834 21496 19654
rect 21560 19446 21588 19722
rect 21548 19440 21600 19446
rect 21548 19382 21600 19388
rect 21456 18828 21508 18834
rect 21456 18770 21508 18776
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21376 17700 21496 17728
rect 21100 17564 21312 17592
rect 21362 17640 21418 17649
rect 21362 17575 21418 17584
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 21008 16794 21036 17478
rect 21100 17202 21128 17564
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21008 16522 21036 16730
rect 21088 16720 21140 16726
rect 21284 16697 21312 17138
rect 21088 16662 21140 16668
rect 21270 16688 21326 16697
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 21008 15570 21036 16458
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20996 15088 21048 15094
rect 20996 15030 21048 15036
rect 21008 14822 21036 15030
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 21008 13870 21036 14010
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 21100 12889 21128 16662
rect 21270 16623 21326 16632
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 21192 16250 21220 16458
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21376 15609 21404 17575
rect 21468 16726 21496 17700
rect 21560 16998 21588 18770
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21456 16720 21508 16726
rect 21456 16662 21508 16668
rect 21454 16416 21510 16425
rect 21454 16351 21510 16360
rect 21468 16114 21496 16351
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21362 15600 21418 15609
rect 21362 15535 21418 15544
rect 21560 14550 21588 16934
rect 21652 16046 21680 24239
rect 22006 24032 22062 24041
rect 22006 23967 22062 23976
rect 21824 23792 21876 23798
rect 21824 23734 21876 23740
rect 21836 23186 21864 23734
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21916 23112 21968 23118
rect 21916 23054 21968 23060
rect 21928 22642 21956 23054
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 21928 22438 21956 22578
rect 21916 22432 21968 22438
rect 21916 22374 21968 22380
rect 21928 22098 21956 22374
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 22020 22030 22048 23967
rect 22204 23225 22232 26200
rect 22848 25906 22876 26200
rect 22836 25900 22888 25906
rect 22836 25842 22888 25848
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23296 23792 23348 23798
rect 23296 23734 23348 23740
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22190 23216 22246 23225
rect 22190 23151 22246 23160
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22204 20482 22232 21830
rect 22296 20942 22324 23462
rect 22388 23322 22416 23598
rect 22376 23316 22428 23322
rect 22376 23258 22428 23264
rect 22388 22710 22416 23258
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22848 22642 22876 23598
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23308 23322 23336 23734
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23308 23050 23336 23258
rect 23296 23044 23348 23050
rect 23296 22986 23348 22992
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22652 22568 22704 22574
rect 22652 22510 22704 22516
rect 22664 22166 22692 22510
rect 22652 22160 22704 22166
rect 22652 22102 22704 22108
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22388 21894 22416 21966
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22388 21078 22416 21830
rect 22848 21690 22876 22578
rect 23492 22438 23520 26200
rect 24032 24200 24084 24206
rect 24032 24142 24084 24148
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23572 23316 23624 23322
rect 23572 23258 23624 23264
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23204 22160 23256 22166
rect 23204 22102 23256 22108
rect 22926 21856 22982 21865
rect 22926 21791 22982 21800
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22940 21622 22968 21791
rect 23216 21729 23244 22102
rect 23202 21720 23258 21729
rect 23202 21655 23258 21664
rect 22928 21616 22980 21622
rect 22928 21558 22980 21564
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22376 21072 22428 21078
rect 22376 21014 22428 21020
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22020 20466 22232 20482
rect 22008 20460 22232 20466
rect 22060 20454 22232 20460
rect 22008 20402 22060 20408
rect 21824 19440 21876 19446
rect 21824 19382 21876 19388
rect 21836 19242 21864 19382
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 21824 19236 21876 19242
rect 21824 19178 21876 19184
rect 21732 17876 21784 17882
rect 21732 17818 21784 17824
rect 21744 17134 21772 17818
rect 21836 17542 21864 19178
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21928 17354 21956 19314
rect 22112 19224 22140 20454
rect 22296 19854 22324 20878
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22560 20800 22612 20806
rect 22560 20742 22612 20748
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22480 20602 22508 20742
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22572 20330 22600 20742
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22664 19446 22692 20742
rect 23400 20466 23428 21490
rect 23584 21146 23612 23258
rect 23768 23254 23796 23462
rect 23756 23248 23808 23254
rect 23756 23190 23808 23196
rect 23940 22976 23992 22982
rect 24044 22953 24072 24142
rect 24136 23089 24164 26200
rect 24308 24064 24360 24070
rect 24308 24006 24360 24012
rect 24122 23080 24178 23089
rect 24122 23015 24178 23024
rect 23940 22918 23992 22924
rect 24030 22944 24086 22953
rect 23664 22704 23716 22710
rect 23664 22646 23716 22652
rect 23676 22030 23704 22646
rect 23952 22574 23980 22918
rect 24030 22879 24086 22888
rect 23940 22568 23992 22574
rect 23940 22510 23992 22516
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23952 21622 23980 22374
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23572 21004 23624 21010
rect 23572 20946 23624 20952
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22836 19984 22888 19990
rect 22836 19926 22888 19932
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22192 19236 22244 19242
rect 22112 19196 22192 19224
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22020 18970 22048 19110
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 22112 18630 22140 19196
rect 22192 19178 22244 19184
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22572 18766 22600 19110
rect 22664 18970 22692 19246
rect 22652 18964 22704 18970
rect 22652 18906 22704 18912
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22006 18456 22062 18465
rect 22006 18391 22062 18400
rect 22020 18290 22048 18391
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 21836 17326 21956 17354
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21652 15706 21680 15982
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21548 14544 21600 14550
rect 21548 14486 21600 14492
rect 21560 14278 21588 14486
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21192 12986 21220 14010
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 21284 12986 21312 13126
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21086 12880 21142 12889
rect 21086 12815 21142 12824
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20916 11898 20944 12582
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 21468 11558 21496 12718
rect 21744 12714 21772 16934
rect 21836 14414 21864 17326
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21928 14890 21956 15302
rect 22020 15026 22048 17614
rect 22112 15609 22140 18566
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22480 18057 22508 18158
rect 22466 18048 22522 18057
rect 22466 17983 22522 17992
rect 22480 17338 22508 17983
rect 22560 17604 22612 17610
rect 22560 17546 22612 17552
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22192 17060 22244 17066
rect 22192 17002 22244 17008
rect 22098 15600 22154 15609
rect 22098 15535 22154 15544
rect 22112 15162 22140 15535
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22204 15094 22232 17002
rect 22480 16776 22508 17274
rect 22572 17270 22600 17546
rect 22560 17264 22612 17270
rect 22560 17206 22612 17212
rect 22756 17218 22784 19722
rect 22848 18086 22876 19926
rect 23584 19786 23612 20946
rect 23676 20806 23704 21082
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23756 20596 23808 20602
rect 23756 20538 23808 20544
rect 23768 19854 23796 20538
rect 23860 19922 23888 20946
rect 24124 20936 24176 20942
rect 24124 20878 24176 20884
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23572 19780 23624 19786
rect 23572 19722 23624 19728
rect 23296 19712 23348 19718
rect 23296 19654 23348 19660
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23308 19514 23336 19654
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23388 19304 23440 19310
rect 23388 19246 23440 19252
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23400 18850 23428 19246
rect 23308 18822 23428 18850
rect 22926 18456 22982 18465
rect 22926 18391 22982 18400
rect 22940 18222 22968 18391
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 22836 18080 22888 18086
rect 22836 18022 22888 18028
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22756 17190 22876 17218
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22572 16998 22600 17070
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22480 16748 22692 16776
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22296 15745 22324 15982
rect 22282 15736 22338 15745
rect 22282 15671 22338 15680
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21836 14006 21864 14350
rect 21928 14346 21956 14826
rect 22020 14482 22048 14962
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 22020 13297 22048 14214
rect 22204 13530 22232 15030
rect 22388 14090 22416 16390
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22296 14062 22416 14090
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22006 13288 22062 13297
rect 22006 13223 22062 13232
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 21732 12708 21784 12714
rect 21732 12650 21784 12656
rect 22020 12646 22048 12922
rect 22008 12640 22060 12646
rect 21836 12600 22008 12628
rect 21836 12170 21864 12600
rect 22008 12582 22060 12588
rect 22204 12628 22232 13330
rect 22296 12918 22324 14062
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22388 13258 22416 13874
rect 22376 13252 22428 13258
rect 22376 13194 22428 13200
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22480 12782 22508 15846
rect 22572 15502 22600 16594
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22572 15162 22600 15438
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22664 15042 22692 16748
rect 22572 15014 22692 15042
rect 22572 13938 22600 15014
rect 22848 14278 22876 17190
rect 23308 17082 23336 18822
rect 23584 18766 23612 19450
rect 23676 18834 23704 19654
rect 23756 19168 23808 19174
rect 23756 19110 23808 19116
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23768 18766 23796 19110
rect 23572 18760 23624 18766
rect 23386 18728 23442 18737
rect 23756 18760 23808 18766
rect 23572 18702 23624 18708
rect 23676 18708 23756 18714
rect 23676 18702 23808 18708
rect 23386 18663 23442 18672
rect 23676 18686 23796 18702
rect 23400 18630 23428 18663
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23492 18358 23520 18566
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23676 17678 23704 18686
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23754 17912 23810 17921
rect 23754 17847 23756 17856
rect 23808 17847 23810 17856
rect 23756 17818 23808 17824
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23768 17270 23796 17682
rect 23756 17264 23808 17270
rect 23756 17206 23808 17212
rect 23756 17128 23808 17134
rect 23308 17054 23428 17082
rect 23860 17116 23888 18566
rect 23952 17241 23980 20742
rect 23938 17232 23994 17241
rect 23938 17167 23994 17176
rect 23808 17088 23888 17116
rect 23756 17070 23808 17076
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23308 16590 23336 16934
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23400 15978 23428 17054
rect 23768 16794 23796 17070
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23676 16114 23704 16526
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23388 15972 23440 15978
rect 23388 15914 23440 15920
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23664 15700 23716 15706
rect 23664 15642 23716 15648
rect 22928 15632 22980 15638
rect 22926 15600 22928 15609
rect 22980 15600 22982 15609
rect 22926 15535 22982 15544
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22572 13530 22600 13874
rect 22744 13796 22796 13802
rect 22744 13738 22796 13744
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22756 13274 22784 13738
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22848 13462 22876 13670
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23308 13530 23336 15438
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23400 15026 23428 15302
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23400 14890 23428 14962
rect 23388 14884 23440 14890
rect 23388 14826 23440 14832
rect 23572 14544 23624 14550
rect 23572 14486 23624 14492
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 22836 13456 22888 13462
rect 23400 13410 23428 14214
rect 22836 13398 22888 13404
rect 23216 13382 23428 13410
rect 23480 13388 23532 13394
rect 23020 13320 23072 13326
rect 22756 13246 22876 13274
rect 23020 13262 23072 13268
rect 23110 13288 23166 13297
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22284 12640 22336 12646
rect 22204 12600 22284 12628
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 21928 12306 21956 12378
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 22204 12238 22232 12600
rect 22284 12582 22336 12588
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 21824 12164 21876 12170
rect 21824 12106 21876 12112
rect 21836 11830 21864 12106
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 21836 11558 21864 11766
rect 22204 11694 22232 12174
rect 22756 11830 22784 12922
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 21192 9926 21220 11018
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21376 10538 21404 10950
rect 21468 10810 21496 11494
rect 21836 11218 21864 11494
rect 21824 11212 21876 11218
rect 21824 11154 21876 11160
rect 21836 11082 21864 11154
rect 21824 11076 21876 11082
rect 21824 11018 21876 11024
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21364 10532 21416 10538
rect 21364 10474 21416 10480
rect 21836 10470 21864 11018
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21836 10266 21864 10406
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21836 10062 21864 10202
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 21192 9518 21220 9862
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 22204 7410 22232 11630
rect 22848 11354 22876 13246
rect 23032 12850 23060 13262
rect 23110 13223 23112 13232
rect 23164 13223 23166 13232
rect 23112 13194 23164 13200
rect 23216 12986 23244 13382
rect 23480 13330 23532 13336
rect 23492 12986 23520 13330
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23584 12918 23612 14486
rect 23572 12912 23624 12918
rect 23572 12854 23624 12860
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 23032 12646 23060 12786
rect 23020 12640 23072 12646
rect 23020 12582 23072 12588
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23020 12164 23072 12170
rect 23020 12106 23072 12112
rect 23032 11812 23060 12106
rect 23112 11824 23164 11830
rect 23032 11784 23112 11812
rect 23112 11766 23164 11772
rect 23124 11558 23152 11766
rect 23676 11694 23704 15642
rect 23768 13802 23796 16594
rect 23848 16448 23900 16454
rect 24136 16425 24164 20878
rect 24214 20768 24270 20777
rect 24214 20703 24270 20712
rect 24228 20466 24256 20703
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 23848 16390 23900 16396
rect 24122 16416 24178 16425
rect 23860 16114 23888 16390
rect 24122 16351 24178 16360
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23940 15428 23992 15434
rect 23940 15370 23992 15376
rect 23952 15026 23980 15370
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23860 14346 23888 14758
rect 23952 14482 23980 14962
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23848 14340 23900 14346
rect 23848 14282 23900 14288
rect 23756 13796 23808 13802
rect 23756 13738 23808 13744
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23768 13258 23796 13330
rect 23756 13252 23808 13258
rect 23756 13194 23808 13200
rect 23860 12918 23888 14282
rect 24044 13870 24072 15982
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 23952 13258 23980 13466
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 23848 12912 23900 12918
rect 23848 12854 23900 12860
rect 23860 12782 23888 12854
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 24044 12102 24072 13806
rect 24136 13530 24164 13874
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 24044 11898 24072 12038
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23112 11552 23164 11558
rect 23756 11552 23808 11558
rect 23112 11494 23164 11500
rect 23400 11512 23756 11540
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22848 10606 22876 11290
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23400 9994 23428 11512
rect 23756 11494 23808 11500
rect 23572 10056 23624 10062
rect 23572 9998 23624 10004
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23400 7750 23428 9454
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17420 2990 17448 4762
rect 17696 4486 17724 5102
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17696 3126 17724 4422
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17880 3058 17908 4966
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 20548 3058 20576 4966
rect 20732 3466 20760 6802
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 21744 5846 21772 6734
rect 22480 5914 22508 7278
rect 22848 6458 22876 7686
rect 23584 7410 23612 9998
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 23768 6866 23796 9522
rect 24320 9081 24348 24006
rect 24780 23497 24808 26200
rect 24964 24206 24992 26302
rect 25410 26200 25466 26302
rect 26054 26330 26110 27000
rect 26698 26330 26754 27000
rect 26054 26302 26188 26330
rect 26054 26200 26110 26302
rect 25596 25832 25648 25838
rect 25596 25774 25648 25780
rect 25608 25022 25636 25774
rect 26160 25022 26188 26302
rect 26698 26302 27292 26330
rect 26698 26200 26754 26302
rect 26792 25900 26844 25906
rect 26792 25842 26844 25848
rect 25596 25016 25648 25022
rect 25596 24958 25648 24964
rect 26148 25016 26200 25022
rect 26148 24958 26200 24964
rect 25044 24812 25096 24818
rect 25044 24754 25096 24760
rect 25056 24274 25084 24754
rect 26240 24744 26292 24750
rect 26240 24686 26292 24692
rect 25688 24608 25740 24614
rect 25688 24550 25740 24556
rect 25700 24410 25728 24550
rect 25688 24404 25740 24410
rect 25688 24346 25740 24352
rect 25872 24404 25924 24410
rect 25872 24346 25924 24352
rect 25044 24268 25096 24274
rect 25044 24210 25096 24216
rect 25320 24268 25372 24274
rect 25320 24210 25372 24216
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 25332 24138 25360 24210
rect 25884 24206 25912 24346
rect 26252 24206 26280 24686
rect 26516 24336 26568 24342
rect 26516 24278 26568 24284
rect 25872 24200 25924 24206
rect 25872 24142 25924 24148
rect 25964 24200 26016 24206
rect 25964 24142 26016 24148
rect 26240 24200 26292 24206
rect 26240 24142 26292 24148
rect 26424 24200 26476 24206
rect 26424 24142 26476 24148
rect 25320 24132 25372 24138
rect 25320 24074 25372 24080
rect 25504 24132 25556 24138
rect 25504 24074 25556 24080
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 24964 23866 24992 24006
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25148 23662 25176 24006
rect 25412 23792 25464 23798
rect 25516 23780 25544 24074
rect 25464 23752 25544 23780
rect 25412 23734 25464 23740
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 25780 23656 25832 23662
rect 25780 23598 25832 23604
rect 24872 23526 24900 23598
rect 24860 23520 24912 23526
rect 24766 23488 24822 23497
rect 24860 23462 24912 23468
rect 24766 23423 24822 23432
rect 25688 23248 25740 23254
rect 25688 23190 25740 23196
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 24400 22704 24452 22710
rect 24400 22646 24452 22652
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24412 21729 24440 22646
rect 24584 22228 24636 22234
rect 24584 22170 24636 22176
rect 24398 21720 24454 21729
rect 24398 21655 24454 21664
rect 24412 21622 24440 21655
rect 24400 21616 24452 21622
rect 24400 21558 24452 21564
rect 24412 20516 24440 21558
rect 24492 20528 24544 20534
rect 24412 20488 24492 20516
rect 24492 20470 24544 20476
rect 24596 20058 24624 22170
rect 24780 22030 24808 22646
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 25056 21865 25084 23054
rect 25148 22778 25176 23122
rect 25700 22778 25728 23190
rect 25792 22778 25820 23598
rect 25976 22982 26004 24142
rect 26436 23866 26464 24142
rect 26528 23905 26556 24278
rect 26514 23896 26570 23905
rect 26424 23860 26476 23866
rect 26514 23831 26570 23840
rect 26424 23802 26476 23808
rect 26516 23792 26568 23798
rect 26516 23734 26568 23740
rect 25964 22976 26016 22982
rect 25964 22918 26016 22924
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 25688 22772 25740 22778
rect 25688 22714 25740 22720
rect 25780 22772 25832 22778
rect 25780 22714 25832 22720
rect 25136 22568 25188 22574
rect 25136 22510 25188 22516
rect 25148 22166 25176 22510
rect 25700 22438 25728 22714
rect 25976 22574 26004 22918
rect 25964 22568 26016 22574
rect 25884 22528 25964 22556
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25136 22160 25188 22166
rect 25136 22102 25188 22108
rect 25042 21856 25098 21865
rect 25042 21791 25098 21800
rect 25056 21690 25084 21791
rect 25044 21684 25096 21690
rect 25044 21626 25096 21632
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 24688 20398 24716 21422
rect 24768 21412 24820 21418
rect 24768 21354 24820 21360
rect 24780 20942 24808 21354
rect 25332 21350 25360 22374
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 25700 21010 25728 21966
rect 25884 21894 25912 22528
rect 25964 22510 26016 22516
rect 26424 22568 26476 22574
rect 26424 22510 26476 22516
rect 26240 22432 26292 22438
rect 26240 22374 26292 22380
rect 25872 21888 25924 21894
rect 25872 21830 25924 21836
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25976 21690 26004 21830
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 26252 21026 26280 22374
rect 26332 21956 26384 21962
rect 26332 21898 26384 21904
rect 26344 21690 26372 21898
rect 26332 21684 26384 21690
rect 26332 21626 26384 21632
rect 25688 21004 25740 21010
rect 25688 20946 25740 20952
rect 26056 21004 26108 21010
rect 26056 20946 26108 20952
rect 26160 20998 26280 21026
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 25700 20777 25728 20946
rect 25872 20936 25924 20942
rect 25872 20878 25924 20884
rect 25686 20768 25742 20777
rect 25686 20703 25742 20712
rect 25884 20466 25912 20878
rect 26068 20602 26096 20946
rect 26056 20596 26108 20602
rect 26056 20538 26108 20544
rect 25872 20460 25924 20466
rect 25872 20402 25924 20408
rect 24676 20392 24728 20398
rect 25964 20392 26016 20398
rect 24676 20334 24728 20340
rect 24766 20360 24822 20369
rect 25964 20334 26016 20340
rect 24766 20295 24822 20304
rect 24584 20052 24636 20058
rect 24584 19994 24636 20000
rect 24780 19854 24808 20295
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24398 18592 24454 18601
rect 24398 18527 24454 18536
rect 24412 18170 24440 18527
rect 24412 18154 24532 18170
rect 24412 18148 24544 18154
rect 24412 18142 24492 18148
rect 24492 18090 24544 18096
rect 24400 17536 24452 17542
rect 24400 17478 24452 17484
rect 24412 17338 24440 17478
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24504 17202 24532 18090
rect 24676 18080 24728 18086
rect 24676 18022 24728 18028
rect 24688 17746 24716 18022
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24688 17202 24716 17682
rect 24872 17354 24900 19246
rect 24872 17326 24992 17354
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24676 17196 24728 17202
rect 24728 17156 24900 17184
rect 24676 17138 24728 17144
rect 24504 16590 24532 17138
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24504 16182 24532 16526
rect 24596 16454 24624 16594
rect 24584 16448 24636 16454
rect 24584 16390 24636 16396
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24596 16182 24624 16390
rect 24492 16176 24544 16182
rect 24492 16118 24544 16124
rect 24584 16176 24636 16182
rect 24584 16118 24636 16124
rect 24596 15706 24624 16118
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24584 14272 24636 14278
rect 24584 14214 24636 14220
rect 24596 14006 24624 14214
rect 24584 14000 24636 14006
rect 24584 13942 24636 13948
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24400 12708 24452 12714
rect 24400 12650 24452 12656
rect 24412 12102 24440 12650
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24412 11626 24440 12038
rect 24400 11620 24452 11626
rect 24400 11562 24452 11568
rect 24596 9654 24624 13670
rect 24688 13394 24716 16390
rect 24872 16114 24900 17156
rect 24964 16250 24992 17326
rect 25056 16590 25084 19654
rect 25240 19174 25268 19858
rect 25504 19440 25556 19446
rect 25504 19382 25556 19388
rect 25320 19236 25372 19242
rect 25320 19178 25372 19184
rect 25228 19168 25280 19174
rect 25228 19110 25280 19116
rect 25136 18896 25188 18902
rect 25136 18838 25188 18844
rect 25148 18766 25176 18838
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25148 18358 25176 18702
rect 25136 18352 25188 18358
rect 25136 18294 25188 18300
rect 25240 18222 25268 19110
rect 25332 18358 25360 19178
rect 25410 18728 25466 18737
rect 25410 18663 25466 18672
rect 25320 18352 25372 18358
rect 25320 18294 25372 18300
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 25148 16726 25176 17546
rect 25424 17082 25452 18663
rect 25240 17054 25452 17082
rect 25136 16720 25188 16726
rect 25136 16662 25188 16668
rect 25240 16658 25268 17054
rect 25320 16992 25372 16998
rect 25320 16934 25372 16940
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25332 16522 25360 16934
rect 25516 16522 25544 19382
rect 25700 18970 25728 20198
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25792 19310 25820 19790
rect 25872 19712 25924 19718
rect 25872 19654 25924 19660
rect 25884 19514 25912 19654
rect 25872 19508 25924 19514
rect 25872 19450 25924 19456
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25792 18834 25820 19246
rect 25780 18828 25832 18834
rect 25780 18770 25832 18776
rect 25792 17746 25820 18770
rect 25976 18698 26004 20334
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 26068 18358 26096 20538
rect 26160 20534 26188 20998
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26148 20528 26200 20534
rect 26148 20470 26200 20476
rect 26148 19780 26200 19786
rect 26148 19722 26200 19728
rect 26160 18970 26188 19722
rect 26252 19514 26280 20810
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26148 18964 26200 18970
rect 26148 18906 26200 18912
rect 26238 18864 26294 18873
rect 26238 18799 26240 18808
rect 26292 18799 26294 18808
rect 26240 18770 26292 18776
rect 26056 18352 26108 18358
rect 26056 18294 26108 18300
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25962 17232 26018 17241
rect 25962 17167 26018 17176
rect 25976 16998 26004 17167
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 25686 16688 25742 16697
rect 25976 16658 26004 16934
rect 25686 16623 25742 16632
rect 25780 16652 25832 16658
rect 25320 16516 25372 16522
rect 25320 16458 25372 16464
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 24964 15162 24992 16186
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 25148 14346 25176 16390
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25136 14340 25188 14346
rect 25136 14282 25188 14288
rect 25148 14006 25176 14282
rect 25136 14000 25188 14006
rect 25056 13960 25136 13988
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 25056 12345 25084 13960
rect 25136 13942 25188 13948
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 25042 12336 25098 12345
rect 25042 12271 25098 12280
rect 25148 11558 25176 13806
rect 25240 13297 25268 15302
rect 25332 14822 25360 16458
rect 25700 16454 25728 16623
rect 25780 16594 25832 16600
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 25688 16448 25740 16454
rect 25688 16390 25740 16396
rect 25792 15570 25820 16594
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25596 15360 25648 15366
rect 25594 15328 25596 15337
rect 25648 15328 25650 15337
rect 25594 15263 25650 15272
rect 25320 14816 25372 14822
rect 25320 14758 25372 14764
rect 25332 14278 25360 14758
rect 25792 14550 25820 15506
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 26160 15366 26188 15438
rect 26148 15360 26200 15366
rect 26148 15302 26200 15308
rect 25780 14544 25832 14550
rect 25780 14486 25832 14492
rect 25596 14476 25648 14482
rect 25596 14418 25648 14424
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 25332 13938 25360 14214
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25226 13288 25282 13297
rect 25226 13223 25282 13232
rect 25608 12442 25636 14418
rect 26160 14346 26188 15302
rect 26148 14340 26200 14346
rect 26148 14282 26200 14288
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25792 14074 25820 14214
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 24584 9648 24636 9654
rect 24584 9590 24636 9596
rect 24306 9072 24362 9081
rect 24306 9007 24362 9016
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 23952 7002 23980 7482
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 22756 5778 22784 6054
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 20904 5704 20956 5710
rect 20904 5646 20956 5652
rect 20916 4826 20944 5646
rect 23400 5642 23428 6598
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 25504 5636 25556 5642
rect 25504 5578 25556 5584
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21376 5234 21404 5510
rect 22204 5234 22232 5578
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 17420 800 17448 2450
rect 17512 2446 17540 2790
rect 20088 2446 20116 2790
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20180 1170 20208 2450
rect 22020 2446 22048 2790
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 25516 2650 25544 5578
rect 25964 5024 26016 5030
rect 25964 4966 26016 4972
rect 25976 4554 26004 4966
rect 26436 4554 26464 22510
rect 26528 22438 26556 23734
rect 26608 23520 26660 23526
rect 26608 23462 26660 23468
rect 26620 22642 26648 23462
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 26516 22432 26568 22438
rect 26516 22374 26568 22380
rect 26528 21962 26556 22374
rect 26804 22098 26832 25842
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 26792 22092 26844 22098
rect 26792 22034 26844 22040
rect 26516 21956 26568 21962
rect 26516 21898 26568 21904
rect 26528 21729 26556 21898
rect 26514 21720 26570 21729
rect 26514 21655 26570 21664
rect 26528 20856 26556 21655
rect 26896 21554 26924 25638
rect 27264 24426 27292 26302
rect 27342 26200 27398 27000
rect 27986 26330 28042 27000
rect 27986 26302 28304 26330
rect 27986 26200 28042 26302
rect 27356 24750 27384 26200
rect 28276 25158 28304 26302
rect 28630 26200 28686 27000
rect 29274 26200 29330 27000
rect 29918 26330 29974 27000
rect 29918 26302 30144 26330
rect 29918 26200 29974 26302
rect 27620 25152 27672 25158
rect 27620 25094 27672 25100
rect 28264 25152 28316 25158
rect 28264 25094 28316 25100
rect 27344 24744 27396 24750
rect 27344 24686 27396 24692
rect 27632 24614 27660 25094
rect 28448 25084 28500 25090
rect 28448 25026 28500 25032
rect 27620 24608 27672 24614
rect 27620 24550 27672 24556
rect 27264 24398 27660 24426
rect 27632 24138 27660 24398
rect 27896 24336 27948 24342
rect 27896 24278 27948 24284
rect 27804 24268 27856 24274
rect 27804 24210 27856 24216
rect 27816 24154 27844 24210
rect 27436 24132 27488 24138
rect 27436 24074 27488 24080
rect 27528 24132 27580 24138
rect 27528 24074 27580 24080
rect 27620 24132 27672 24138
rect 27620 24074 27672 24080
rect 27724 24126 27844 24154
rect 27068 23792 27120 23798
rect 27068 23734 27120 23740
rect 27080 22930 27108 23734
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 27172 23186 27200 23598
rect 27252 23520 27304 23526
rect 27252 23462 27304 23468
rect 27160 23180 27212 23186
rect 27160 23122 27212 23128
rect 27080 22902 27200 22930
rect 27172 22094 27200 22902
rect 27264 22574 27292 23462
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27252 22568 27304 22574
rect 27252 22510 27304 22516
rect 27356 22273 27384 22578
rect 27448 22506 27476 24074
rect 27436 22500 27488 22506
rect 27436 22442 27488 22448
rect 27342 22264 27398 22273
rect 27342 22199 27398 22208
rect 27448 22166 27476 22442
rect 27436 22160 27488 22166
rect 27436 22102 27488 22108
rect 27172 22066 27292 22094
rect 26884 21548 26936 21554
rect 26884 21490 26936 21496
rect 26608 21480 26660 21486
rect 26608 21422 26660 21428
rect 26620 21321 26648 21422
rect 26606 21312 26662 21321
rect 26606 21247 26662 21256
rect 26608 20868 26660 20874
rect 26528 20828 26608 20856
rect 26528 20262 26556 20828
rect 26608 20810 26660 20816
rect 26516 20256 26568 20262
rect 26568 20216 26648 20244
rect 26516 20198 26568 20204
rect 26620 19786 26648 20216
rect 26608 19780 26660 19786
rect 26608 19722 26660 19728
rect 26620 19446 26648 19722
rect 26608 19440 26660 19446
rect 26608 19382 26660 19388
rect 26896 19310 26924 21490
rect 27264 20602 27292 22066
rect 27344 21956 27396 21962
rect 27344 21898 27396 21904
rect 27356 21554 27384 21898
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 27160 20596 27212 20602
rect 27160 20538 27212 20544
rect 27252 20596 27304 20602
rect 27252 20538 27304 20544
rect 27172 19514 27200 20538
rect 27540 20466 27568 24074
rect 27724 23798 27752 24126
rect 27908 24052 27936 24278
rect 27816 24024 27936 24052
rect 28356 24064 28408 24070
rect 27712 23792 27764 23798
rect 27712 23734 27764 23740
rect 27620 23180 27672 23186
rect 27620 23122 27672 23128
rect 27632 22710 27660 23122
rect 27816 23050 27844 24024
rect 28356 24006 28408 24012
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27804 23044 27856 23050
rect 27804 22986 27856 22992
rect 28368 22982 28396 24006
rect 28356 22976 28408 22982
rect 28356 22918 28408 22924
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 28460 22794 28488 25026
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28552 23118 28580 23666
rect 28644 23254 28672 26200
rect 29184 25832 29236 25838
rect 29184 25774 29236 25780
rect 28724 25152 28776 25158
rect 28724 25094 28776 25100
rect 28736 23254 28764 25094
rect 29000 25016 29052 25022
rect 29000 24958 29052 24964
rect 29012 24206 29040 24958
rect 29092 24404 29144 24410
rect 29092 24346 29144 24352
rect 29000 24200 29052 24206
rect 29000 24142 29052 24148
rect 28816 23520 28868 23526
rect 28816 23462 28868 23468
rect 28828 23322 28856 23462
rect 29104 23322 29132 24346
rect 28816 23316 28868 23322
rect 28816 23258 28868 23264
rect 29092 23316 29144 23322
rect 29092 23258 29144 23264
rect 28632 23248 28684 23254
rect 28632 23190 28684 23196
rect 28724 23248 28776 23254
rect 28724 23190 28776 23196
rect 28540 23112 28592 23118
rect 28592 23072 28672 23100
rect 28540 23054 28592 23060
rect 28368 22766 28488 22794
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 27804 22228 27856 22234
rect 27804 22170 27856 22176
rect 27620 21412 27672 21418
rect 27620 21354 27672 21360
rect 27632 21010 27660 21354
rect 27816 21146 27844 22170
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 28368 21672 28396 22766
rect 28644 22710 28672 23072
rect 28828 22778 28856 23258
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 28816 22772 28868 22778
rect 28816 22714 28868 22720
rect 28632 22704 28684 22710
rect 28632 22646 28684 22652
rect 28816 22432 28868 22438
rect 28814 22400 28816 22409
rect 28868 22400 28870 22409
rect 28814 22335 28870 22344
rect 28920 22234 28948 23054
rect 29000 22432 29052 22438
rect 29000 22374 29052 22380
rect 28448 22228 28500 22234
rect 28448 22170 28500 22176
rect 28908 22228 28960 22234
rect 28908 22170 28960 22176
rect 28276 21644 28396 21672
rect 27896 21548 27948 21554
rect 27896 21490 27948 21496
rect 27908 21146 27936 21490
rect 27712 21140 27764 21146
rect 27712 21082 27764 21088
rect 27804 21140 27856 21146
rect 27804 21082 27856 21088
rect 27896 21140 27948 21146
rect 27896 21082 27948 21088
rect 27620 21004 27672 21010
rect 27620 20946 27672 20952
rect 27528 20460 27580 20466
rect 27528 20402 27580 20408
rect 27540 19938 27568 20402
rect 27632 20330 27660 20946
rect 27620 20324 27672 20330
rect 27620 20266 27672 20272
rect 27724 20262 27752 21082
rect 28276 21078 28304 21644
rect 28460 21486 28488 22170
rect 28538 21992 28594 22001
rect 28538 21927 28594 21936
rect 28448 21480 28500 21486
rect 28368 21440 28448 21468
rect 28264 21072 28316 21078
rect 28264 21014 28316 21020
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 28368 20398 28396 21440
rect 28448 21422 28500 21428
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28356 20392 28408 20398
rect 28356 20334 28408 20340
rect 27896 20324 27948 20330
rect 27896 20266 27948 20272
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27540 19910 27660 19938
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27160 19508 27212 19514
rect 27160 19450 27212 19456
rect 27264 19446 27292 19790
rect 26976 19440 27028 19446
rect 26976 19382 27028 19388
rect 27252 19440 27304 19446
rect 27252 19382 27304 19388
rect 26884 19304 26936 19310
rect 26884 19246 26936 19252
rect 26608 19168 26660 19174
rect 26608 19110 26660 19116
rect 26514 18864 26570 18873
rect 26514 18799 26570 18808
rect 26528 16697 26556 18799
rect 26620 17814 26648 19110
rect 26792 18896 26844 18902
rect 26792 18838 26844 18844
rect 26804 18154 26832 18838
rect 26988 18698 27016 19382
rect 27434 19272 27490 19281
rect 27434 19207 27436 19216
rect 27488 19207 27490 19216
rect 27436 19178 27488 19184
rect 27632 19174 27660 19910
rect 27908 19718 27936 20266
rect 27988 19984 28040 19990
rect 27988 19926 28040 19932
rect 28000 19854 28028 19926
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 27896 19712 27948 19718
rect 27896 19654 27948 19660
rect 28356 19712 28408 19718
rect 28356 19654 28408 19660
rect 28460 19666 28488 20878
rect 28552 19854 28580 21927
rect 28632 21888 28684 21894
rect 28632 21830 28684 21836
rect 28644 20913 28672 21830
rect 29012 21622 29040 22374
rect 29196 22094 29224 25774
rect 29288 24274 29316 26200
rect 29552 24744 29604 24750
rect 29552 24686 29604 24692
rect 29276 24268 29328 24274
rect 29276 24210 29328 24216
rect 29564 23866 29592 24686
rect 30012 24676 30064 24682
rect 30012 24618 30064 24624
rect 30024 24274 30052 24618
rect 30012 24268 30064 24274
rect 30012 24210 30064 24216
rect 29552 23860 29604 23866
rect 29552 23802 29604 23808
rect 29564 23730 29592 23802
rect 30116 23798 30144 26302
rect 30562 26200 30618 27000
rect 31206 26200 31262 27000
rect 31850 26200 31906 27000
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26330 33838 27000
rect 33782 26302 34100 26330
rect 33782 26200 33838 26302
rect 30288 25220 30340 25226
rect 30288 25162 30340 25168
rect 30196 24200 30248 24206
rect 30196 24142 30248 24148
rect 30104 23792 30156 23798
rect 30104 23734 30156 23740
rect 29552 23724 29604 23730
rect 29552 23666 29604 23672
rect 29734 23488 29790 23497
rect 29734 23423 29790 23432
rect 29748 23254 29776 23423
rect 29736 23248 29788 23254
rect 29736 23190 29788 23196
rect 29828 22976 29880 22982
rect 29828 22918 29880 22924
rect 29840 22098 29868 22918
rect 29104 22066 29224 22094
rect 29828 22092 29880 22098
rect 30116 22094 30144 23734
rect 30208 23361 30236 24142
rect 30300 23730 30328 25162
rect 30472 24812 30524 24818
rect 30472 24754 30524 24760
rect 30380 24336 30432 24342
rect 30380 24278 30432 24284
rect 30392 24070 30420 24278
rect 30380 24064 30432 24070
rect 30380 24006 30432 24012
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 30194 23352 30250 23361
rect 30194 23287 30250 23296
rect 30484 23202 30512 24754
rect 30576 24206 30604 26200
rect 30564 24200 30616 24206
rect 30564 24142 30616 24148
rect 30562 23896 30618 23905
rect 30562 23831 30618 23840
rect 30576 23662 30604 23831
rect 30944 23684 31156 23712
rect 30564 23656 30616 23662
rect 30944 23610 30972 23684
rect 30564 23598 30616 23604
rect 30852 23594 30972 23610
rect 30840 23588 30972 23594
rect 30892 23582 30972 23588
rect 31024 23588 31076 23594
rect 30840 23530 30892 23536
rect 31024 23530 31076 23536
rect 30484 23174 30604 23202
rect 30286 23080 30342 23089
rect 30286 23015 30288 23024
rect 30340 23015 30342 23024
rect 30288 22986 30340 22992
rect 30576 22778 30604 23174
rect 30840 22976 30892 22982
rect 30840 22918 30892 22924
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 30852 22574 30880 22918
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30840 22568 30892 22574
rect 30840 22510 30892 22516
rect 28724 21616 28776 21622
rect 28724 21558 28776 21564
rect 29000 21616 29052 21622
rect 29000 21558 29052 21564
rect 28736 21486 28764 21558
rect 28724 21480 28776 21486
rect 28724 21422 28776 21428
rect 28816 21480 28868 21486
rect 28868 21428 28948 21434
rect 28816 21422 28948 21428
rect 28736 21321 28764 21422
rect 28828 21406 28948 21422
rect 28722 21312 28778 21321
rect 28722 21247 28778 21256
rect 28920 21146 28948 21406
rect 28908 21140 28960 21146
rect 28908 21082 28960 21088
rect 28630 20904 28686 20913
rect 28630 20839 28686 20848
rect 28632 20256 28684 20262
rect 28632 20198 28684 20204
rect 28540 19848 28592 19854
rect 28540 19790 28592 19796
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 27804 19304 27856 19310
rect 27804 19246 27856 19252
rect 27620 19168 27672 19174
rect 27620 19110 27672 19116
rect 27252 18964 27304 18970
rect 27252 18906 27304 18912
rect 26976 18692 27028 18698
rect 26976 18634 27028 18640
rect 26988 18426 27016 18634
rect 27264 18465 27292 18906
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 27250 18456 27306 18465
rect 26976 18420 27028 18426
rect 27250 18391 27306 18400
rect 26976 18362 27028 18368
rect 26792 18148 26844 18154
rect 26792 18090 26844 18096
rect 26608 17808 26660 17814
rect 26608 17750 26660 17756
rect 26988 17610 27016 18362
rect 27068 18216 27120 18222
rect 27068 18158 27120 18164
rect 26976 17604 27028 17610
rect 26976 17546 27028 17552
rect 26988 17270 27016 17546
rect 26976 17264 27028 17270
rect 26976 17206 27028 17212
rect 26514 16688 26570 16697
rect 26514 16623 26570 16632
rect 26988 16250 27016 17206
rect 27080 16658 27108 18158
rect 27344 18080 27396 18086
rect 27344 18022 27396 18028
rect 27356 17610 27384 18022
rect 27344 17604 27396 17610
rect 27344 17546 27396 17552
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27160 16992 27212 16998
rect 27160 16934 27212 16940
rect 27172 16658 27200 16934
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 26976 16244 27028 16250
rect 26976 16186 27028 16192
rect 26988 16130 27016 16186
rect 26988 16102 27108 16130
rect 26884 15360 26936 15366
rect 26884 15302 26936 15308
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26620 14482 26648 14758
rect 26896 14550 26924 15302
rect 27080 15162 27108 16102
rect 27172 16046 27200 16594
rect 27632 16590 27660 17070
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27160 16040 27212 16046
rect 27160 15982 27212 15988
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 26884 14544 26936 14550
rect 26884 14486 26936 14492
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 27528 13252 27580 13258
rect 27528 13194 27580 13200
rect 27540 11218 27568 13194
rect 27528 11212 27580 11218
rect 27632 11200 27660 16186
rect 27724 11665 27752 18702
rect 27816 18290 27844 19246
rect 28368 19174 28396 19654
rect 28460 19638 28580 19666
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 27804 18284 27856 18290
rect 27804 18226 27856 18232
rect 27816 17746 27844 18226
rect 27804 17740 27856 17746
rect 27804 17682 27856 17688
rect 27816 17202 27844 17682
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 28368 17218 28396 19110
rect 28448 17808 28500 17814
rect 28448 17750 28500 17756
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 28276 17190 28396 17218
rect 28276 16454 28304 17190
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 28368 16250 28396 16526
rect 28460 16522 28488 17750
rect 28552 16561 28580 19638
rect 28644 19446 28672 20198
rect 28724 19916 28776 19922
rect 28724 19858 28776 19864
rect 28632 19440 28684 19446
rect 28632 19382 28684 19388
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 28644 18358 28672 19110
rect 28632 18352 28684 18358
rect 28632 18294 28684 18300
rect 28736 16658 28764 19858
rect 28724 16652 28776 16658
rect 28724 16594 28776 16600
rect 28538 16552 28594 16561
rect 28448 16516 28500 16522
rect 28538 16487 28594 16496
rect 28448 16458 28500 16464
rect 28540 16448 28592 16454
rect 28540 16390 28592 16396
rect 28356 16244 28408 16250
rect 28356 16186 28408 16192
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27710 11656 27766 11665
rect 27710 11591 27766 11600
rect 27632 11172 27752 11200
rect 27528 11154 27580 11160
rect 27620 11076 27672 11082
rect 27620 11018 27672 11024
rect 27632 7546 27660 11018
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27724 7426 27752 11172
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 28448 9580 28500 9586
rect 28448 9522 28500 9528
rect 28460 9382 28488 9522
rect 28448 9376 28500 9382
rect 28448 9318 28500 9324
rect 28460 9178 28488 9318
rect 28448 9172 28500 9178
rect 28448 9114 28500 9120
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27632 7398 27752 7426
rect 27160 5636 27212 5642
rect 27160 5578 27212 5584
rect 27172 5370 27200 5578
rect 27632 5574 27660 7398
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27620 5568 27672 5574
rect 27620 5510 27672 5516
rect 27160 5364 27212 5370
rect 27160 5306 27212 5312
rect 25964 4548 26016 4554
rect 25964 4490 26016 4496
rect 26424 4548 26476 4554
rect 26424 4490 26476 4496
rect 27528 4548 27580 4554
rect 27528 4490 27580 4496
rect 27540 3602 27568 4490
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 27632 3534 27660 5510
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 28552 5302 28580 16390
rect 28920 5778 28948 21082
rect 29104 21010 29132 22066
rect 29828 22034 29880 22040
rect 30024 22066 30144 22094
rect 30748 22094 30800 22098
rect 30852 22094 30880 22510
rect 30944 22409 30972 22578
rect 30930 22400 30986 22409
rect 30930 22335 30986 22344
rect 30930 22264 30986 22273
rect 30930 22199 30986 22208
rect 30748 22092 30880 22094
rect 29276 21956 29328 21962
rect 29276 21898 29328 21904
rect 29092 21004 29144 21010
rect 29092 20946 29144 20952
rect 29288 20942 29316 21898
rect 29840 21729 29868 22034
rect 29826 21720 29882 21729
rect 29826 21655 29882 21664
rect 29840 21554 29868 21655
rect 29828 21548 29880 21554
rect 29828 21490 29880 21496
rect 29276 20936 29328 20942
rect 29276 20878 29328 20884
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 29564 20602 29592 20878
rect 29552 20596 29604 20602
rect 29552 20538 29604 20544
rect 29092 17672 29144 17678
rect 29092 17614 29144 17620
rect 29104 17338 29132 17614
rect 29092 17332 29144 17338
rect 29092 17274 29144 17280
rect 29564 16017 29592 20538
rect 29736 20460 29788 20466
rect 29840 20448 29868 21490
rect 30024 21146 30052 22066
rect 30800 22066 30880 22092
rect 30748 22034 30800 22040
rect 30748 21956 30800 21962
rect 30748 21898 30800 21904
rect 30104 21888 30156 21894
rect 30104 21830 30156 21836
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 30116 21350 30144 21830
rect 30104 21344 30156 21350
rect 30104 21286 30156 21292
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 30012 21140 30064 21146
rect 30012 21082 30064 21088
rect 30104 21140 30156 21146
rect 30104 21082 30156 21088
rect 30116 20505 30144 21082
rect 29788 20420 29868 20448
rect 30102 20496 30158 20505
rect 30102 20431 30158 20440
rect 29736 20402 29788 20408
rect 29644 19984 29696 19990
rect 29748 19972 29776 20402
rect 30208 20398 30236 21286
rect 30484 21010 30512 21830
rect 30656 21344 30708 21350
rect 30656 21286 30708 21292
rect 30472 21004 30524 21010
rect 30472 20946 30524 20952
rect 30196 20392 30248 20398
rect 30196 20334 30248 20340
rect 30288 20392 30340 20398
rect 30288 20334 30340 20340
rect 30196 20256 30248 20262
rect 30196 20198 30248 20204
rect 29696 19944 29776 19972
rect 29644 19926 29696 19932
rect 29656 19378 29684 19926
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 29656 18358 29684 19314
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29736 18624 29788 18630
rect 29736 18566 29788 18572
rect 29644 18352 29696 18358
rect 29644 18294 29696 18300
rect 29656 17746 29684 18294
rect 29644 17740 29696 17746
rect 29644 17682 29696 17688
rect 29656 17610 29684 17682
rect 29644 17604 29696 17610
rect 29644 17546 29696 17552
rect 29656 17338 29684 17546
rect 29644 17332 29696 17338
rect 29644 17274 29696 17280
rect 29550 16008 29606 16017
rect 29550 15943 29606 15952
rect 29748 15638 29776 18566
rect 29840 18086 29868 18702
rect 29828 18080 29880 18086
rect 29828 18022 29880 18028
rect 29736 15632 29788 15638
rect 29736 15574 29788 15580
rect 29932 15473 29960 19790
rect 30208 18834 30236 20198
rect 30300 19174 30328 20334
rect 30484 19718 30512 20946
rect 30668 20806 30696 21286
rect 30656 20800 30708 20806
rect 30656 20742 30708 20748
rect 30472 19712 30524 19718
rect 30472 19654 30524 19660
rect 30654 19408 30710 19417
rect 30654 19343 30656 19352
rect 30708 19343 30710 19352
rect 30656 19314 30708 19320
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 30656 18692 30708 18698
rect 30656 18634 30708 18640
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 30116 18426 30144 18566
rect 30668 18426 30696 18634
rect 30104 18420 30156 18426
rect 30104 18362 30156 18368
rect 30656 18420 30708 18426
rect 30656 18362 30708 18368
rect 30656 18284 30708 18290
rect 30656 18226 30708 18232
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 30392 18034 30420 18090
rect 30300 18006 30420 18034
rect 30300 17746 30328 18006
rect 30668 17921 30696 18226
rect 30654 17912 30710 17921
rect 30654 17847 30710 17856
rect 30288 17740 30340 17746
rect 30288 17682 30340 17688
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30208 17338 30236 17478
rect 30196 17332 30248 17338
rect 30196 17274 30248 17280
rect 30208 17066 30236 17274
rect 30300 17134 30328 17682
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30196 17060 30248 17066
rect 30196 17002 30248 17008
rect 30208 16794 30236 17002
rect 30196 16788 30248 16794
rect 30196 16730 30248 16736
rect 29918 15464 29974 15473
rect 29918 15399 29974 15408
rect 30760 13433 30788 21898
rect 30944 20602 30972 22199
rect 30932 20596 30984 20602
rect 30932 20538 30984 20544
rect 30840 20052 30892 20058
rect 30840 19994 30892 20000
rect 30852 19786 30880 19994
rect 30840 19780 30892 19786
rect 30840 19722 30892 19728
rect 30840 19304 30892 19310
rect 30840 19246 30892 19252
rect 30852 18834 30880 19246
rect 30840 18828 30892 18834
rect 30840 18770 30892 18776
rect 31036 18290 31064 23530
rect 31128 22273 31156 23684
rect 31220 22574 31248 26200
rect 31298 24712 31354 24721
rect 31298 24647 31354 24656
rect 31312 23526 31340 24647
rect 31864 24206 31892 26200
rect 32220 25356 32272 25362
rect 32220 25298 32272 25304
rect 31576 24200 31628 24206
rect 31576 24142 31628 24148
rect 31852 24200 31904 24206
rect 31852 24142 31904 24148
rect 31392 23724 31444 23730
rect 31392 23666 31444 23672
rect 31404 23526 31432 23666
rect 31300 23520 31352 23526
rect 31300 23462 31352 23468
rect 31392 23520 31444 23526
rect 31392 23462 31444 23468
rect 31298 23352 31354 23361
rect 31298 23287 31300 23296
rect 31352 23287 31354 23296
rect 31300 23258 31352 23264
rect 31404 23186 31432 23462
rect 31392 23180 31444 23186
rect 31392 23122 31444 23128
rect 31484 23112 31536 23118
rect 31484 23054 31536 23060
rect 31300 22636 31352 22642
rect 31300 22578 31352 22584
rect 31208 22568 31260 22574
rect 31208 22510 31260 22516
rect 31312 22409 31340 22578
rect 31298 22400 31354 22409
rect 31298 22335 31354 22344
rect 31114 22264 31170 22273
rect 31114 22199 31170 22208
rect 31114 21448 31170 21457
rect 31114 21383 31170 21392
rect 31128 20942 31156 21383
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 31208 20800 31260 20806
rect 31208 20742 31260 20748
rect 31220 18329 31248 20742
rect 31206 18320 31262 18329
rect 31024 18284 31076 18290
rect 31206 18255 31262 18264
rect 31024 18226 31076 18232
rect 31312 17678 31340 22335
rect 31496 21729 31524 23054
rect 31482 21720 31538 21729
rect 31482 21655 31538 21664
rect 31496 21554 31524 21655
rect 31484 21548 31536 21554
rect 31484 21490 31536 21496
rect 31392 21412 31444 21418
rect 31392 21354 31444 21360
rect 31404 21146 31432 21354
rect 31392 21140 31444 21146
rect 31392 21082 31444 21088
rect 31496 20398 31524 21490
rect 31588 21486 31616 24142
rect 31852 24064 31904 24070
rect 31852 24006 31904 24012
rect 31668 23656 31720 23662
rect 31668 23598 31720 23604
rect 31680 23497 31708 23598
rect 31666 23488 31722 23497
rect 31666 23423 31722 23432
rect 31680 22234 31708 23423
rect 31864 23118 31892 24006
rect 32036 23724 32088 23730
rect 32036 23666 32088 23672
rect 31944 23180 31996 23186
rect 31944 23122 31996 23128
rect 31852 23112 31904 23118
rect 31852 23054 31904 23060
rect 31852 22976 31904 22982
rect 31772 22936 31852 22964
rect 31668 22228 31720 22234
rect 31668 22170 31720 22176
rect 31668 21888 31720 21894
rect 31668 21830 31720 21836
rect 31576 21480 31628 21486
rect 31576 21422 31628 21428
rect 31680 21010 31708 21830
rect 31772 21350 31800 22936
rect 31852 22918 31904 22924
rect 31956 22506 31984 23122
rect 31944 22500 31996 22506
rect 31944 22442 31996 22448
rect 31852 22160 31904 22166
rect 31852 22102 31904 22108
rect 31760 21344 31812 21350
rect 31760 21286 31812 21292
rect 31864 21049 31892 22102
rect 31850 21040 31906 21049
rect 31668 21004 31720 21010
rect 31850 20975 31906 20984
rect 31668 20946 31720 20952
rect 31852 20868 31904 20874
rect 31852 20810 31904 20816
rect 31484 20392 31536 20398
rect 31484 20334 31536 20340
rect 31864 19961 31892 20810
rect 31944 20800 31996 20806
rect 31944 20742 31996 20748
rect 31850 19952 31906 19961
rect 31850 19887 31906 19896
rect 30840 17672 30892 17678
rect 30840 17614 30892 17620
rect 31300 17672 31352 17678
rect 31956 17649 31984 20742
rect 32048 19446 32076 23666
rect 32232 23662 32260 25298
rect 32508 24682 32536 26200
rect 32864 25424 32916 25430
rect 32864 25366 32916 25372
rect 32588 25288 32640 25294
rect 32588 25230 32640 25236
rect 32496 24676 32548 24682
rect 32496 24618 32548 24624
rect 32312 24064 32364 24070
rect 32312 24006 32364 24012
rect 32324 23905 32352 24006
rect 32310 23896 32366 23905
rect 32310 23831 32366 23840
rect 32220 23656 32272 23662
rect 32220 23598 32272 23604
rect 32220 23520 32272 23526
rect 32220 23462 32272 23468
rect 32496 23520 32548 23526
rect 32496 23462 32548 23468
rect 32232 22710 32260 23462
rect 32404 23044 32456 23050
rect 32404 22986 32456 22992
rect 32220 22704 32272 22710
rect 32220 22646 32272 22652
rect 32312 22636 32364 22642
rect 32312 22578 32364 22584
rect 32324 21894 32352 22578
rect 32416 22166 32444 22986
rect 32508 22930 32536 23462
rect 32600 23254 32628 25230
rect 32680 24200 32732 24206
rect 32680 24142 32732 24148
rect 32588 23248 32640 23254
rect 32588 23190 32640 23196
rect 32508 22902 32628 22930
rect 32494 22536 32550 22545
rect 32494 22471 32550 22480
rect 32508 22438 32536 22471
rect 32496 22432 32548 22438
rect 32496 22374 32548 22380
rect 32404 22160 32456 22166
rect 32404 22102 32456 22108
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 32312 21888 32364 21894
rect 32312 21830 32364 21836
rect 32220 21548 32272 21554
rect 32220 21490 32272 21496
rect 32232 19825 32260 21490
rect 32218 19816 32274 19825
rect 32218 19751 32274 19760
rect 32036 19440 32088 19446
rect 32036 19382 32088 19388
rect 31300 17614 31352 17620
rect 31942 17640 31998 17649
rect 30852 17338 30880 17614
rect 30932 17604 30984 17610
rect 31942 17575 31998 17584
rect 30932 17546 30984 17552
rect 30944 17338 30972 17546
rect 30840 17332 30892 17338
rect 30840 17274 30892 17280
rect 30932 17332 30984 17338
rect 30932 17274 30984 17280
rect 30852 16658 30880 17274
rect 30944 17066 30972 17274
rect 31760 17196 31812 17202
rect 31760 17138 31812 17144
rect 30932 17060 30984 17066
rect 30932 17002 30984 17008
rect 30840 16652 30892 16658
rect 30840 16594 30892 16600
rect 30746 13424 30802 13433
rect 30746 13359 30802 13368
rect 31772 11354 31800 17138
rect 32324 12434 32352 21830
rect 32416 21418 32444 21966
rect 32404 21412 32456 21418
rect 32404 21354 32456 21360
rect 32496 21344 32548 21350
rect 32496 21286 32548 21292
rect 32508 13530 32536 21286
rect 32600 21146 32628 22902
rect 32692 22094 32720 24142
rect 32876 23798 32904 25366
rect 33152 24698 33180 26200
rect 33692 25764 33744 25770
rect 33692 25706 33744 25712
rect 33600 25560 33652 25566
rect 33600 25502 33652 25508
rect 33508 24880 33560 24886
rect 33508 24822 33560 24828
rect 33152 24670 33364 24698
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 33336 24206 33364 24670
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 32864 23792 32916 23798
rect 32864 23734 32916 23740
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 33048 23316 33100 23322
rect 33048 23258 33100 23264
rect 32956 22976 33008 22982
rect 32956 22918 33008 22924
rect 32968 22778 32996 22918
rect 33060 22778 33088 23258
rect 33336 23202 33364 24142
rect 33416 24064 33468 24070
rect 33416 24006 33468 24012
rect 33428 23769 33456 24006
rect 33414 23760 33470 23769
rect 33414 23695 33470 23704
rect 33520 23254 33548 24822
rect 33612 23866 33640 25502
rect 33600 23860 33652 23866
rect 33600 23802 33652 23808
rect 33704 23254 33732 25706
rect 34072 24206 34100 26302
rect 34426 26200 34482 27000
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26200 36414 27000
rect 37002 26330 37058 27000
rect 37002 26302 37228 26330
rect 37002 26200 37058 26302
rect 34152 24608 34204 24614
rect 34152 24550 34204 24556
rect 34164 24410 34192 24550
rect 34152 24404 34204 24410
rect 34440 24392 34468 26200
rect 34796 25628 34848 25634
rect 34796 25570 34848 25576
rect 34440 24364 34560 24392
rect 34152 24346 34204 24352
rect 34060 24200 34112 24206
rect 34060 24142 34112 24148
rect 34532 24138 34560 24364
rect 34520 24132 34572 24138
rect 34520 24074 34572 24080
rect 34808 23866 34836 25570
rect 35084 24290 35112 26200
rect 35624 25492 35676 25498
rect 35624 25434 35676 25440
rect 35084 24262 35204 24290
rect 35070 24168 35126 24177
rect 34980 24132 35032 24138
rect 35176 24138 35204 24262
rect 35070 24103 35126 24112
rect 35164 24132 35216 24138
rect 34980 24074 35032 24080
rect 34796 23860 34848 23866
rect 34796 23802 34848 23808
rect 34704 23724 34756 23730
rect 34704 23666 34756 23672
rect 34520 23656 34572 23662
rect 34520 23598 34572 23604
rect 33508 23248 33560 23254
rect 33336 23174 33456 23202
rect 33508 23190 33560 23196
rect 33692 23248 33744 23254
rect 33692 23190 33744 23196
rect 33324 23044 33376 23050
rect 33324 22986 33376 22992
rect 32956 22772 33008 22778
rect 32956 22714 33008 22720
rect 33048 22772 33100 22778
rect 33048 22714 33100 22720
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 33232 22228 33284 22234
rect 33232 22170 33284 22176
rect 32772 22094 32824 22098
rect 32692 22092 32824 22094
rect 32692 22066 32772 22092
rect 32772 22034 32824 22040
rect 32864 22024 32916 22030
rect 32864 21966 32916 21972
rect 32588 21140 32640 21146
rect 32588 21082 32640 21088
rect 32680 20936 32732 20942
rect 32680 20878 32732 20884
rect 32692 18193 32720 20878
rect 32678 18184 32734 18193
rect 32678 18119 32734 18128
rect 32496 13524 32548 13530
rect 32496 13466 32548 13472
rect 32324 12406 32444 12434
rect 31760 11348 31812 11354
rect 31760 11290 31812 11296
rect 31300 11076 31352 11082
rect 31300 11018 31352 11024
rect 31312 9654 31340 11018
rect 31300 9648 31352 9654
rect 31300 9590 31352 9596
rect 32416 8634 32444 12406
rect 32404 8628 32456 8634
rect 32404 8570 32456 8576
rect 32876 8362 32904 21966
rect 33244 21690 33272 22170
rect 33336 22030 33364 22986
rect 33428 22506 33456 23174
rect 33508 23044 33560 23050
rect 33508 22986 33560 22992
rect 33416 22500 33468 22506
rect 33416 22442 33468 22448
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 33232 21684 33284 21690
rect 33232 21626 33284 21632
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 33336 15065 33364 21966
rect 33416 21344 33468 21350
rect 33416 21286 33468 21292
rect 33428 21078 33456 21286
rect 33416 21072 33468 21078
rect 33416 21014 33468 21020
rect 33520 19990 33548 22986
rect 33874 22672 33930 22681
rect 33874 22607 33876 22616
rect 33928 22607 33930 22616
rect 33876 22578 33928 22584
rect 33600 22568 33652 22574
rect 33600 22510 33652 22516
rect 33612 22137 33640 22510
rect 33598 22128 33654 22137
rect 33598 22063 33654 22072
rect 34532 21622 34560 23598
rect 34716 22778 34744 23666
rect 34992 23254 35020 24074
rect 35084 24070 35112 24103
rect 35164 24074 35216 24080
rect 35072 24064 35124 24070
rect 35072 24006 35124 24012
rect 35636 23798 35664 25434
rect 35728 24426 35756 26200
rect 35990 24848 36046 24857
rect 35990 24783 36046 24792
rect 35728 24398 35940 24426
rect 35808 24336 35860 24342
rect 35808 24278 35860 24284
rect 35716 24132 35768 24138
rect 35716 24074 35768 24080
rect 35728 23798 35756 24074
rect 35624 23792 35676 23798
rect 35624 23734 35676 23740
rect 35716 23792 35768 23798
rect 35716 23734 35768 23740
rect 34888 23248 34940 23254
rect 34886 23216 34888 23225
rect 34980 23248 35032 23254
rect 34940 23216 34942 23225
rect 34980 23190 35032 23196
rect 34886 23151 34942 23160
rect 35072 23112 35124 23118
rect 35070 23080 35072 23089
rect 35716 23112 35768 23118
rect 35124 23080 35126 23089
rect 34992 23038 35070 23066
rect 34704 22772 34756 22778
rect 34704 22714 34756 22720
rect 34992 22642 35020 23038
rect 35716 23054 35768 23060
rect 35070 23015 35126 23024
rect 35532 22976 35584 22982
rect 35532 22918 35584 22924
rect 35072 22772 35124 22778
rect 35072 22714 35124 22720
rect 34980 22636 35032 22642
rect 34980 22578 35032 22584
rect 34520 21616 34572 21622
rect 34520 21558 34572 21564
rect 33508 19984 33560 19990
rect 33508 19926 33560 19932
rect 33322 15056 33378 15065
rect 33322 14991 33378 15000
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 35084 14618 35112 22714
rect 35544 21554 35572 22918
rect 35728 22438 35756 23054
rect 35716 22432 35768 22438
rect 35716 22374 35768 22380
rect 35820 21962 35848 24278
rect 35912 24206 35940 24398
rect 35900 24200 35952 24206
rect 35900 24142 35952 24148
rect 36004 24070 36032 24783
rect 36268 24676 36320 24682
rect 36268 24618 36320 24624
rect 35992 24064 36044 24070
rect 35992 24006 36044 24012
rect 36280 23730 36308 24618
rect 36372 23730 36400 26200
rect 36912 24336 36964 24342
rect 36912 24278 36964 24284
rect 36820 24200 36872 24206
rect 36820 24142 36872 24148
rect 36452 24064 36504 24070
rect 36452 24006 36504 24012
rect 36268 23724 36320 23730
rect 36268 23666 36320 23672
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 36084 23520 36136 23526
rect 36084 23462 36136 23468
rect 36096 23186 36124 23462
rect 36280 23322 36308 23666
rect 36268 23316 36320 23322
rect 36268 23258 36320 23264
rect 36084 23180 36136 23186
rect 36084 23122 36136 23128
rect 36176 22976 36228 22982
rect 36176 22918 36228 22924
rect 35808 21956 35860 21962
rect 35808 21898 35860 21904
rect 36188 21593 36216 22918
rect 36174 21584 36230 21593
rect 35532 21548 35584 21554
rect 36174 21519 36230 21528
rect 35532 21490 35584 21496
rect 36464 21010 36492 24006
rect 36832 23322 36860 24142
rect 36820 23316 36872 23322
rect 36820 23258 36872 23264
rect 36452 21004 36504 21010
rect 36452 20946 36504 20952
rect 36924 20466 36952 24278
rect 37200 24188 37228 26302
rect 37646 26200 37702 27000
rect 38290 26330 38346 27000
rect 38934 26330 38990 27000
rect 38290 26302 38516 26330
rect 38290 26200 38346 26302
rect 37280 24200 37332 24206
rect 37200 24160 37280 24188
rect 37280 24142 37332 24148
rect 37188 23588 37240 23594
rect 37188 23530 37240 23536
rect 36912 20460 36964 20466
rect 36912 20402 36964 20408
rect 37200 19854 37228 23530
rect 37292 23322 37320 24142
rect 37660 23730 37688 26200
rect 38488 24206 38516 26302
rect 38934 26302 39252 26330
rect 38934 26200 38990 26302
rect 38658 24984 38714 24993
rect 38658 24919 38714 24928
rect 38672 24342 38700 24919
rect 38660 24336 38712 24342
rect 38660 24278 38712 24284
rect 39224 24206 39252 26302
rect 39578 26200 39634 27000
rect 40222 26330 40278 27000
rect 40222 26302 40356 26330
rect 40222 26200 40278 26302
rect 39304 24948 39356 24954
rect 39304 24890 39356 24896
rect 39316 24410 39344 24890
rect 39304 24404 39356 24410
rect 39304 24346 39356 24352
rect 39592 24274 39620 26200
rect 40130 24304 40186 24313
rect 39580 24268 39632 24274
rect 40130 24239 40132 24248
rect 39580 24210 39632 24216
rect 40184 24239 40186 24248
rect 40132 24210 40184 24216
rect 38476 24200 38528 24206
rect 38476 24142 38528 24148
rect 39212 24200 39264 24206
rect 39212 24142 39264 24148
rect 38292 24132 38344 24138
rect 38292 24074 38344 24080
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 38304 23866 38332 24074
rect 38488 23866 38516 24142
rect 39224 23866 39252 24142
rect 39592 23866 39620 24210
rect 40328 23866 40356 26302
rect 40866 26200 40922 27000
rect 41510 26200 41566 27000
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43442 26330 43498 27000
rect 43442 26302 43852 26330
rect 43442 26200 43498 26302
rect 40684 24336 40736 24342
rect 40684 24278 40736 24284
rect 40696 23866 40724 24278
rect 38292 23860 38344 23866
rect 38292 23802 38344 23808
rect 38476 23860 38528 23866
rect 38476 23802 38528 23808
rect 39212 23860 39264 23866
rect 39212 23802 39264 23808
rect 39580 23860 39632 23866
rect 39580 23802 39632 23808
rect 40316 23860 40368 23866
rect 40316 23802 40368 23808
rect 40684 23860 40736 23866
rect 40684 23802 40736 23808
rect 37648 23724 37700 23730
rect 40880 23712 40908 26200
rect 41524 24206 41552 26200
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 41512 24200 41564 24206
rect 41512 24142 41564 24148
rect 42064 24064 42116 24070
rect 42064 24006 42116 24012
rect 43720 24064 43772 24070
rect 43720 24006 43772 24012
rect 42076 23730 42104 24006
rect 43732 23730 43760 24006
rect 43824 23730 43852 26302
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26330 45430 27000
rect 45374 26302 45508 26330
rect 45374 26200 45430 26302
rect 44100 23746 44128 26200
rect 44744 24410 44772 26200
rect 44732 24404 44784 24410
rect 44732 24346 44784 24352
rect 44744 24206 44772 24346
rect 45480 24290 45508 26302
rect 46018 26200 46074 27000
rect 46662 26200 46718 27000
rect 47306 26200 47362 27000
rect 47950 26200 48006 27000
rect 48594 26200 48650 27000
rect 45480 24262 45600 24290
rect 45572 24206 45600 24262
rect 46032 24206 46060 26200
rect 44364 24200 44416 24206
rect 44364 24142 44416 24148
rect 44732 24200 44784 24206
rect 44732 24142 44784 24148
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 45928 24200 45980 24206
rect 45928 24142 45980 24148
rect 46020 24200 46072 24206
rect 46020 24142 46072 24148
rect 44180 23792 44232 23798
rect 44100 23740 44180 23746
rect 44100 23734 44232 23740
rect 40960 23724 41012 23730
rect 40880 23684 40960 23712
rect 37648 23666 37700 23672
rect 40960 23666 41012 23672
rect 42064 23724 42116 23730
rect 42064 23666 42116 23672
rect 43720 23724 43772 23730
rect 43720 23666 43772 23672
rect 43812 23724 43864 23730
rect 44100 23718 44220 23734
rect 43812 23666 43864 23672
rect 38568 23656 38620 23662
rect 38568 23598 38620 23604
rect 37372 23520 37424 23526
rect 37372 23462 37424 23468
rect 37280 23316 37332 23322
rect 37280 23258 37332 23264
rect 37188 19848 37240 19854
rect 37188 19790 37240 19796
rect 37384 17678 37412 23462
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37740 22432 37792 22438
rect 37740 22374 37792 22380
rect 37752 18222 37780 22374
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 38580 18426 38608 23598
rect 41420 23588 41472 23594
rect 41420 23530 41472 23536
rect 41432 23118 41460 23530
rect 43352 23520 43404 23526
rect 43352 23462 43404 23468
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 43364 23118 43392 23462
rect 44376 23322 44404 24142
rect 45376 24064 45428 24070
rect 45376 24006 45428 24012
rect 44640 23724 44692 23730
rect 44640 23666 44692 23672
rect 44652 23322 44680 23666
rect 44364 23316 44416 23322
rect 44364 23258 44416 23264
rect 44640 23316 44692 23322
rect 44640 23258 44692 23264
rect 41420 23112 41472 23118
rect 41420 23054 41472 23060
rect 43352 23112 43404 23118
rect 43352 23054 43404 23060
rect 39948 22976 40000 22982
rect 39948 22918 40000 22924
rect 39960 22778 39988 22918
rect 39948 22772 40000 22778
rect 39948 22714 40000 22720
rect 44732 22636 44784 22642
rect 44732 22578 44784 22584
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 44744 21894 44772 22578
rect 44732 21888 44784 21894
rect 44732 21830 44784 21836
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 44824 21140 44876 21146
rect 44824 21082 44876 21088
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 38568 18420 38620 18426
rect 38568 18362 38620 18368
rect 37740 18216 37792 18222
rect 37740 18158 37792 18164
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 37372 17672 37424 17678
rect 37372 17614 37424 17620
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 37280 17264 37332 17270
rect 37280 17206 37332 17212
rect 37292 15502 37320 17206
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 37280 15496 37332 15502
rect 37280 15438 37332 15444
rect 44836 15366 44864 21082
rect 45388 18737 45416 24006
rect 45940 23866 45968 24142
rect 45928 23860 45980 23866
rect 45928 23802 45980 23808
rect 46676 23730 46704 26200
rect 47320 24206 47348 26200
rect 47308 24200 47360 24206
rect 47308 24142 47360 24148
rect 46848 24064 46900 24070
rect 46848 24006 46900 24012
rect 47124 24064 47176 24070
rect 47124 24006 47176 24012
rect 46664 23724 46716 23730
rect 46664 23666 46716 23672
rect 45744 23520 45796 23526
rect 45744 23462 45796 23468
rect 45756 18873 45784 23462
rect 45742 18864 45798 18873
rect 45742 18799 45798 18808
rect 45374 18728 45430 18737
rect 45374 18663 45430 18672
rect 46860 17241 46888 24006
rect 46940 23520 46992 23526
rect 46940 23462 46992 23468
rect 47032 23520 47084 23526
rect 47032 23462 47084 23468
rect 46952 18834 46980 23462
rect 47044 18970 47072 23462
rect 47032 18964 47084 18970
rect 47032 18906 47084 18912
rect 46940 18828 46992 18834
rect 46940 18770 46992 18776
rect 46846 17232 46902 17241
rect 46846 17167 46902 17176
rect 47136 16998 47164 24006
rect 47320 23866 47348 24142
rect 47964 24052 47992 26200
rect 48318 24848 48374 24857
rect 48318 24783 48374 24792
rect 47872 24024 47992 24052
rect 47308 23860 47360 23866
rect 47308 23802 47360 23808
rect 47768 23724 47820 23730
rect 47768 23666 47820 23672
rect 47492 22976 47544 22982
rect 47492 22918 47544 22924
rect 47400 22500 47452 22506
rect 47400 22442 47452 22448
rect 47412 17066 47440 22442
rect 47504 21146 47532 22918
rect 47780 22778 47808 23666
rect 47872 23118 47900 24024
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 48226 23760 48282 23769
rect 48332 23730 48360 24783
rect 48608 24290 48636 26200
rect 48516 24262 48636 24290
rect 48226 23695 48282 23704
rect 48320 23724 48372 23730
rect 47860 23112 47912 23118
rect 47860 23054 47912 23060
rect 48240 23066 48268 23695
rect 48320 23666 48372 23672
rect 48516 23118 48544 24262
rect 48596 24200 48648 24206
rect 48596 24142 48648 24148
rect 48608 23322 48636 24142
rect 48688 24064 48740 24070
rect 48688 24006 48740 24012
rect 48700 23730 48728 24006
rect 48688 23724 48740 23730
rect 48688 23666 48740 23672
rect 48688 23520 48740 23526
rect 48688 23462 48740 23468
rect 48596 23316 48648 23322
rect 48596 23258 48648 23264
rect 48504 23112 48556 23118
rect 48240 23038 48360 23066
rect 48504 23054 48556 23060
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 47768 22772 47820 22778
rect 47768 22714 47820 22720
rect 48332 22642 48360 23038
rect 48320 22636 48372 22642
rect 48320 22578 48372 22584
rect 48504 22432 48556 22438
rect 48504 22374 48556 22380
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 47860 21548 47912 21554
rect 47860 21490 47912 21496
rect 47872 21350 47900 21490
rect 47860 21344 47912 21350
rect 47860 21286 47912 21292
rect 47492 21140 47544 21146
rect 47492 21082 47544 21088
rect 47400 17060 47452 17066
rect 47400 17002 47452 17008
rect 47124 16992 47176 16998
rect 47124 16934 47176 16940
rect 44824 15360 44876 15366
rect 44824 15302 44876 15308
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 35072 14612 35124 14618
rect 35072 14554 35124 14560
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 47872 11082 47900 21286
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 48516 17270 48544 22374
rect 48700 22030 48728 23462
rect 49054 22944 49110 22953
rect 49054 22879 49110 22888
rect 49068 22642 49096 22879
rect 49056 22636 49108 22642
rect 49056 22578 49108 22584
rect 48688 22024 48740 22030
rect 49056 22024 49108 22030
rect 48688 21966 48740 21972
rect 49054 21992 49056 22001
rect 49108 21992 49110 22001
rect 49054 21927 49110 21936
rect 49068 21146 49096 21927
rect 49240 21888 49292 21894
rect 49240 21830 49292 21836
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 49056 21140 49108 21146
rect 49056 21082 49108 21088
rect 49160 21049 49188 21422
rect 49146 21040 49202 21049
rect 49146 20975 49202 20984
rect 49252 20058 49280 21830
rect 49240 20052 49292 20058
rect 49240 19994 49292 20000
rect 48504 17264 48556 17270
rect 48504 17206 48556 17212
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47860 11076 47912 11082
rect 47860 11018 47912 11024
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 32864 8356 32916 8362
rect 32864 8298 32916 8304
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 28724 5772 28776 5778
rect 28724 5714 28776 5720
rect 28908 5772 28960 5778
rect 28908 5714 28960 5720
rect 28540 5296 28592 5302
rect 28540 5238 28592 5244
rect 27804 4684 27856 4690
rect 27804 4626 27856 4632
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27816 2650 27844 4626
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28736 2650 28764 5714
rect 28816 5160 28868 5166
rect 28816 5102 28868 5108
rect 28828 4826 28856 5102
rect 28816 4820 28868 4826
rect 28816 4762 28868 4768
rect 28920 3670 28948 5714
rect 33508 5092 33560 5098
rect 33508 5034 33560 5040
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 33520 2650 33548 5034
rect 25504 2644 25556 2650
rect 25504 2586 25556 2592
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 28724 2644 28776 2650
rect 28724 2586 28776 2592
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 36372 2514 36400 9114
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 41420 5160 41472 5166
rect 41420 5102 41472 5108
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 38752 3460 38804 3466
rect 38752 3402 38804 3408
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 36360 2508 36412 2514
rect 36360 2450 36412 2456
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 20088 1142 20208 1170
rect 20088 800 20116 1142
rect 22756 800 22784 2450
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 25424 800 25452 2382
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28092 870 28212 898
rect 28092 800 28120 870
rect 1398 0 1454 800
rect 4066 0 4122 800
rect 6734 0 6790 800
rect 9402 0 9458 800
rect 12070 0 12126 800
rect 14738 0 14794 800
rect 17406 0 17462 800
rect 20074 0 20130 800
rect 22742 0 22798 800
rect 25410 0 25466 800
rect 28078 0 28134 800
rect 28184 762 28212 870
rect 28368 762 28396 2382
rect 30760 800 30788 2382
rect 33428 800 33456 2382
rect 36096 800 36124 2382
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38764 800 38792 3402
rect 41432 800 41460 5102
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 44088 3664 44140 3670
rect 44088 3606 44140 3612
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 44100 800 44128 3606
rect 46756 3596 46808 3602
rect 46756 3538 46808 3544
rect 46768 800 46796 3538
rect 49424 3528 49476 3534
rect 49424 3470 49476 3476
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49436 800 49464 3470
rect 28184 734 28396 762
rect 30746 0 30802 800
rect 33414 0 33470 800
rect 36082 0 36138 800
rect 38750 0 38806 800
rect 41418 0 41474 800
rect 44086 0 44142 800
rect 46754 0 46810 800
rect 49422 0 49478 800
<< via2 >>
rect 1306 20712 1362 20768
rect 1214 17040 1270 17096
rect 1306 16632 1362 16688
rect 1306 16224 1362 16280
rect 1306 15816 1362 15872
rect 1306 15408 1362 15464
rect 1306 15000 1362 15056
rect 1306 14592 1362 14648
rect 1306 14184 1362 14240
rect 1214 13368 1270 13424
rect 1306 12144 1362 12200
rect 1398 11736 1454 11792
rect 1674 21800 1730 21856
rect 2134 23432 2190 23488
rect 2134 22344 2190 22400
rect 2778 24384 2834 24440
rect 2042 19896 2098 19952
rect 2226 17720 2282 17776
rect 2042 17448 2098 17504
rect 1766 13932 1822 13968
rect 1766 13912 1768 13932
rect 1768 13912 1820 13932
rect 1820 13912 1822 13932
rect 1766 13268 1768 13288
rect 1768 13268 1820 13288
rect 1820 13268 1822 13288
rect 1766 13232 1822 13268
rect 1674 10920 1730 10976
rect 1582 9696 1638 9752
rect 2042 13776 2098 13832
rect 2042 12552 2098 12608
rect 1766 8880 1822 8936
rect 1306 7656 1362 7712
rect 2226 7792 2282 7848
rect 1306 6432 1362 6488
rect 1306 6024 1362 6080
rect 1306 5652 1308 5672
rect 1308 5652 1360 5672
rect 1360 5652 1362 5672
rect 1306 5616 1362 5652
rect 1306 5228 1362 5264
rect 1306 5208 1308 5228
rect 1308 5208 1360 5228
rect 1360 5208 1362 5228
rect 1306 4800 1362 4856
rect 1306 3168 1362 3224
rect 1306 2760 1362 2816
rect 1214 2352 1270 2408
rect 1306 1944 1362 2000
rect 3054 24792 3110 24848
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 3790 25608 3846 25664
rect 3698 25200 3754 25256
rect 3698 23160 3754 23216
rect 3606 23060 3608 23080
rect 3608 23060 3660 23080
rect 3660 23060 3662 23080
rect 3606 23024 3662 23060
rect 2778 21120 2834 21176
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2962 21528 3018 21584
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2778 19488 2834 19544
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 3606 21392 3662 21448
rect 2962 19216 3018 19272
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 3330 18672 3386 18728
rect 2870 18264 2926 18320
rect 2778 17856 2834 17912
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 4066 23976 4122 24032
rect 3882 23568 3938 23624
rect 4802 24656 4858 24712
rect 4250 24148 4252 24168
rect 4252 24148 4304 24168
rect 4304 24148 4306 24168
rect 4250 24112 4306 24148
rect 4158 22480 4214 22536
rect 3606 19488 3662 19544
rect 3514 16768 3570 16824
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2778 10648 2834 10704
rect 2778 10512 2834 10568
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 3422 12960 3478 13016
rect 2962 12280 3018 12336
rect 3330 12280 3386 12336
rect 3974 21664 4030 21720
rect 4526 22924 4528 22944
rect 4528 22924 4580 22944
rect 4580 22924 4582 22944
rect 4526 22888 4582 22924
rect 4250 21004 4306 21040
rect 4250 20984 4252 21004
rect 4252 20984 4304 21004
rect 4304 20984 4306 21004
rect 3882 20340 3884 20360
rect 3884 20340 3936 20360
rect 3936 20340 3938 20360
rect 3882 20304 3938 20340
rect 3790 17720 3846 17776
rect 4066 20848 4122 20904
rect 4066 19080 4122 19136
rect 3974 17992 4030 18048
rect 4066 17604 4122 17640
rect 4066 17584 4068 17604
rect 4068 17584 4120 17604
rect 4120 17584 4122 17604
rect 4066 17040 4122 17096
rect 3790 15308 3792 15328
rect 3792 15308 3844 15328
rect 3844 15308 3846 15328
rect 3790 15272 3846 15308
rect 4434 18808 4490 18864
rect 4434 17176 4490 17232
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 3606 12144 3662 12200
rect 3514 11192 3570 11248
rect 3698 11192 3754 11248
rect 2870 10104 2926 10160
rect 3422 10104 3478 10160
rect 2778 9288 2834 9344
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2870 8472 2926 8528
rect 2778 8064 2834 8120
rect 3330 8916 3332 8936
rect 3332 8916 3384 8936
rect 3384 8916 3386 8936
rect 3330 8880 3386 8916
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2870 7248 2926 7304
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3698 10376 3754 10432
rect 3698 10104 3754 10160
rect 3606 9444 3662 9480
rect 3606 9424 3608 9444
rect 3608 9424 3660 9444
rect 3660 9424 3662 9444
rect 4618 21936 4674 21992
rect 4986 22752 5042 22808
rect 6550 23468 6552 23488
rect 6552 23468 6604 23488
rect 6604 23468 6606 23488
rect 6550 23432 6606 23468
rect 4802 17856 4858 17912
rect 4894 15680 4950 15736
rect 4802 14048 4858 14104
rect 4250 12280 4306 12336
rect 4158 11328 4214 11384
rect 4434 10648 4490 10704
rect 4250 8492 4306 8528
rect 4250 8472 4252 8492
rect 4252 8472 4304 8492
rect 4304 8472 4306 8492
rect 3606 6840 3662 6896
rect 4710 13132 4712 13152
rect 4712 13132 4764 13152
rect 4764 13132 4766 13152
rect 4710 13096 4766 13132
rect 4618 11056 4674 11112
rect 5262 19372 5318 19408
rect 5262 19352 5264 19372
rect 5264 19352 5316 19372
rect 5316 19352 5318 19372
rect 5630 21256 5686 21312
rect 5722 20712 5778 20768
rect 5630 18284 5686 18320
rect 5630 18264 5632 18284
rect 5632 18264 5684 18284
rect 5684 18264 5686 18284
rect 5630 16632 5686 16688
rect 6182 21528 6238 21584
rect 6090 20304 6146 20360
rect 6090 18400 6146 18456
rect 5906 18164 5908 18184
rect 5908 18164 5960 18184
rect 5960 18164 5962 18184
rect 5906 18128 5962 18164
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 4158 4392 4214 4448
rect 4066 3984 4122 4040
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2870 3576 2926 3632
rect 5722 15000 5778 15056
rect 5354 11464 5410 11520
rect 5446 11056 5502 11112
rect 7102 23568 7158 23624
rect 6642 22072 6698 22128
rect 6458 20304 6514 20360
rect 6458 18128 6514 18184
rect 6182 17448 6238 17504
rect 5538 9560 5594 9616
rect 6458 16496 6514 16552
rect 6734 19896 6790 19952
rect 6734 18284 6790 18320
rect 6734 18264 6736 18284
rect 6736 18264 6788 18284
rect 6788 18264 6790 18284
rect 6458 15408 6514 15464
rect 6918 20712 6974 20768
rect 6458 14476 6514 14512
rect 7194 20712 7250 20768
rect 7378 21256 7434 21312
rect 7286 17856 7342 17912
rect 7194 17604 7250 17640
rect 7194 17584 7196 17604
rect 7196 17584 7248 17604
rect 7248 17584 7250 17604
rect 7470 19352 7526 19408
rect 7378 16088 7434 16144
rect 7378 15272 7434 15328
rect 6458 14456 6460 14476
rect 6460 14456 6512 14476
rect 6512 14456 6514 14476
rect 6458 14320 6514 14376
rect 6550 14068 6606 14104
rect 6550 14048 6552 14068
rect 6552 14048 6604 14068
rect 6604 14048 6606 14068
rect 6182 11872 6238 11928
rect 6366 9560 6422 9616
rect 7286 12688 7342 12744
rect 6734 11600 6790 11656
rect 6918 11464 6974 11520
rect 7194 11076 7250 11112
rect 7194 11056 7196 11076
rect 7196 11056 7248 11076
rect 7248 11056 7250 11076
rect 7010 10648 7066 10704
rect 6918 9968 6974 10024
rect 6642 8628 6698 8664
rect 6642 8608 6644 8628
rect 6644 8608 6696 8628
rect 6696 8608 6698 8628
rect 7378 12280 7434 12336
rect 7562 12416 7618 12472
rect 7378 10376 7434 10432
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7930 23432 7986 23488
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 8022 21564 8024 21584
rect 8024 21564 8076 21584
rect 8076 21564 8078 21584
rect 8022 21528 8078 21564
rect 8206 21528 8262 21584
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 9678 24248 9734 24304
rect 8758 24112 8814 24168
rect 8298 19216 8354 19272
rect 8574 19896 8630 19952
rect 9310 21936 9366 21992
rect 9494 21936 9550 21992
rect 8758 19352 8814 19408
rect 8574 19080 8630 19136
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 8022 17856 8078 17912
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 8114 16768 8170 16824
rect 8206 16516 8262 16552
rect 8206 16496 8208 16516
rect 8208 16496 8260 16516
rect 8260 16496 8262 16516
rect 8390 16632 8446 16688
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7930 16088 7986 16144
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7838 14864 7894 14920
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 8574 17076 8576 17096
rect 8576 17076 8628 17096
rect 8628 17076 8630 17096
rect 8574 17040 8630 17076
rect 8942 17040 8998 17096
rect 8850 16632 8906 16688
rect 8482 15408 8538 15464
rect 8666 15408 8722 15464
rect 8574 15000 8630 15056
rect 8482 14340 8538 14376
rect 8482 14320 8484 14340
rect 8484 14320 8536 14340
rect 8536 14320 8538 14340
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 8850 14864 8906 14920
rect 7746 9016 7802 9072
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 2870 1536 2926 1592
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 8666 9560 8722 9616
rect 11794 23976 11850 24032
rect 12070 23568 12126 23624
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12346 23704 12402 23760
rect 9310 20576 9366 20632
rect 9218 20168 9274 20224
rect 9310 18128 9366 18184
rect 9678 20712 9734 20768
rect 9586 17720 9642 17776
rect 9862 18400 9918 18456
rect 9218 15580 9220 15600
rect 9220 15580 9272 15600
rect 9272 15580 9274 15600
rect 9218 15544 9274 15580
rect 9862 16496 9918 16552
rect 10966 21800 11022 21856
rect 10506 21392 10562 21448
rect 11426 20848 11482 20904
rect 11334 20712 11390 20768
rect 10874 19508 10930 19544
rect 10874 19488 10876 19508
rect 10876 19488 10928 19508
rect 10928 19488 10930 19508
rect 10138 17876 10194 17912
rect 10138 17856 10140 17876
rect 10140 17856 10192 17876
rect 10192 17856 10194 17876
rect 9770 14728 9826 14784
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 9402 13388 9458 13424
rect 9402 13368 9404 13388
rect 9404 13368 9456 13388
rect 9456 13368 9458 13388
rect 9494 11500 9496 11520
rect 9496 11500 9548 11520
rect 9548 11500 9550 11520
rect 9494 11464 9550 11500
rect 10046 11056 10102 11112
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 10598 19216 10654 19272
rect 10506 18536 10562 18592
rect 10414 18400 10470 18456
rect 10598 17856 10654 17912
rect 10598 16244 10654 16280
rect 10598 16224 10600 16244
rect 10600 16224 10652 16244
rect 10652 16224 10654 16244
rect 10690 15816 10746 15872
rect 11058 18808 11114 18864
rect 11426 19388 11428 19408
rect 11428 19388 11480 19408
rect 11480 19388 11482 19408
rect 11426 19352 11482 19388
rect 10966 16088 11022 16144
rect 10966 15972 11022 16008
rect 10966 15952 10968 15972
rect 10968 15952 11020 15972
rect 11020 15952 11022 15972
rect 10322 14728 10378 14784
rect 10322 12552 10378 12608
rect 10782 15272 10838 15328
rect 10690 12844 10746 12880
rect 10690 12824 10692 12844
rect 10692 12824 10744 12844
rect 10744 12824 10746 12844
rect 10966 12552 11022 12608
rect 11518 18944 11574 19000
rect 11518 18672 11574 18728
rect 12254 21256 12310 21312
rect 12622 23024 12678 23080
rect 11794 20576 11850 20632
rect 11794 19760 11850 19816
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12714 22752 12770 22808
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 13726 23296 13782 23352
rect 13910 23060 13912 23080
rect 13912 23060 13964 23080
rect 13964 23060 13966 23080
rect 13910 23024 13966 23060
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12530 20168 12586 20224
rect 12438 19488 12494 19544
rect 11518 17584 11574 17640
rect 11886 17992 11942 18048
rect 11886 17756 11888 17776
rect 11888 17756 11940 17776
rect 11940 17756 11942 17776
rect 11886 17720 11942 17756
rect 11518 16904 11574 16960
rect 11794 16632 11850 16688
rect 12070 15408 12126 15464
rect 11978 15020 12034 15056
rect 11978 15000 11980 15020
rect 11980 15000 12032 15020
rect 12032 15000 12034 15020
rect 11426 11464 11482 11520
rect 11518 11056 11574 11112
rect 11058 10512 11114 10568
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 11518 10512 11574 10568
rect 11426 9832 11482 9888
rect 11886 14456 11942 14512
rect 12530 17448 12586 17504
rect 12530 16904 12586 16960
rect 12254 15136 12310 15192
rect 12438 12688 12494 12744
rect 12254 11872 12310 11928
rect 11978 11328 12034 11384
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 13174 18536 13230 18592
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 13266 17756 13268 17776
rect 13268 17756 13320 17776
rect 13320 17756 13322 17776
rect 13266 17720 13322 17756
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13910 21120 13966 21176
rect 13910 20748 13912 20768
rect 13912 20748 13964 20768
rect 13964 20748 13966 20768
rect 13910 20712 13966 20748
rect 13818 20440 13874 20496
rect 13634 18536 13690 18592
rect 12806 16768 12862 16824
rect 13358 16768 13414 16824
rect 12990 16668 12992 16688
rect 12992 16668 13044 16688
rect 13044 16668 13046 16688
rect 12990 16632 13046 16668
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 13358 15680 13414 15736
rect 14462 23976 14518 24032
rect 14462 23432 14518 23488
rect 14370 23296 14426 23352
rect 14370 21956 14426 21992
rect 14370 21936 14372 21956
rect 14372 21936 14424 21956
rect 14424 21936 14426 21956
rect 14922 24248 14978 24304
rect 14922 23568 14978 23624
rect 14922 21956 14978 21992
rect 14922 21936 14924 21956
rect 14924 21936 14976 21956
rect 14976 21936 14978 21956
rect 14922 21392 14978 21448
rect 14830 20576 14886 20632
rect 13726 16940 13728 16960
rect 13728 16940 13780 16960
rect 13780 16940 13782 16960
rect 13726 16904 13782 16940
rect 12438 11736 12494 11792
rect 12346 11056 12402 11112
rect 12254 10784 12310 10840
rect 12070 9424 12126 9480
rect 13266 15136 13322 15192
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12898 14320 12954 14376
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13082 11736 13138 11792
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12898 10784 12954 10840
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 14462 18672 14518 18728
rect 14922 19252 14924 19272
rect 14924 19252 14976 19272
rect 14976 19252 14978 19272
rect 14922 19216 14978 19252
rect 14738 17992 14794 18048
rect 14462 17584 14518 17640
rect 14370 16496 14426 16552
rect 14002 13096 14058 13152
rect 13818 10784 13874 10840
rect 15014 18808 15070 18864
rect 15566 21412 15622 21448
rect 15566 21392 15568 21412
rect 15568 21392 15620 21412
rect 15620 21392 15622 21412
rect 15750 21528 15806 21584
rect 16026 23704 16082 23760
rect 16210 25200 16266 25256
rect 15382 19216 15438 19272
rect 15566 19216 15622 19272
rect 15198 18400 15254 18456
rect 15750 18944 15806 19000
rect 15934 21564 15936 21584
rect 15936 21564 15988 21584
rect 15988 21564 15990 21584
rect 15934 21528 15990 21564
rect 16946 22616 17002 22672
rect 16578 21256 16634 21312
rect 16118 19488 16174 19544
rect 15382 15816 15438 15872
rect 15566 14728 15622 14784
rect 15290 13096 15346 13152
rect 15198 12552 15254 12608
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 14738 9460 14740 9480
rect 14740 9460 14792 9480
rect 14792 9460 14794 9480
rect 14738 9424 14794 9460
rect 16578 19116 16580 19136
rect 16580 19116 16632 19136
rect 16632 19116 16634 19136
rect 16578 19080 16634 19116
rect 16394 18264 16450 18320
rect 16578 16632 16634 16688
rect 15842 14320 15898 14376
rect 16210 14320 16266 14376
rect 15474 10240 15530 10296
rect 16578 15852 16580 15872
rect 16580 15852 16632 15872
rect 16632 15852 16634 15872
rect 16578 15816 16634 15852
rect 16486 11076 16542 11112
rect 16486 11056 16488 11076
rect 16488 11056 16540 11076
rect 16540 11056 16542 11076
rect 16578 10260 16634 10296
rect 16578 10240 16580 10260
rect 16580 10240 16632 10260
rect 16632 10240 16634 10260
rect 16946 20032 17002 20088
rect 16854 18944 16910 19000
rect 17038 18536 17094 18592
rect 16854 17992 16910 18048
rect 17222 22616 17278 22672
rect 17222 21800 17278 21856
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 18970 25200 19026 25256
rect 18418 24384 18474 24440
rect 18418 23976 18474 24032
rect 17406 20884 17408 20904
rect 17408 20884 17460 20904
rect 17460 20884 17462 20904
rect 17406 20848 17462 20884
rect 17222 19932 17224 19952
rect 17224 19932 17276 19952
rect 17276 19932 17278 19952
rect 17222 19896 17278 19932
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18418 21120 18474 21176
rect 17130 17856 17186 17912
rect 16946 16768 17002 16824
rect 16946 16360 17002 16416
rect 17130 16244 17186 16280
rect 17130 16224 17132 16244
rect 17132 16224 17184 16244
rect 17184 16224 17186 16244
rect 17406 19116 17408 19136
rect 17408 19116 17460 19136
rect 17460 19116 17462 19136
rect 17406 19080 17462 19116
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17774 19488 17830 19544
rect 17682 19080 17738 19136
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17590 18264 17646 18320
rect 18326 18264 18382 18320
rect 17130 14864 17186 14920
rect 17498 16360 17554 16416
rect 17498 15272 17554 15328
rect 17774 17720 17830 17776
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17774 16632 17830 16688
rect 18326 17040 18382 17096
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18602 18944 18658 19000
rect 18602 16632 18658 16688
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17314 11892 17370 11928
rect 17314 11872 17316 11892
rect 17316 11872 17368 11892
rect 17368 11872 17370 11892
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18878 18536 18934 18592
rect 18878 17856 18934 17912
rect 18970 16632 19026 16688
rect 18786 14728 18842 14784
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18602 12688 18658 12744
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 17590 9424 17646 9480
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 19246 22072 19302 22128
rect 19522 21972 19524 21992
rect 19524 21972 19576 21992
rect 19576 21972 19578 21992
rect 19522 21936 19578 21972
rect 19522 20032 19578 20088
rect 19246 18672 19302 18728
rect 19522 19216 19578 19272
rect 19522 18672 19578 18728
rect 19430 18400 19486 18456
rect 19338 16088 19394 16144
rect 19614 17176 19670 17232
rect 19522 15272 19578 15328
rect 19338 14864 19394 14920
rect 19154 12552 19210 12608
rect 19154 11192 19210 11248
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 20166 21936 20222 21992
rect 20718 24792 20774 24848
rect 20534 24384 20590 24440
rect 20166 21256 20222 21312
rect 20074 16904 20130 16960
rect 20166 16768 20222 16824
rect 20626 22208 20682 22264
rect 21178 24656 21234 24712
rect 21638 24248 21694 24304
rect 20534 17584 20590 17640
rect 19890 13912 19946 13968
rect 19614 12300 19670 12336
rect 19614 12280 19616 12300
rect 19616 12280 19668 12300
rect 19668 12280 19670 12300
rect 20718 14356 20720 14376
rect 20720 14356 20772 14376
rect 20772 14356 20774 14376
rect 20718 14320 20774 14356
rect 21086 17992 21142 18048
rect 21362 17584 21418 17640
rect 21270 16632 21326 16688
rect 21454 16360 21510 16416
rect 21362 15544 21418 15600
rect 22006 23976 22062 24032
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22190 23160 22246 23216
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22926 21800 22982 21856
rect 23202 21664 23258 21720
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 24122 23024 24178 23080
rect 24030 22888 24086 22944
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22006 18400 22062 18456
rect 21086 12824 21142 12880
rect 22466 17992 22522 18048
rect 22098 15544 22154 15600
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22926 18400 22982 18456
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22282 15680 22338 15736
rect 22006 13232 22062 13288
rect 23386 18672 23442 18728
rect 23754 17876 23810 17912
rect 23754 17856 23756 17876
rect 23756 17856 23808 17876
rect 23808 17856 23810 17876
rect 23938 17176 23994 17232
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22926 15580 22928 15600
rect 22928 15580 22980 15600
rect 22980 15580 22982 15600
rect 22926 15544 22982 15580
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 23110 13252 23166 13288
rect 23110 13232 23112 13252
rect 23112 13232 23164 13252
rect 23164 13232 23166 13252
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 24214 20712 24270 20768
rect 24122 16360 24178 16416
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 24766 23432 24822 23488
rect 24398 21664 24454 21720
rect 26514 23840 26570 23896
rect 25042 21800 25098 21856
rect 25686 20712 25742 20768
rect 24766 20304 24822 20360
rect 24398 18536 24454 18592
rect 25410 18672 25466 18728
rect 26238 18828 26294 18864
rect 26238 18808 26240 18828
rect 26240 18808 26292 18828
rect 26292 18808 26294 18828
rect 25962 17176 26018 17232
rect 25686 16632 25742 16688
rect 25042 12280 25098 12336
rect 25594 15308 25596 15328
rect 25596 15308 25648 15328
rect 25648 15308 25650 15328
rect 25594 15272 25650 15308
rect 25226 13232 25282 13288
rect 24306 9016 24362 9072
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 26514 21664 26570 21720
rect 27342 22208 27398 22264
rect 26606 21256 26662 21312
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 28814 22380 28816 22400
rect 28816 22380 28868 22400
rect 28868 22380 28870 22400
rect 28814 22344 28870 22380
rect 28538 21936 28594 21992
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 26514 18808 26570 18864
rect 27434 19236 27490 19272
rect 27434 19216 27436 19236
rect 27436 19216 27488 19236
rect 27488 19216 27490 19236
rect 29734 23432 29790 23488
rect 30194 23296 30250 23352
rect 30562 23840 30618 23896
rect 30286 23044 30342 23080
rect 30286 23024 30288 23044
rect 30288 23024 30340 23044
rect 30340 23024 30342 23044
rect 28722 21256 28778 21312
rect 28630 20848 28686 20904
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27250 18400 27306 18456
rect 26514 16632 26570 16688
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 28538 16496 28594 16552
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27710 11600 27766 11656
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 30930 22344 30986 22400
rect 30930 22208 30986 22264
rect 29826 21664 29882 21720
rect 30102 20440 30158 20496
rect 29550 15952 29606 16008
rect 30654 19372 30710 19408
rect 30654 19352 30656 19372
rect 30656 19352 30708 19372
rect 30708 19352 30710 19372
rect 30654 17856 30710 17912
rect 29918 15408 29974 15464
rect 31298 24656 31354 24712
rect 31298 23316 31354 23352
rect 31298 23296 31300 23316
rect 31300 23296 31352 23316
rect 31352 23296 31354 23316
rect 31298 22344 31354 22400
rect 31114 22208 31170 22264
rect 31114 21392 31170 21448
rect 31206 18264 31262 18320
rect 31482 21664 31538 21720
rect 31666 23432 31722 23488
rect 31850 20984 31906 21040
rect 31850 19896 31906 19952
rect 32310 23840 32366 23896
rect 32494 22480 32550 22536
rect 32218 19760 32274 19816
rect 31942 17584 31998 17640
rect 30746 13368 30802 13424
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 33414 23704 33470 23760
rect 35070 24112 35126 24168
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32678 18128 32734 18184
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 33874 22636 33930 22672
rect 33874 22616 33876 22636
rect 33876 22616 33928 22636
rect 33928 22616 33930 22636
rect 33598 22072 33654 22128
rect 35990 24792 36046 24848
rect 34886 23196 34888 23216
rect 34888 23196 34940 23216
rect 34940 23196 34942 23216
rect 34886 23160 34942 23196
rect 35070 23060 35072 23080
rect 35072 23060 35124 23080
rect 35124 23060 35126 23080
rect 35070 23024 35126 23060
rect 33322 15000 33378 15056
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 36174 21528 36230 21584
rect 38658 24928 38714 24984
rect 40130 24268 40186 24304
rect 40130 24248 40132 24268
rect 40132 24248 40184 24268
rect 40184 24248 40186 24268
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 45742 18808 45798 18864
rect 45374 18672 45430 18728
rect 46846 17176 46902 17232
rect 48318 24792 48374 24848
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 48226 23704 48282 23760
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 49054 22888 49110 22944
rect 49054 21972 49056 21992
rect 49056 21972 49108 21992
rect 49108 21972 49110 21992
rect 49054 21936 49110 21972
rect 49146 20984 49202 21040
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 0 25666 800 25696
rect 3785 25666 3851 25669
rect 0 25664 3851 25666
rect 0 25608 3790 25664
rect 3846 25608 3851 25664
rect 0 25606 3851 25608
rect 0 25576 800 25606
rect 3785 25603 3851 25606
rect 0 25258 800 25288
rect 3693 25258 3759 25261
rect 0 25256 3759 25258
rect 0 25200 3698 25256
rect 3754 25200 3759 25256
rect 0 25198 3759 25200
rect 0 25168 800 25198
rect 3693 25195 3759 25198
rect 16205 25258 16271 25261
rect 18965 25258 19031 25261
rect 16205 25256 19031 25258
rect 16205 25200 16210 25256
rect 16266 25200 18970 25256
rect 19026 25200 19031 25256
rect 16205 25198 19031 25200
rect 16205 25195 16271 25198
rect 18965 25195 19031 25198
rect 16982 24924 16988 24988
rect 17052 24986 17058 24988
rect 38653 24986 38719 24989
rect 17052 24984 38719 24986
rect 17052 24928 38658 24984
rect 38714 24928 38719 24984
rect 17052 24926 38719 24928
rect 17052 24924 17058 24926
rect 38653 24923 38719 24926
rect 0 24850 800 24880
rect 3049 24850 3115 24853
rect 0 24848 3115 24850
rect 0 24792 3054 24848
rect 3110 24792 3115 24848
rect 0 24790 3115 24792
rect 0 24760 800 24790
rect 3049 24787 3115 24790
rect 20713 24850 20779 24853
rect 35985 24850 36051 24853
rect 20713 24848 36051 24850
rect 20713 24792 20718 24848
rect 20774 24792 35990 24848
rect 36046 24792 36051 24848
rect 20713 24790 36051 24792
rect 20713 24787 20779 24790
rect 35985 24787 36051 24790
rect 48313 24850 48379 24853
rect 50200 24850 51000 24880
rect 48313 24848 51000 24850
rect 48313 24792 48318 24848
rect 48374 24792 51000 24848
rect 48313 24790 51000 24792
rect 48313 24787 48379 24790
rect 50200 24760 51000 24790
rect 4797 24714 4863 24717
rect 21173 24714 21239 24717
rect 31293 24714 31359 24717
rect 4797 24712 21239 24714
rect 4797 24656 4802 24712
rect 4858 24656 21178 24712
rect 21234 24656 21239 24712
rect 4797 24654 21239 24656
rect 4797 24651 4863 24654
rect 21173 24651 21239 24654
rect 22050 24712 31359 24714
rect 22050 24656 31298 24712
rect 31354 24656 31359 24712
rect 22050 24654 31359 24656
rect 14406 24516 14412 24580
rect 14476 24578 14482 24580
rect 22050 24578 22110 24654
rect 31293 24651 31359 24654
rect 14476 24518 22110 24578
rect 14476 24516 14482 24518
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 2773 24442 2839 24445
rect 18413 24442 18479 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 14782 24440 18479 24442
rect 14782 24384 18418 24440
rect 18474 24384 18479 24440
rect 14782 24382 18479 24384
rect 9673 24306 9739 24309
rect 14782 24306 14842 24382
rect 18413 24379 18479 24382
rect 20529 24442 20595 24445
rect 20529 24440 22110 24442
rect 20529 24384 20534 24440
rect 20590 24384 22110 24440
rect 20529 24382 22110 24384
rect 20529 24379 20595 24382
rect 9673 24304 14842 24306
rect 9673 24248 9678 24304
rect 9734 24248 14842 24304
rect 9673 24246 14842 24248
rect 14917 24306 14983 24309
rect 21633 24306 21699 24309
rect 14917 24304 21699 24306
rect 14917 24248 14922 24304
rect 14978 24248 21638 24304
rect 21694 24248 21699 24304
rect 14917 24246 21699 24248
rect 22050 24306 22110 24382
rect 40125 24306 40191 24309
rect 22050 24304 40191 24306
rect 22050 24248 40130 24304
rect 40186 24248 40191 24304
rect 22050 24246 40191 24248
rect 9673 24243 9739 24246
rect 14917 24243 14983 24246
rect 21633 24243 21699 24246
rect 40125 24243 40191 24246
rect 4245 24170 4311 24173
rect 5574 24170 5580 24172
rect 4245 24168 5580 24170
rect 4245 24112 4250 24168
rect 4306 24112 5580 24168
rect 4245 24110 5580 24112
rect 4245 24107 4311 24110
rect 5574 24108 5580 24110
rect 5644 24108 5650 24172
rect 8753 24170 8819 24173
rect 35065 24170 35131 24173
rect 8753 24168 35131 24170
rect 8753 24112 8758 24168
rect 8814 24112 35070 24168
rect 35126 24112 35131 24168
rect 8753 24110 35131 24112
rect 8753 24107 8819 24110
rect 35065 24107 35131 24110
rect 0 24034 800 24064
rect 4061 24034 4127 24037
rect 0 24032 4127 24034
rect 0 23976 4066 24032
rect 4122 23976 4127 24032
rect 0 23974 4127 23976
rect 0 23944 800 23974
rect 4061 23971 4127 23974
rect 11789 24034 11855 24037
rect 14457 24034 14523 24037
rect 11789 24032 14523 24034
rect 11789 23976 11794 24032
rect 11850 23976 14462 24032
rect 14518 23976 14523 24032
rect 11789 23974 14523 23976
rect 11789 23971 11855 23974
rect 14457 23971 14523 23974
rect 18413 24034 18479 24037
rect 22001 24034 22067 24037
rect 18413 24032 22067 24034
rect 18413 23976 18418 24032
rect 18474 23976 22006 24032
rect 22062 23976 22067 24032
rect 18413 23974 22067 23976
rect 18413 23971 18479 23974
rect 22001 23971 22067 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 26509 23898 26575 23901
rect 18462 23896 26575 23898
rect 18462 23840 26514 23896
rect 26570 23840 26575 23896
rect 18462 23838 26575 23840
rect 12341 23762 12407 23765
rect 16021 23762 16087 23765
rect 18462 23762 18522 23838
rect 26509 23835 26575 23838
rect 30557 23898 30623 23901
rect 32305 23898 32371 23901
rect 50200 23898 51000 23928
rect 30557 23896 32371 23898
rect 30557 23840 30562 23896
rect 30618 23840 32310 23896
rect 32366 23840 32371 23896
rect 30557 23838 32371 23840
rect 30557 23835 30623 23838
rect 32305 23835 32371 23838
rect 48454 23838 51000 23898
rect 33409 23762 33475 23765
rect 12341 23760 15210 23762
rect 12341 23704 12346 23760
rect 12402 23704 15210 23760
rect 12341 23702 15210 23704
rect 12341 23699 12407 23702
rect 0 23626 800 23656
rect 3877 23626 3943 23629
rect 0 23624 3943 23626
rect 0 23568 3882 23624
rect 3938 23568 3943 23624
rect 0 23566 3943 23568
rect 0 23536 800 23566
rect 3877 23563 3943 23566
rect 4286 23564 4292 23628
rect 4356 23626 4362 23628
rect 7097 23626 7163 23629
rect 4356 23624 7163 23626
rect 4356 23568 7102 23624
rect 7158 23568 7163 23624
rect 4356 23566 7163 23568
rect 4356 23564 4362 23566
rect 7097 23563 7163 23566
rect 12065 23626 12131 23629
rect 14917 23626 14983 23629
rect 12065 23624 14983 23626
rect 12065 23568 12070 23624
rect 12126 23568 14922 23624
rect 14978 23568 14983 23624
rect 12065 23566 14983 23568
rect 15150 23626 15210 23702
rect 16021 23760 18522 23762
rect 16021 23704 16026 23760
rect 16082 23704 18522 23760
rect 16021 23702 18522 23704
rect 22050 23760 33475 23762
rect 22050 23704 33414 23760
rect 33470 23704 33475 23760
rect 22050 23702 33475 23704
rect 16021 23699 16087 23702
rect 22050 23626 22110 23702
rect 33409 23699 33475 23702
rect 48221 23762 48287 23765
rect 48454 23762 48514 23838
rect 50200 23808 51000 23838
rect 48221 23760 48514 23762
rect 48221 23704 48226 23760
rect 48282 23704 48514 23760
rect 48221 23702 48514 23704
rect 48221 23699 48287 23702
rect 15150 23566 22110 23626
rect 22694 23566 23490 23626
rect 12065 23563 12131 23566
rect 14917 23563 14983 23566
rect 2129 23490 2195 23493
rect 2262 23490 2268 23492
rect 2129 23488 2268 23490
rect 2129 23432 2134 23488
rect 2190 23432 2268 23488
rect 2129 23430 2268 23432
rect 2129 23427 2195 23430
rect 2262 23428 2268 23430
rect 2332 23428 2338 23492
rect 5390 23428 5396 23492
rect 5460 23490 5466 23492
rect 6545 23490 6611 23493
rect 5460 23488 6611 23490
rect 5460 23432 6550 23488
rect 6606 23432 6611 23488
rect 5460 23430 6611 23432
rect 5460 23428 5466 23430
rect 6545 23427 6611 23430
rect 7598 23428 7604 23492
rect 7668 23490 7674 23492
rect 7925 23490 7991 23493
rect 7668 23488 7991 23490
rect 7668 23432 7930 23488
rect 7986 23432 7991 23488
rect 7668 23430 7991 23432
rect 7668 23428 7674 23430
rect 7925 23427 7991 23430
rect 14457 23490 14523 23493
rect 22694 23490 22754 23566
rect 14457 23488 22754 23490
rect 14457 23432 14462 23488
rect 14518 23432 22754 23488
rect 14457 23430 22754 23432
rect 23430 23490 23490 23566
rect 24761 23490 24827 23493
rect 23430 23488 24827 23490
rect 23430 23432 24766 23488
rect 24822 23432 24827 23488
rect 23430 23430 24827 23432
rect 14457 23427 14523 23430
rect 24761 23427 24827 23430
rect 29729 23490 29795 23493
rect 31661 23490 31727 23493
rect 29729 23488 31727 23490
rect 29729 23432 29734 23488
rect 29790 23432 31666 23488
rect 31722 23432 31727 23488
rect 29729 23430 31727 23432
rect 29729 23427 29795 23430
rect 31661 23427 31727 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 13721 23354 13787 23357
rect 14365 23354 14431 23357
rect 30189 23354 30255 23357
rect 31293 23354 31359 23357
rect 13721 23352 22754 23354
rect 13721 23296 13726 23352
rect 13782 23296 14370 23352
rect 14426 23296 22754 23352
rect 13721 23294 22754 23296
rect 13721 23291 13787 23294
rect 14365 23291 14431 23294
rect 0 23218 800 23248
rect 3693 23218 3759 23221
rect 22185 23220 22251 23221
rect 0 23216 3759 23218
rect 0 23160 3698 23216
rect 3754 23160 3759 23216
rect 0 23158 3759 23160
rect 0 23128 800 23158
rect 3693 23155 3759 23158
rect 5574 23156 5580 23220
rect 5644 23218 5650 23220
rect 22134 23218 22140 23220
rect 5644 23158 18706 23218
rect 22094 23158 22140 23218
rect 22204 23216 22251 23220
rect 22246 23160 22251 23216
rect 5644 23156 5650 23158
rect 3601 23082 3667 23085
rect 12617 23082 12683 23085
rect 3601 23080 12683 23082
rect 3601 23024 3606 23080
rect 3662 23024 12622 23080
rect 12678 23024 12683 23080
rect 3601 23022 12683 23024
rect 3601 23019 3667 23022
rect 12617 23019 12683 23022
rect 13905 23082 13971 23085
rect 18646 23082 18706 23158
rect 22134 23156 22140 23158
rect 22204 23156 22251 23160
rect 22694 23218 22754 23294
rect 30189 23352 31359 23354
rect 30189 23296 30194 23352
rect 30250 23296 31298 23352
rect 31354 23296 31359 23352
rect 30189 23294 31359 23296
rect 30189 23291 30255 23294
rect 31293 23291 31359 23294
rect 34881 23218 34947 23221
rect 22694 23216 34947 23218
rect 22694 23160 34886 23216
rect 34942 23160 34947 23216
rect 22694 23158 34947 23160
rect 22185 23155 22251 23156
rect 34881 23155 34947 23158
rect 24117 23082 24183 23085
rect 13905 23080 18522 23082
rect 13905 23024 13910 23080
rect 13966 23024 18522 23080
rect 13905 23022 18522 23024
rect 18646 23080 24183 23082
rect 18646 23024 24122 23080
rect 24178 23024 24183 23080
rect 18646 23022 24183 23024
rect 13905 23019 13971 23022
rect 4521 22946 4587 22949
rect 4654 22946 4660 22948
rect 4521 22944 4660 22946
rect 4521 22888 4526 22944
rect 4582 22888 4660 22944
rect 4521 22886 4660 22888
rect 4521 22883 4587 22886
rect 4654 22884 4660 22886
rect 4724 22884 4730 22948
rect 18462 22946 18522 23022
rect 24117 23019 24183 23022
rect 30281 23082 30347 23085
rect 35065 23082 35131 23085
rect 30281 23080 35131 23082
rect 30281 23024 30286 23080
rect 30342 23024 35070 23080
rect 35126 23024 35131 23080
rect 30281 23022 35131 23024
rect 30281 23019 30347 23022
rect 35065 23019 35131 23022
rect 24025 22946 24091 22949
rect 18462 22944 24091 22946
rect 18462 22888 24030 22944
rect 24086 22888 24091 22944
rect 18462 22886 24091 22888
rect 24025 22883 24091 22886
rect 49049 22946 49115 22949
rect 50200 22946 51000 22976
rect 49049 22944 51000 22946
rect 49049 22888 49054 22944
rect 49110 22888 51000 22944
rect 49049 22886 51000 22888
rect 49049 22883 49115 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 50200 22856 51000 22886
rect 47946 22815 48262 22816
rect 4981 22810 5047 22813
rect 0 22808 5047 22810
rect 0 22752 4986 22808
rect 5042 22752 5047 22808
rect 0 22750 5047 22752
rect 0 22720 800 22750
rect 4981 22747 5047 22750
rect 12709 22810 12775 22813
rect 17166 22810 17172 22812
rect 12709 22808 17172 22810
rect 12709 22752 12714 22808
rect 12770 22752 17172 22808
rect 12709 22750 17172 22752
rect 12709 22747 12775 22750
rect 17166 22748 17172 22750
rect 17236 22748 17242 22812
rect 16941 22674 17007 22677
rect 17217 22674 17283 22677
rect 33869 22674 33935 22677
rect 16941 22672 33935 22674
rect 16941 22616 16946 22672
rect 17002 22616 17222 22672
rect 17278 22616 33874 22672
rect 33930 22616 33935 22672
rect 16941 22614 33935 22616
rect 16941 22611 17007 22614
rect 17217 22611 17283 22614
rect 33869 22611 33935 22614
rect 4153 22540 4219 22541
rect 4102 22538 4108 22540
rect 4062 22478 4108 22538
rect 4172 22536 4219 22540
rect 4214 22480 4219 22536
rect 4102 22476 4108 22478
rect 4172 22476 4219 22480
rect 17166 22476 17172 22540
rect 17236 22538 17242 22540
rect 32489 22538 32555 22541
rect 17236 22536 32555 22538
rect 17236 22480 32494 22536
rect 32550 22480 32555 22536
rect 17236 22478 32555 22480
rect 17236 22476 17242 22478
rect 4153 22475 4219 22476
rect 32489 22475 32555 22478
rect 0 22402 800 22432
rect 2129 22402 2195 22405
rect 0 22400 2195 22402
rect 0 22344 2134 22400
rect 2190 22344 2195 22400
rect 0 22342 2195 22344
rect 0 22312 800 22342
rect 2129 22339 2195 22342
rect 28809 22402 28875 22405
rect 30925 22402 30991 22405
rect 31293 22402 31359 22405
rect 28809 22400 31359 22402
rect 28809 22344 28814 22400
rect 28870 22344 30930 22400
rect 30986 22344 31298 22400
rect 31354 22344 31359 22400
rect 28809 22342 31359 22344
rect 28809 22339 28875 22342
rect 30925 22339 30991 22342
rect 31293 22339 31359 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 20621 22266 20687 22269
rect 27337 22266 27403 22269
rect 30925 22266 30991 22269
rect 31109 22266 31175 22269
rect 20621 22264 22110 22266
rect 20621 22208 20626 22264
rect 20682 22208 22110 22264
rect 20621 22206 22110 22208
rect 20621 22203 20687 22206
rect 6637 22132 6703 22133
rect 6637 22130 6684 22132
rect 6556 22128 6684 22130
rect 6748 22130 6754 22132
rect 19241 22130 19307 22133
rect 6748 22128 19307 22130
rect 6556 22072 6642 22128
rect 6748 22072 19246 22128
rect 19302 22072 19307 22128
rect 6556 22070 6684 22072
rect 6637 22068 6684 22070
rect 6748 22070 19307 22072
rect 22050 22130 22110 22206
rect 27337 22264 31175 22266
rect 27337 22208 27342 22264
rect 27398 22208 30930 22264
rect 30986 22208 31114 22264
rect 31170 22208 31175 22264
rect 27337 22206 31175 22208
rect 27337 22203 27403 22206
rect 30925 22203 30991 22206
rect 31109 22203 31175 22206
rect 33593 22130 33659 22133
rect 22050 22128 33659 22130
rect 22050 22072 33598 22128
rect 33654 22072 33659 22128
rect 22050 22070 33659 22072
rect 6748 22068 6754 22070
rect 6637 22067 6703 22068
rect 19241 22067 19307 22070
rect 33593 22067 33659 22070
rect 0 21994 800 22024
rect 4613 21994 4679 21997
rect 9305 21994 9371 21997
rect 0 21992 4679 21994
rect 0 21936 4618 21992
rect 4674 21936 4679 21992
rect 0 21934 4679 21936
rect 0 21904 800 21934
rect 4613 21931 4679 21934
rect 7790 21992 9371 21994
rect 7790 21936 9310 21992
rect 9366 21936 9371 21992
rect 7790 21934 9371 21936
rect 1669 21858 1735 21861
rect 7790 21858 7850 21934
rect 9305 21931 9371 21934
rect 9489 21994 9555 21997
rect 14365 21996 14431 21997
rect 14365 21994 14412 21996
rect 9489 21992 14412 21994
rect 14476 21994 14482 21996
rect 14917 21994 14983 21997
rect 19517 21994 19583 21997
rect 9489 21936 9494 21992
rect 9550 21936 14370 21992
rect 9489 21934 14412 21936
rect 9489 21931 9555 21934
rect 14365 21932 14412 21934
rect 14476 21934 14522 21994
rect 14917 21992 19583 21994
rect 14917 21936 14922 21992
rect 14978 21936 19522 21992
rect 19578 21936 19583 21992
rect 14917 21934 19583 21936
rect 14476 21932 14482 21934
rect 14365 21931 14431 21932
rect 14917 21931 14983 21934
rect 19517 21931 19583 21934
rect 20161 21994 20227 21997
rect 28533 21994 28599 21997
rect 20161 21992 28599 21994
rect 20161 21936 20166 21992
rect 20222 21936 28538 21992
rect 28594 21936 28599 21992
rect 20161 21934 28599 21936
rect 20161 21931 20227 21934
rect 28533 21931 28599 21934
rect 49049 21994 49115 21997
rect 50200 21994 51000 22024
rect 49049 21992 51000 21994
rect 49049 21936 49054 21992
rect 49110 21936 51000 21992
rect 49049 21934 51000 21936
rect 49049 21931 49115 21934
rect 50200 21904 51000 21934
rect 1669 21856 7850 21858
rect 1669 21800 1674 21856
rect 1730 21800 7850 21856
rect 1669 21798 7850 21800
rect 10961 21858 11027 21861
rect 17217 21858 17283 21861
rect 10961 21856 17283 21858
rect 10961 21800 10966 21856
rect 11022 21800 17222 21856
rect 17278 21800 17283 21856
rect 10961 21798 17283 21800
rect 1669 21795 1735 21798
rect 10961 21795 11027 21798
rect 17217 21795 17283 21798
rect 22921 21858 22987 21861
rect 25037 21858 25103 21861
rect 22921 21856 25103 21858
rect 22921 21800 22926 21856
rect 22982 21800 25042 21856
rect 25098 21800 25103 21856
rect 22921 21798 25103 21800
rect 22921 21795 22987 21798
rect 25037 21795 25103 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 3969 21724 4035 21725
rect 3918 21660 3924 21724
rect 3988 21722 4035 21724
rect 3988 21720 4080 21722
rect 4030 21664 4080 21720
rect 3988 21662 4080 21664
rect 3988 21660 4035 21662
rect 22686 21660 22692 21724
rect 22756 21722 22762 21724
rect 23197 21722 23263 21725
rect 22756 21720 23263 21722
rect 22756 21664 23202 21720
rect 23258 21664 23263 21720
rect 22756 21662 23263 21664
rect 22756 21660 22762 21662
rect 3969 21659 4035 21660
rect 23197 21659 23263 21662
rect 24393 21722 24459 21725
rect 26509 21722 26575 21725
rect 24393 21720 26575 21722
rect 24393 21664 24398 21720
rect 24454 21664 26514 21720
rect 26570 21664 26575 21720
rect 24393 21662 26575 21664
rect 24393 21659 24459 21662
rect 26509 21659 26575 21662
rect 29821 21722 29887 21725
rect 31477 21722 31543 21725
rect 29821 21720 31543 21722
rect 29821 21664 29826 21720
rect 29882 21664 31482 21720
rect 31538 21664 31543 21720
rect 29821 21662 31543 21664
rect 29821 21659 29887 21662
rect 31477 21659 31543 21662
rect 0 21586 800 21616
rect 2957 21586 3023 21589
rect 0 21584 3023 21586
rect 0 21528 2962 21584
rect 3018 21528 3023 21584
rect 0 21526 3023 21528
rect 0 21496 800 21526
rect 2957 21523 3023 21526
rect 6177 21586 6243 21589
rect 8017 21586 8083 21589
rect 6177 21584 8083 21586
rect 6177 21528 6182 21584
rect 6238 21528 8022 21584
rect 8078 21528 8083 21584
rect 6177 21526 8083 21528
rect 6177 21523 6243 21526
rect 8017 21523 8083 21526
rect 8201 21586 8267 21589
rect 15745 21586 15811 21589
rect 8201 21584 15811 21586
rect 8201 21528 8206 21584
rect 8262 21528 15750 21584
rect 15806 21528 15811 21584
rect 8201 21526 15811 21528
rect 8201 21523 8267 21526
rect 15745 21523 15811 21526
rect 15929 21586 15995 21589
rect 36169 21586 36235 21589
rect 15929 21584 36235 21586
rect 15929 21528 15934 21584
rect 15990 21528 36174 21584
rect 36230 21528 36235 21584
rect 15929 21526 36235 21528
rect 15929 21523 15995 21526
rect 36169 21523 36235 21526
rect 3601 21450 3667 21453
rect 10501 21450 10567 21453
rect 14917 21450 14983 21453
rect 3601 21448 10567 21450
rect 3601 21392 3606 21448
rect 3662 21392 10506 21448
rect 10562 21392 10567 21448
rect 3601 21390 10567 21392
rect 3601 21387 3667 21390
rect 10501 21387 10567 21390
rect 12390 21448 14983 21450
rect 12390 21392 14922 21448
rect 14978 21392 14983 21448
rect 12390 21390 14983 21392
rect 5625 21314 5691 21317
rect 5942 21314 5948 21316
rect 5625 21312 5948 21314
rect 5625 21256 5630 21312
rect 5686 21256 5948 21312
rect 5625 21254 5948 21256
rect 5625 21251 5691 21254
rect 5942 21252 5948 21254
rect 6012 21252 6018 21316
rect 7373 21314 7439 21317
rect 12249 21314 12315 21317
rect 7373 21312 12315 21314
rect 7373 21256 7378 21312
rect 7434 21256 12254 21312
rect 12310 21256 12315 21312
rect 7373 21254 12315 21256
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 5950 21178 6010 21252
rect 7373 21251 7439 21254
rect 12249 21251 12315 21254
rect 12390 21178 12450 21390
rect 14917 21387 14983 21390
rect 15561 21450 15627 21453
rect 31109 21450 31175 21453
rect 15561 21448 31175 21450
rect 15561 21392 15566 21448
rect 15622 21392 31114 21448
rect 31170 21392 31175 21448
rect 15561 21390 31175 21392
rect 15561 21387 15627 21390
rect 31109 21387 31175 21390
rect 16573 21314 16639 21317
rect 20161 21314 20227 21317
rect 16573 21312 20227 21314
rect 16573 21256 16578 21312
rect 16634 21256 20166 21312
rect 20222 21256 20227 21312
rect 16573 21254 20227 21256
rect 16573 21251 16639 21254
rect 20161 21251 20227 21254
rect 26601 21314 26667 21317
rect 28717 21314 28783 21317
rect 26601 21312 28783 21314
rect 26601 21256 26606 21312
rect 26662 21256 28722 21312
rect 28778 21256 28783 21312
rect 26601 21254 28783 21256
rect 26601 21251 26667 21254
rect 28717 21251 28783 21254
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 5950 21118 12450 21178
rect 13905 21178 13971 21181
rect 18413 21178 18479 21181
rect 13905 21176 18479 21178
rect 13905 21120 13910 21176
rect 13966 21120 18418 21176
rect 18474 21120 18479 21176
rect 13905 21118 18479 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 13905 21115 13971 21118
rect 18413 21115 18479 21118
rect 4245 21042 4311 21045
rect 31845 21042 31911 21045
rect 4245 21040 31911 21042
rect 4245 20984 4250 21040
rect 4306 20984 31850 21040
rect 31906 20984 31911 21040
rect 4245 20982 31911 20984
rect 4245 20979 4311 20982
rect 31845 20979 31911 20982
rect 49141 21042 49207 21045
rect 50200 21042 51000 21072
rect 49141 21040 51000 21042
rect 49141 20984 49146 21040
rect 49202 20984 51000 21040
rect 49141 20982 51000 20984
rect 49141 20979 49207 20982
rect 50200 20952 51000 20982
rect 4061 20906 4127 20909
rect 11421 20906 11487 20909
rect 4061 20904 11487 20906
rect 4061 20848 4066 20904
rect 4122 20848 11426 20904
rect 11482 20848 11487 20904
rect 4061 20846 11487 20848
rect 4061 20843 4127 20846
rect 11421 20843 11487 20846
rect 17401 20906 17467 20909
rect 28625 20906 28691 20909
rect 17401 20904 28691 20906
rect 17401 20848 17406 20904
rect 17462 20848 28630 20904
rect 28686 20848 28691 20904
rect 17401 20846 28691 20848
rect 17401 20843 17467 20846
rect 28625 20843 28691 20846
rect 0 20770 800 20800
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 800 20710
rect 1301 20707 1367 20710
rect 5717 20772 5783 20773
rect 6913 20772 6979 20773
rect 5717 20768 5764 20772
rect 5828 20770 5834 20772
rect 6862 20770 6868 20772
rect 5717 20712 5722 20768
rect 5717 20708 5764 20712
rect 5828 20710 5874 20770
rect 6822 20710 6868 20770
rect 6932 20768 6979 20772
rect 6974 20712 6979 20768
rect 5828 20708 5834 20710
rect 6862 20708 6868 20710
rect 6932 20708 6979 20712
rect 7046 20708 7052 20772
rect 7116 20770 7122 20772
rect 7189 20770 7255 20773
rect 7116 20768 7255 20770
rect 7116 20712 7194 20768
rect 7250 20712 7255 20768
rect 7116 20710 7255 20712
rect 7116 20708 7122 20710
rect 5717 20707 5783 20708
rect 6913 20707 6979 20708
rect 7189 20707 7255 20710
rect 9673 20770 9739 20773
rect 10542 20770 10548 20772
rect 9673 20768 10548 20770
rect 9673 20712 9678 20768
rect 9734 20712 10548 20768
rect 9673 20710 10548 20712
rect 9673 20707 9739 20710
rect 10542 20708 10548 20710
rect 10612 20708 10618 20772
rect 11094 20708 11100 20772
rect 11164 20770 11170 20772
rect 11329 20770 11395 20773
rect 13905 20772 13971 20773
rect 11164 20768 11395 20770
rect 11164 20712 11334 20768
rect 11390 20712 11395 20768
rect 11164 20710 11395 20712
rect 11164 20708 11170 20710
rect 11329 20707 11395 20710
rect 13854 20708 13860 20772
rect 13924 20770 13971 20772
rect 24209 20770 24275 20773
rect 25681 20770 25747 20773
rect 13924 20768 14016 20770
rect 13966 20712 14016 20768
rect 13924 20710 14016 20712
rect 24209 20768 25747 20770
rect 24209 20712 24214 20768
rect 24270 20712 25686 20768
rect 25742 20712 25747 20768
rect 24209 20710 25747 20712
rect 13924 20708 13971 20710
rect 13905 20707 13971 20708
rect 24209 20707 24275 20710
rect 25681 20707 25747 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 9305 20634 9371 20637
rect 11789 20634 11855 20637
rect 14825 20634 14891 20637
rect 9305 20632 14891 20634
rect 9305 20576 9310 20632
rect 9366 20576 11794 20632
rect 11850 20576 14830 20632
rect 14886 20576 14891 20632
rect 9305 20574 14891 20576
rect 9305 20571 9371 20574
rect 11789 20571 11855 20574
rect 14825 20571 14891 20574
rect 13813 20498 13879 20501
rect 30097 20498 30163 20501
rect 13813 20496 30163 20498
rect 13813 20440 13818 20496
rect 13874 20440 30102 20496
rect 30158 20440 30163 20496
rect 13813 20438 30163 20440
rect 13813 20435 13879 20438
rect 30097 20435 30163 20438
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 6085 20362 6151 20365
rect 6453 20362 6519 20365
rect 24761 20362 24827 20365
rect 6085 20360 24827 20362
rect 6085 20304 6090 20360
rect 6146 20304 6458 20360
rect 6514 20304 24766 20360
rect 24822 20304 24827 20360
rect 6085 20302 24827 20304
rect 6085 20299 6151 20302
rect 6453 20299 6519 20302
rect 24761 20299 24827 20302
rect 9213 20226 9279 20229
rect 12525 20226 12591 20229
rect 9213 20224 12591 20226
rect 9213 20168 9218 20224
rect 9274 20168 12530 20224
rect 12586 20168 12591 20224
rect 9213 20166 12591 20168
rect 9213 20163 9279 20166
rect 12525 20163 12591 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 16941 20090 17007 20093
rect 19517 20090 19583 20093
rect 16941 20088 19583 20090
rect 16941 20032 16946 20088
rect 17002 20032 19522 20088
rect 19578 20032 19583 20088
rect 16941 20030 19583 20032
rect 16941 20027 17007 20030
rect 19517 20027 19583 20030
rect 0 19954 800 19984
rect 2037 19954 2103 19957
rect 0 19952 2103 19954
rect 0 19896 2042 19952
rect 2098 19896 2103 19952
rect 0 19894 2103 19896
rect 0 19864 800 19894
rect 2037 19891 2103 19894
rect 6729 19954 6795 19957
rect 8569 19954 8635 19957
rect 6729 19952 8635 19954
rect 6729 19896 6734 19952
rect 6790 19896 8574 19952
rect 8630 19896 8635 19952
rect 6729 19894 8635 19896
rect 6729 19891 6795 19894
rect 8569 19891 8635 19894
rect 17217 19954 17283 19957
rect 31845 19954 31911 19957
rect 17217 19952 31911 19954
rect 17217 19896 17222 19952
rect 17278 19896 31850 19952
rect 31906 19896 31911 19952
rect 17217 19894 31911 19896
rect 17217 19891 17283 19894
rect 31845 19891 31911 19894
rect 11789 19818 11855 19821
rect 32213 19818 32279 19821
rect 11789 19816 32279 19818
rect 11789 19760 11794 19816
rect 11850 19760 32218 19816
rect 32274 19760 32279 19816
rect 11789 19758 32279 19760
rect 11789 19755 11855 19758
rect 32213 19755 32279 19758
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 2773 19546 2839 19549
rect 3601 19546 3667 19549
rect 0 19544 2839 19546
rect 0 19488 2778 19544
rect 2834 19488 2839 19544
rect 0 19486 2839 19488
rect 0 19456 800 19486
rect 2773 19483 2839 19486
rect 3558 19544 3667 19546
rect 3558 19488 3606 19544
rect 3662 19488 3667 19544
rect 3558 19483 3667 19488
rect 10869 19546 10935 19549
rect 12433 19546 12499 19549
rect 10869 19544 12499 19546
rect 10869 19488 10874 19544
rect 10930 19488 12438 19544
rect 12494 19488 12499 19544
rect 10869 19486 12499 19488
rect 10869 19483 10935 19486
rect 12433 19483 12499 19486
rect 16113 19546 16179 19549
rect 17769 19546 17835 19549
rect 16113 19544 17835 19546
rect 16113 19488 16118 19544
rect 16174 19488 17774 19544
rect 17830 19488 17835 19544
rect 16113 19486 17835 19488
rect 16113 19483 16179 19486
rect 17769 19483 17835 19486
rect 2957 19274 3023 19277
rect 2730 19272 3023 19274
rect 2730 19216 2962 19272
rect 3018 19216 3023 19272
rect 2730 19214 3023 19216
rect 0 19138 800 19168
rect 2730 19138 2790 19214
rect 2957 19211 3023 19214
rect 0 19078 2790 19138
rect 0 19048 800 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 3558 19002 3618 19483
rect 5257 19410 5323 19413
rect 7465 19410 7531 19413
rect 5257 19408 7531 19410
rect 5257 19352 5262 19408
rect 5318 19352 7470 19408
rect 7526 19352 7531 19408
rect 5257 19350 7531 19352
rect 5257 19347 5323 19350
rect 7465 19347 7531 19350
rect 8753 19410 8819 19413
rect 9622 19410 9628 19412
rect 8753 19408 9628 19410
rect 8753 19352 8758 19408
rect 8814 19352 9628 19408
rect 8753 19350 9628 19352
rect 8753 19347 8819 19350
rect 9622 19348 9628 19350
rect 9692 19348 9698 19412
rect 11421 19410 11487 19413
rect 30649 19410 30715 19413
rect 11421 19408 30715 19410
rect 11421 19352 11426 19408
rect 11482 19352 30654 19408
rect 30710 19352 30715 19408
rect 11421 19350 30715 19352
rect 11421 19347 11487 19350
rect 30649 19347 30715 19350
rect 7414 19212 7420 19276
rect 7484 19274 7490 19276
rect 8293 19274 8359 19277
rect 7484 19272 8359 19274
rect 7484 19216 8298 19272
rect 8354 19216 8359 19272
rect 7484 19214 8359 19216
rect 7484 19212 7490 19214
rect 8293 19211 8359 19214
rect 10593 19274 10659 19277
rect 14917 19274 14983 19277
rect 10593 19272 14983 19274
rect 10593 19216 10598 19272
rect 10654 19216 14922 19272
rect 14978 19216 14983 19272
rect 10593 19214 14983 19216
rect 10593 19211 10659 19214
rect 14917 19211 14983 19214
rect 15377 19274 15443 19277
rect 15561 19274 15627 19277
rect 19517 19274 19583 19277
rect 27429 19274 27495 19277
rect 15377 19272 19583 19274
rect 15377 19216 15382 19272
rect 15438 19216 15566 19272
rect 15622 19216 19522 19272
rect 19578 19216 19583 19272
rect 15377 19214 19583 19216
rect 15377 19211 15443 19214
rect 15561 19211 15627 19214
rect 19517 19211 19583 19214
rect 22050 19272 27495 19274
rect 22050 19216 27434 19272
rect 27490 19216 27495 19272
rect 22050 19214 27495 19216
rect 4061 19138 4127 19141
rect 8569 19138 8635 19141
rect 4061 19136 8635 19138
rect 4061 19080 4066 19136
rect 4122 19080 8574 19136
rect 8630 19080 8635 19136
rect 4061 19078 8635 19080
rect 4061 19075 4127 19078
rect 8569 19075 8635 19078
rect 16573 19138 16639 19141
rect 17401 19138 17467 19141
rect 16573 19136 17467 19138
rect 16573 19080 16578 19136
rect 16634 19080 17406 19136
rect 17462 19080 17467 19136
rect 16573 19078 17467 19080
rect 16573 19075 16639 19078
rect 17401 19075 17467 19078
rect 17534 19076 17540 19140
rect 17604 19138 17610 19140
rect 17677 19138 17743 19141
rect 22050 19138 22110 19214
rect 27429 19211 27495 19214
rect 17604 19136 22110 19138
rect 17604 19080 17682 19136
rect 17738 19080 22110 19136
rect 17604 19078 22110 19080
rect 17604 19076 17610 19078
rect 17677 19075 17743 19078
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 3734 19002 3740 19004
rect 3558 18942 3740 19002
rect 3734 18940 3740 18942
rect 3804 19002 3810 19004
rect 11513 19002 11579 19005
rect 15745 19002 15811 19005
rect 3804 19000 11579 19002
rect 3804 18944 11518 19000
rect 11574 18944 11579 19000
rect 3804 18942 11579 18944
rect 3804 18940 3810 18942
rect 11513 18939 11579 18942
rect 14046 19000 15811 19002
rect 14046 18944 15750 19000
rect 15806 18944 15811 19000
rect 14046 18942 15811 18944
rect 4429 18866 4495 18869
rect 11053 18866 11119 18869
rect 14046 18866 14106 18942
rect 15745 18939 15811 18942
rect 16849 19002 16915 19005
rect 18597 19002 18663 19005
rect 16849 19000 18663 19002
rect 16849 18944 16854 19000
rect 16910 18944 18602 19000
rect 18658 18944 18663 19000
rect 16849 18942 18663 18944
rect 16849 18939 16915 18942
rect 18597 18939 18663 18942
rect 4429 18864 11119 18866
rect 4429 18808 4434 18864
rect 4490 18808 11058 18864
rect 11114 18808 11119 18864
rect 4429 18806 11119 18808
rect 4429 18803 4495 18806
rect 11053 18803 11119 18806
rect 11286 18806 14106 18866
rect 15009 18866 15075 18869
rect 26233 18866 26299 18869
rect 15009 18864 26299 18866
rect 15009 18808 15014 18864
rect 15070 18808 26238 18864
rect 26294 18808 26299 18864
rect 15009 18806 26299 18808
rect 0 18730 800 18760
rect 3325 18730 3391 18733
rect 0 18728 3391 18730
rect 0 18672 3330 18728
rect 3386 18672 3391 18728
rect 0 18670 3391 18672
rect 0 18640 800 18670
rect 3325 18667 3391 18670
rect 3550 18668 3556 18732
rect 3620 18730 3626 18732
rect 11286 18730 11346 18806
rect 15009 18803 15075 18806
rect 26233 18803 26299 18806
rect 26509 18866 26575 18869
rect 45737 18866 45803 18869
rect 26509 18864 45803 18866
rect 26509 18808 26514 18864
rect 26570 18808 45742 18864
rect 45798 18808 45803 18864
rect 26509 18806 45803 18808
rect 26509 18803 26575 18806
rect 45737 18803 45803 18806
rect 3620 18670 11346 18730
rect 11513 18730 11579 18733
rect 14457 18730 14523 18733
rect 19241 18730 19307 18733
rect 11513 18728 14523 18730
rect 11513 18672 11518 18728
rect 11574 18672 14462 18728
rect 14518 18672 14523 18728
rect 11513 18670 14523 18672
rect 3620 18668 3626 18670
rect 11513 18667 11579 18670
rect 14457 18667 14523 18670
rect 17174 18728 19307 18730
rect 17174 18672 19246 18728
rect 19302 18672 19307 18728
rect 17174 18670 19307 18672
rect 10501 18594 10567 18597
rect 13169 18594 13235 18597
rect 10501 18592 13235 18594
rect 10501 18536 10506 18592
rect 10562 18536 13174 18592
rect 13230 18536 13235 18592
rect 10501 18534 13235 18536
rect 10501 18531 10567 18534
rect 13169 18531 13235 18534
rect 13629 18594 13695 18597
rect 17033 18594 17099 18597
rect 13629 18592 17099 18594
rect 13629 18536 13634 18592
rect 13690 18536 17038 18592
rect 17094 18536 17099 18592
rect 13629 18534 17099 18536
rect 13629 18531 13695 18534
rect 17033 18531 17099 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 6085 18460 6151 18461
rect 6085 18458 6132 18460
rect 5950 18456 6132 18458
rect 6196 18458 6202 18460
rect 9857 18458 9923 18461
rect 10409 18458 10475 18461
rect 15193 18458 15259 18461
rect 17174 18458 17234 18670
rect 19241 18667 19307 18670
rect 19517 18730 19583 18733
rect 23381 18730 23447 18733
rect 19517 18728 23447 18730
rect 19517 18672 19522 18728
rect 19578 18672 23386 18728
rect 23442 18672 23447 18728
rect 19517 18670 23447 18672
rect 19517 18667 19583 18670
rect 23381 18667 23447 18670
rect 25405 18730 25471 18733
rect 45369 18730 45435 18733
rect 25405 18728 45435 18730
rect 25405 18672 25410 18728
rect 25466 18672 45374 18728
rect 45430 18672 45435 18728
rect 25405 18670 45435 18672
rect 25405 18667 25471 18670
rect 45369 18667 45435 18670
rect 18873 18594 18939 18597
rect 24393 18594 24459 18597
rect 18873 18592 24459 18594
rect 18873 18536 18878 18592
rect 18934 18536 24398 18592
rect 24454 18536 24459 18592
rect 18873 18534 24459 18536
rect 18873 18531 18939 18534
rect 24393 18531 24459 18534
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 47946 18463 48262 18464
rect 5950 18400 6090 18456
rect 5950 18398 6132 18400
rect 0 18322 800 18352
rect 2865 18322 2931 18325
rect 0 18320 2931 18322
rect 0 18264 2870 18320
rect 2926 18264 2931 18320
rect 0 18262 2931 18264
rect 0 18232 800 18262
rect 2865 18259 2931 18262
rect 5625 18322 5691 18325
rect 5950 18322 6010 18398
rect 6085 18396 6132 18398
rect 6196 18398 6278 18458
rect 9857 18456 15259 18458
rect 9857 18400 9862 18456
rect 9918 18400 10414 18456
rect 10470 18400 15198 18456
rect 15254 18400 15259 18456
rect 9857 18398 15259 18400
rect 6196 18396 6202 18398
rect 6085 18395 6151 18396
rect 9857 18395 9923 18398
rect 10409 18395 10475 18398
rect 15193 18395 15259 18398
rect 15334 18398 17234 18458
rect 19425 18458 19491 18461
rect 22001 18458 22067 18461
rect 19425 18456 22067 18458
rect 19425 18400 19430 18456
rect 19486 18400 22006 18456
rect 22062 18400 22067 18456
rect 19425 18398 22067 18400
rect 5625 18320 6010 18322
rect 5625 18264 5630 18320
rect 5686 18264 6010 18320
rect 5625 18262 6010 18264
rect 6729 18322 6795 18325
rect 15334 18322 15394 18398
rect 19425 18395 19491 18398
rect 22001 18395 22067 18398
rect 22921 18458 22987 18461
rect 27245 18458 27311 18461
rect 22921 18456 27311 18458
rect 22921 18400 22926 18456
rect 22982 18400 27250 18456
rect 27306 18400 27311 18456
rect 22921 18398 27311 18400
rect 22921 18395 22987 18398
rect 27245 18395 27311 18398
rect 6729 18320 15394 18322
rect 6729 18264 6734 18320
rect 6790 18264 15394 18320
rect 6729 18262 15394 18264
rect 16389 18322 16455 18325
rect 17585 18322 17651 18325
rect 16389 18320 17651 18322
rect 16389 18264 16394 18320
rect 16450 18264 17590 18320
rect 17646 18264 17651 18320
rect 16389 18262 17651 18264
rect 5625 18259 5691 18262
rect 6729 18259 6795 18262
rect 16389 18259 16455 18262
rect 17585 18259 17651 18262
rect 18321 18322 18387 18325
rect 31201 18322 31267 18325
rect 18321 18320 31267 18322
rect 18321 18264 18326 18320
rect 18382 18264 31206 18320
rect 31262 18264 31267 18320
rect 18321 18262 31267 18264
rect 18321 18259 18387 18262
rect 31201 18259 31267 18262
rect 5901 18186 5967 18189
rect 6453 18186 6519 18189
rect 9305 18186 9371 18189
rect 32673 18186 32739 18189
rect 5901 18184 9371 18186
rect 5901 18128 5906 18184
rect 5962 18128 6458 18184
rect 6514 18128 9310 18184
rect 9366 18128 9371 18184
rect 5901 18126 9371 18128
rect 5901 18123 5967 18126
rect 6453 18123 6519 18126
rect 9305 18123 9371 18126
rect 12390 18184 32739 18186
rect 12390 18128 32678 18184
rect 32734 18128 32739 18184
rect 12390 18126 32739 18128
rect 3366 17988 3372 18052
rect 3436 18050 3442 18052
rect 3969 18050 4035 18053
rect 3436 18048 4035 18050
rect 3436 17992 3974 18048
rect 4030 17992 4035 18048
rect 3436 17990 4035 17992
rect 3436 17988 3442 17990
rect 3969 17987 4035 17990
rect 11881 18050 11947 18053
rect 12390 18050 12450 18126
rect 32673 18123 32739 18126
rect 11881 18048 12450 18050
rect 11881 17992 11886 18048
rect 11942 17992 12450 18048
rect 11881 17990 12450 17992
rect 14733 18050 14799 18053
rect 16849 18050 16915 18053
rect 21081 18050 21147 18053
rect 22461 18050 22527 18053
rect 14733 18048 16915 18050
rect 14733 17992 14738 18048
rect 14794 17992 16854 18048
rect 16910 17992 16915 18048
rect 14733 17990 16915 17992
rect 11881 17987 11947 17990
rect 14733 17987 14799 17990
rect 16849 17987 16915 17990
rect 19290 18048 22527 18050
rect 19290 17992 21086 18048
rect 21142 17992 22466 18048
rect 22522 17992 22527 18048
rect 19290 17990 22527 17992
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 2773 17914 2839 17917
rect 0 17912 2839 17914
rect 0 17856 2778 17912
rect 2834 17856 2839 17912
rect 0 17854 2839 17856
rect 0 17824 800 17854
rect 2773 17851 2839 17854
rect 4797 17914 4863 17917
rect 7281 17914 7347 17917
rect 8017 17914 8083 17917
rect 4797 17912 8083 17914
rect 4797 17856 4802 17912
rect 4858 17856 7286 17912
rect 7342 17856 8022 17912
rect 8078 17856 8083 17912
rect 4797 17854 8083 17856
rect 4797 17851 4863 17854
rect 7281 17851 7347 17854
rect 8017 17851 8083 17854
rect 10133 17914 10199 17917
rect 10593 17914 10659 17917
rect 10133 17912 10659 17914
rect 10133 17856 10138 17912
rect 10194 17856 10598 17912
rect 10654 17856 10659 17912
rect 10133 17854 10659 17856
rect 10133 17851 10199 17854
rect 10593 17851 10659 17854
rect 17125 17914 17191 17917
rect 18873 17914 18939 17917
rect 17125 17912 18939 17914
rect 17125 17856 17130 17912
rect 17186 17856 18878 17912
rect 18934 17856 18939 17912
rect 17125 17854 18939 17856
rect 17125 17851 17191 17854
rect 18873 17851 18939 17854
rect 2221 17778 2287 17781
rect 3785 17778 3851 17781
rect 9581 17778 9647 17781
rect 2221 17776 9647 17778
rect 2221 17720 2226 17776
rect 2282 17720 3790 17776
rect 3846 17720 9586 17776
rect 9642 17720 9647 17776
rect 2221 17718 9647 17720
rect 2221 17715 2287 17718
rect 3785 17715 3851 17718
rect 9581 17715 9647 17718
rect 11881 17778 11947 17781
rect 13261 17778 13327 17781
rect 11881 17776 13327 17778
rect 11881 17720 11886 17776
rect 11942 17720 13266 17776
rect 13322 17720 13327 17776
rect 11881 17718 13327 17720
rect 11881 17715 11947 17718
rect 13261 17715 13327 17718
rect 17769 17778 17835 17781
rect 19290 17778 19350 17990
rect 21081 17987 21147 17990
rect 22461 17987 22527 17990
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 23749 17914 23815 17917
rect 30649 17914 30715 17917
rect 23749 17912 30715 17914
rect 23749 17856 23754 17912
rect 23810 17856 30654 17912
rect 30710 17856 30715 17912
rect 23749 17854 30715 17856
rect 23749 17851 23815 17854
rect 30649 17851 30715 17854
rect 17769 17776 19350 17778
rect 17769 17720 17774 17776
rect 17830 17720 19350 17776
rect 17769 17718 19350 17720
rect 17769 17715 17835 17718
rect 4061 17642 4127 17645
rect 7189 17642 7255 17645
rect 11513 17642 11579 17645
rect 14457 17642 14523 17645
rect 20529 17642 20595 17645
rect 4061 17640 11579 17642
rect 4061 17584 4066 17640
rect 4122 17584 7194 17640
rect 7250 17584 11518 17640
rect 11574 17584 11579 17640
rect 4061 17582 11579 17584
rect 4061 17579 4127 17582
rect 7189 17579 7255 17582
rect 11513 17579 11579 17582
rect 12390 17640 14523 17642
rect 12390 17584 14462 17640
rect 14518 17584 14523 17640
rect 12390 17582 14523 17584
rect 0 17506 800 17536
rect 2037 17506 2103 17509
rect 0 17504 2103 17506
rect 0 17448 2042 17504
rect 2098 17448 2103 17504
rect 0 17446 2103 17448
rect 0 17416 800 17446
rect 2037 17443 2103 17446
rect 5942 17444 5948 17508
rect 6012 17506 6018 17508
rect 6177 17506 6243 17509
rect 6012 17504 6243 17506
rect 6012 17448 6182 17504
rect 6238 17448 6243 17504
rect 6012 17446 6243 17448
rect 6012 17444 6018 17446
rect 6177 17443 6243 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 12390 17370 12450 17582
rect 14457 17579 14523 17582
rect 14598 17640 20595 17642
rect 14598 17584 20534 17640
rect 20590 17584 20595 17640
rect 14598 17582 20595 17584
rect 12525 17506 12591 17509
rect 14598 17506 14658 17582
rect 20529 17579 20595 17582
rect 21357 17642 21423 17645
rect 31937 17642 32003 17645
rect 21357 17640 32003 17642
rect 21357 17584 21362 17640
rect 21418 17584 31942 17640
rect 31998 17584 32003 17640
rect 21357 17582 32003 17584
rect 21357 17579 21423 17582
rect 31937 17579 32003 17582
rect 12525 17504 14658 17506
rect 12525 17448 12530 17504
rect 12586 17448 14658 17504
rect 12525 17446 14658 17448
rect 12525 17443 12591 17446
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 8342 17310 12450 17370
rect 4429 17234 4495 17237
rect 8342 17234 8402 17310
rect 18454 17234 18460 17236
rect 4429 17232 8402 17234
rect 4429 17176 4434 17232
rect 4490 17176 8402 17232
rect 4429 17174 8402 17176
rect 8710 17174 18460 17234
rect 4429 17171 4495 17174
rect 0 17098 800 17128
rect 1209 17098 1275 17101
rect 0 17096 1275 17098
rect 0 17040 1214 17096
rect 1270 17040 1275 17096
rect 0 17038 1275 17040
rect 0 17008 800 17038
rect 1209 17035 1275 17038
rect 4061 17098 4127 17101
rect 8569 17098 8635 17101
rect 8710 17098 8770 17174
rect 18454 17172 18460 17174
rect 18524 17172 18530 17236
rect 19609 17234 19675 17237
rect 23933 17234 23999 17237
rect 19609 17232 23999 17234
rect 19609 17176 19614 17232
rect 19670 17176 23938 17232
rect 23994 17176 23999 17232
rect 19609 17174 23999 17176
rect 19609 17171 19675 17174
rect 23933 17171 23999 17174
rect 25957 17234 26023 17237
rect 46841 17234 46907 17237
rect 25957 17232 46907 17234
rect 25957 17176 25962 17232
rect 26018 17176 46846 17232
rect 46902 17176 46907 17232
rect 25957 17174 46907 17176
rect 25957 17171 26023 17174
rect 46841 17171 46907 17174
rect 4061 17096 8770 17098
rect 4061 17040 4066 17096
rect 4122 17040 8574 17096
rect 8630 17040 8770 17096
rect 4061 17038 8770 17040
rect 8937 17098 9003 17101
rect 18321 17098 18387 17101
rect 8937 17096 18387 17098
rect 8937 17040 8942 17096
rect 8998 17040 18326 17096
rect 18382 17040 18387 17096
rect 8937 17038 18387 17040
rect 4061 17035 4127 17038
rect 8569 17035 8635 17038
rect 8937 17035 9003 17038
rect 18321 17035 18387 17038
rect 11513 16962 11579 16965
rect 12525 16962 12591 16965
rect 11513 16960 12591 16962
rect 11513 16904 11518 16960
rect 11574 16904 12530 16960
rect 12586 16904 12591 16960
rect 11513 16902 12591 16904
rect 11513 16899 11579 16902
rect 12525 16899 12591 16902
rect 13721 16962 13787 16965
rect 20069 16962 20135 16965
rect 13721 16960 20135 16962
rect 13721 16904 13726 16960
rect 13782 16904 20074 16960
rect 20130 16904 20135 16960
rect 13721 16902 20135 16904
rect 13721 16899 13787 16902
rect 20069 16899 20135 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 3509 16826 3575 16829
rect 8109 16826 8175 16829
rect 12801 16826 12867 16829
rect 3509 16824 12867 16826
rect 3509 16768 3514 16824
rect 3570 16768 8114 16824
rect 8170 16768 12806 16824
rect 12862 16768 12867 16824
rect 3509 16766 12867 16768
rect 3509 16763 3575 16766
rect 8109 16763 8175 16766
rect 12801 16763 12867 16766
rect 13353 16826 13419 16829
rect 16941 16826 17007 16829
rect 20161 16826 20227 16829
rect 13353 16824 16866 16826
rect 13353 16768 13358 16824
rect 13414 16768 16866 16824
rect 13353 16766 16866 16768
rect 13353 16763 13419 16766
rect 0 16690 800 16720
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 800 16630
rect 1301 16627 1367 16630
rect 5625 16690 5691 16693
rect 5758 16690 5764 16692
rect 5625 16688 5764 16690
rect 5625 16632 5630 16688
rect 5686 16632 5764 16688
rect 5625 16630 5764 16632
rect 5625 16627 5691 16630
rect 5758 16628 5764 16630
rect 5828 16628 5834 16692
rect 8385 16690 8451 16693
rect 8518 16690 8524 16692
rect 8385 16688 8524 16690
rect 8385 16632 8390 16688
rect 8446 16632 8524 16688
rect 8385 16630 8524 16632
rect 8385 16627 8451 16630
rect 8518 16628 8524 16630
rect 8588 16628 8594 16692
rect 8845 16690 8911 16693
rect 11789 16690 11855 16693
rect 8845 16688 11855 16690
rect 8845 16632 8850 16688
rect 8906 16632 11794 16688
rect 11850 16632 11855 16688
rect 8845 16630 11855 16632
rect 8845 16627 8911 16630
rect 11789 16627 11855 16630
rect 12985 16690 13051 16693
rect 16573 16690 16639 16693
rect 12985 16688 16639 16690
rect 12985 16632 12990 16688
rect 13046 16632 16578 16688
rect 16634 16632 16639 16688
rect 12985 16630 16639 16632
rect 16806 16690 16866 16766
rect 16941 16824 20227 16826
rect 16941 16768 16946 16824
rect 17002 16768 20166 16824
rect 20222 16768 20227 16824
rect 16941 16766 20227 16768
rect 16941 16763 17007 16766
rect 20161 16763 20227 16766
rect 17769 16690 17835 16693
rect 16806 16688 17835 16690
rect 16806 16632 17774 16688
rect 17830 16632 17835 16688
rect 16806 16630 17835 16632
rect 12985 16627 13051 16630
rect 16573 16627 16639 16630
rect 17769 16627 17835 16630
rect 18597 16690 18663 16693
rect 18965 16690 19031 16693
rect 21265 16690 21331 16693
rect 18597 16688 21331 16690
rect 18597 16632 18602 16688
rect 18658 16632 18970 16688
rect 19026 16632 21270 16688
rect 21326 16632 21331 16688
rect 18597 16630 21331 16632
rect 18597 16627 18663 16630
rect 18965 16627 19031 16630
rect 21265 16627 21331 16630
rect 25681 16690 25747 16693
rect 26509 16690 26575 16693
rect 25681 16688 26575 16690
rect 25681 16632 25686 16688
rect 25742 16632 26514 16688
rect 26570 16632 26575 16688
rect 25681 16630 26575 16632
rect 25681 16627 25747 16630
rect 26509 16627 26575 16630
rect 6453 16554 6519 16557
rect 8201 16554 8267 16557
rect 6453 16552 8267 16554
rect 6453 16496 6458 16552
rect 6514 16496 8206 16552
rect 8262 16496 8267 16552
rect 6453 16494 8267 16496
rect 6453 16491 6519 16494
rect 8201 16491 8267 16494
rect 8334 16492 8340 16556
rect 8404 16554 8410 16556
rect 9857 16554 9923 16557
rect 8404 16552 9923 16554
rect 8404 16496 9862 16552
rect 9918 16496 9923 16552
rect 8404 16494 9923 16496
rect 8404 16492 8410 16494
rect 9857 16491 9923 16494
rect 14365 16554 14431 16557
rect 28533 16554 28599 16557
rect 14365 16552 28599 16554
rect 14365 16496 14370 16552
rect 14426 16496 28538 16552
rect 28594 16496 28599 16552
rect 14365 16494 28599 16496
rect 14365 16491 14431 16494
rect 28533 16491 28599 16494
rect 16941 16420 17007 16421
rect 17493 16420 17559 16421
rect 16941 16418 16988 16420
rect 16896 16416 16988 16418
rect 16896 16360 16946 16416
rect 16896 16358 16988 16360
rect 16941 16356 16988 16358
rect 17052 16356 17058 16420
rect 17493 16416 17540 16420
rect 17604 16418 17610 16420
rect 21449 16418 21515 16421
rect 24117 16418 24183 16421
rect 17493 16360 17498 16416
rect 17493 16356 17540 16360
rect 17604 16358 17650 16418
rect 21449 16416 24183 16418
rect 21449 16360 21454 16416
rect 21510 16360 24122 16416
rect 24178 16360 24183 16416
rect 21449 16358 24183 16360
rect 17604 16356 17610 16358
rect 16941 16355 17007 16356
rect 17493 16355 17559 16356
rect 21449 16355 21515 16358
rect 24117 16355 24183 16358
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 9622 16220 9628 16284
rect 9692 16282 9698 16284
rect 10593 16282 10659 16285
rect 17125 16284 17191 16285
rect 17125 16282 17172 16284
rect 9692 16280 10659 16282
rect 9692 16224 10598 16280
rect 10654 16224 10659 16280
rect 9692 16222 10659 16224
rect 17080 16280 17172 16282
rect 17080 16224 17130 16280
rect 17080 16222 17172 16224
rect 9692 16220 9698 16222
rect 10593 16219 10659 16222
rect 17125 16220 17172 16222
rect 17236 16220 17242 16284
rect 17125 16219 17191 16220
rect 7373 16146 7439 16149
rect 7925 16146 7991 16149
rect 10961 16146 11027 16149
rect 19333 16146 19399 16149
rect 7373 16144 7991 16146
rect 7373 16088 7378 16144
rect 7434 16088 7930 16144
rect 7986 16088 7991 16144
rect 7373 16086 7991 16088
rect 7373 16083 7439 16086
rect 7925 16083 7991 16086
rect 9630 16144 19399 16146
rect 9630 16088 10966 16144
rect 11022 16088 19338 16144
rect 19394 16088 19399 16144
rect 9630 16086 19399 16088
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 4889 15738 4955 15741
rect 9630 15738 9690 16086
rect 10961 16083 11027 16086
rect 19333 16083 19399 16086
rect 10961 16010 11027 16013
rect 29545 16010 29611 16013
rect 10961 16008 29611 16010
rect 10961 15952 10966 16008
rect 11022 15952 29550 16008
rect 29606 15952 29611 16008
rect 10961 15950 29611 15952
rect 10961 15947 11027 15950
rect 29545 15947 29611 15950
rect 9806 15812 9812 15876
rect 9876 15874 9882 15876
rect 10542 15874 10548 15876
rect 9876 15814 10548 15874
rect 9876 15812 9882 15814
rect 10542 15812 10548 15814
rect 10612 15874 10618 15876
rect 10685 15874 10751 15877
rect 10612 15872 10751 15874
rect 10612 15816 10690 15872
rect 10746 15816 10751 15872
rect 10612 15814 10751 15816
rect 10612 15812 10618 15814
rect 10685 15811 10751 15814
rect 15377 15874 15443 15877
rect 16573 15874 16639 15877
rect 15377 15872 16639 15874
rect 15377 15816 15382 15872
rect 15438 15816 16578 15872
rect 16634 15816 16639 15872
rect 15377 15814 16639 15816
rect 15377 15811 15443 15814
rect 16573 15811 16639 15814
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 4889 15736 9690 15738
rect 4889 15680 4894 15736
rect 4950 15680 9690 15736
rect 4889 15678 9690 15680
rect 13353 15738 13419 15741
rect 22277 15738 22343 15741
rect 13353 15736 22343 15738
rect 13353 15680 13358 15736
rect 13414 15680 22282 15736
rect 22338 15680 22343 15736
rect 13353 15678 22343 15680
rect 4889 15675 4955 15678
rect 3918 15540 3924 15604
rect 3988 15602 3994 15604
rect 3988 15542 6746 15602
rect 3988 15540 3994 15542
rect 0 15466 800 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 800 15406
rect 1301 15403 1367 15406
rect 3918 15404 3924 15468
rect 3988 15466 3994 15468
rect 6453 15466 6519 15469
rect 3988 15464 6519 15466
rect 3988 15408 6458 15464
rect 6514 15408 6519 15464
rect 3988 15406 6519 15408
rect 6686 15466 6746 15542
rect 8664 15469 8724 15678
rect 13353 15675 13419 15678
rect 22277 15675 22343 15678
rect 9213 15602 9279 15605
rect 21357 15602 21423 15605
rect 9213 15600 21423 15602
rect 9213 15544 9218 15600
rect 9274 15544 21362 15600
rect 21418 15544 21423 15600
rect 9213 15542 21423 15544
rect 9213 15539 9279 15542
rect 21357 15539 21423 15542
rect 22093 15602 22159 15605
rect 22921 15602 22987 15605
rect 22093 15600 22987 15602
rect 22093 15544 22098 15600
rect 22154 15544 22926 15600
rect 22982 15544 22987 15600
rect 22093 15542 22987 15544
rect 22093 15539 22159 15542
rect 22921 15539 22987 15542
rect 8477 15466 8543 15469
rect 6686 15464 8543 15466
rect 6686 15408 8482 15464
rect 8538 15408 8543 15464
rect 6686 15406 8543 15408
rect 3988 15404 3994 15406
rect 6453 15403 6519 15406
rect 8477 15403 8543 15406
rect 8661 15464 8727 15469
rect 8661 15408 8666 15464
rect 8722 15408 8727 15464
rect 8661 15403 8727 15408
rect 12065 15466 12131 15469
rect 29913 15466 29979 15469
rect 12065 15464 29979 15466
rect 12065 15408 12070 15464
rect 12126 15408 29918 15464
rect 29974 15408 29979 15464
rect 12065 15406 29979 15408
rect 12065 15403 12131 15406
rect 29913 15403 29979 15406
rect 3785 15330 3851 15333
rect 7373 15330 7439 15333
rect 3785 15328 7439 15330
rect 3785 15272 3790 15328
rect 3846 15272 7378 15328
rect 7434 15272 7439 15328
rect 3785 15270 7439 15272
rect 3785 15267 3851 15270
rect 7373 15267 7439 15270
rect 10777 15330 10843 15333
rect 17493 15330 17559 15333
rect 10777 15328 17559 15330
rect 10777 15272 10782 15328
rect 10838 15272 17498 15328
rect 17554 15272 17559 15328
rect 10777 15270 17559 15272
rect 10777 15267 10843 15270
rect 17493 15267 17559 15270
rect 19517 15330 19583 15333
rect 25589 15330 25655 15333
rect 19517 15328 25655 15330
rect 19517 15272 19522 15328
rect 19578 15272 25594 15328
rect 25650 15272 25655 15328
rect 19517 15270 25655 15272
rect 19517 15267 19583 15270
rect 25589 15267 25655 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 12249 15194 12315 15197
rect 13261 15194 13327 15197
rect 12249 15192 13327 15194
rect 12249 15136 12254 15192
rect 12310 15136 13266 15192
rect 13322 15136 13327 15192
rect 12249 15134 13327 15136
rect 12249 15131 12315 15134
rect 13261 15131 13327 15134
rect 0 15058 800 15088
rect 1301 15058 1367 15061
rect 0 15056 1367 15058
rect 0 15000 1306 15056
rect 1362 15000 1367 15056
rect 0 14998 1367 15000
rect 0 14968 800 14998
rect 1301 14995 1367 14998
rect 5717 15058 5783 15061
rect 8569 15058 8635 15061
rect 5717 15056 8635 15058
rect 5717 15000 5722 15056
rect 5778 15000 8574 15056
rect 8630 15000 8635 15056
rect 5717 14998 8635 15000
rect 5717 14995 5783 14998
rect 8569 14995 8635 14998
rect 11973 15058 12039 15061
rect 33317 15058 33383 15061
rect 11973 15056 33383 15058
rect 11973 15000 11978 15056
rect 12034 15000 33322 15056
rect 33378 15000 33383 15056
rect 11973 14998 33383 15000
rect 11973 14995 12039 14998
rect 33317 14995 33383 14998
rect 7833 14922 7899 14925
rect 8845 14922 8911 14925
rect 7833 14920 8911 14922
rect 7833 14864 7838 14920
rect 7894 14864 8850 14920
rect 8906 14864 8911 14920
rect 7833 14862 8911 14864
rect 7833 14859 7899 14862
rect 8845 14859 8911 14862
rect 17125 14922 17191 14925
rect 19333 14922 19399 14925
rect 17125 14920 19399 14922
rect 17125 14864 17130 14920
rect 17186 14864 19338 14920
rect 19394 14864 19399 14920
rect 17125 14862 19399 14864
rect 17125 14859 17191 14862
rect 19333 14859 19399 14862
rect 9765 14786 9831 14789
rect 10317 14786 10383 14789
rect 9765 14784 10383 14786
rect 9765 14728 9770 14784
rect 9826 14728 10322 14784
rect 10378 14728 10383 14784
rect 9765 14726 10383 14728
rect 9765 14723 9831 14726
rect 10317 14723 10383 14726
rect 15561 14786 15627 14789
rect 18781 14786 18847 14789
rect 15561 14784 18847 14786
rect 15561 14728 15566 14784
rect 15622 14728 18786 14784
rect 18842 14728 18847 14784
rect 15561 14726 18847 14728
rect 15561 14723 15627 14726
rect 18781 14723 18847 14726
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 1301 14650 1367 14653
rect 0 14648 1367 14650
rect 0 14592 1306 14648
rect 1362 14592 1367 14648
rect 0 14590 1367 14592
rect 0 14560 800 14590
rect 1301 14587 1367 14590
rect 6453 14514 6519 14517
rect 11881 14514 11947 14517
rect 6453 14512 12450 14514
rect 6453 14456 6458 14512
rect 6514 14456 11886 14512
rect 11942 14456 12450 14512
rect 6453 14454 12450 14456
rect 6453 14451 6519 14454
rect 11881 14451 11947 14454
rect 6453 14378 6519 14381
rect 8477 14378 8543 14381
rect 6453 14376 8543 14378
rect 6453 14320 6458 14376
rect 6514 14320 8482 14376
rect 8538 14320 8543 14376
rect 6453 14318 8543 14320
rect 12390 14378 12450 14454
rect 12893 14378 12959 14381
rect 12390 14376 12959 14378
rect 12390 14320 12898 14376
rect 12954 14320 12959 14376
rect 12390 14318 12959 14320
rect 6453 14315 6519 14318
rect 8477 14315 8543 14318
rect 12893 14315 12959 14318
rect 15837 14378 15903 14381
rect 16205 14378 16271 14381
rect 20713 14378 20779 14381
rect 15837 14376 20779 14378
rect 15837 14320 15842 14376
rect 15898 14320 16210 14376
rect 16266 14320 20718 14376
rect 20774 14320 20779 14376
rect 15837 14318 20779 14320
rect 15837 14315 15903 14318
rect 16205 14315 16271 14318
rect 20713 14315 20779 14318
rect 0 14242 800 14272
rect 1301 14242 1367 14245
rect 0 14240 1367 14242
rect 0 14184 1306 14240
rect 1362 14184 1367 14240
rect 0 14182 1367 14184
rect 0 14152 800 14182
rect 1301 14179 1367 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 4797 14106 4863 14109
rect 6545 14106 6611 14109
rect 4797 14104 6611 14106
rect 4797 14048 4802 14104
rect 4858 14048 6550 14104
rect 6606 14048 6611 14104
rect 4797 14046 6611 14048
rect 4797 14043 4863 14046
rect 6545 14043 6611 14046
rect 1761 13970 1827 13973
rect 19885 13970 19951 13973
rect 1761 13968 19951 13970
rect 1761 13912 1766 13968
rect 1822 13912 19890 13968
rect 19946 13912 19951 13968
rect 1761 13910 19951 13912
rect 1761 13907 1827 13910
rect 19885 13907 19951 13910
rect 0 13834 800 13864
rect 2037 13834 2103 13837
rect 0 13832 2103 13834
rect 0 13776 2042 13832
rect 2098 13776 2103 13832
rect 0 13774 2103 13776
rect 0 13744 800 13774
rect 2037 13771 2103 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 0 13426 800 13456
rect 1209 13426 1275 13429
rect 0 13424 1275 13426
rect 0 13368 1214 13424
rect 1270 13368 1275 13424
rect 0 13366 1275 13368
rect 0 13336 800 13366
rect 1209 13363 1275 13366
rect 9397 13426 9463 13429
rect 30741 13426 30807 13429
rect 9397 13424 30807 13426
rect 9397 13368 9402 13424
rect 9458 13368 30746 13424
rect 30802 13368 30807 13424
rect 9397 13366 30807 13368
rect 9397 13363 9463 13366
rect 30741 13363 30807 13366
rect 1761 13290 1827 13293
rect 22001 13290 22067 13293
rect 1761 13288 22067 13290
rect 1761 13232 1766 13288
rect 1822 13232 22006 13288
rect 22062 13232 22067 13288
rect 1761 13230 22067 13232
rect 1761 13227 1827 13230
rect 22001 13227 22067 13230
rect 23105 13290 23171 13293
rect 25221 13290 25287 13293
rect 23105 13288 25287 13290
rect 23105 13232 23110 13288
rect 23166 13232 25226 13288
rect 25282 13232 25287 13288
rect 23105 13230 25287 13232
rect 23105 13227 23171 13230
rect 25221 13227 25287 13230
rect 4705 13154 4771 13157
rect 6126 13154 6132 13156
rect 4705 13152 6132 13154
rect 4705 13096 4710 13152
rect 4766 13096 6132 13152
rect 4705 13094 6132 13096
rect 4705 13091 4771 13094
rect 6126 13092 6132 13094
rect 6196 13092 6202 13156
rect 13997 13154 14063 13157
rect 15285 13154 15351 13157
rect 13997 13152 15351 13154
rect 13997 13096 14002 13152
rect 14058 13096 15290 13152
rect 15346 13096 15351 13152
rect 13997 13094 15351 13096
rect 13997 13091 14063 13094
rect 15285 13091 15351 13094
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 3417 13018 3483 13021
rect 0 13016 3483 13018
rect 0 12960 3422 13016
rect 3478 12960 3483 13016
rect 0 12958 3483 12960
rect 0 12928 800 12958
rect 3417 12955 3483 12958
rect 10685 12882 10751 12885
rect 21081 12882 21147 12885
rect 10685 12880 21147 12882
rect 10685 12824 10690 12880
rect 10746 12824 21086 12880
rect 21142 12824 21147 12880
rect 10685 12822 21147 12824
rect 10685 12819 10751 12822
rect 21081 12819 21147 12822
rect 7281 12746 7347 12749
rect 12433 12746 12499 12749
rect 7281 12744 12499 12746
rect 7281 12688 7286 12744
rect 7342 12688 12438 12744
rect 12494 12688 12499 12744
rect 7281 12686 12499 12688
rect 7281 12683 7347 12686
rect 12433 12683 12499 12686
rect 18454 12684 18460 12748
rect 18524 12746 18530 12748
rect 18597 12746 18663 12749
rect 18524 12744 18663 12746
rect 18524 12688 18602 12744
rect 18658 12688 18663 12744
rect 18524 12686 18663 12688
rect 18524 12684 18530 12686
rect 18597 12683 18663 12686
rect 0 12610 800 12640
rect 2037 12610 2103 12613
rect 0 12608 2103 12610
rect 0 12552 2042 12608
rect 2098 12552 2103 12608
rect 0 12550 2103 12552
rect 0 12520 800 12550
rect 2037 12547 2103 12550
rect 10317 12610 10383 12613
rect 10961 12610 11027 12613
rect 10317 12608 11027 12610
rect 10317 12552 10322 12608
rect 10378 12552 10966 12608
rect 11022 12552 11027 12608
rect 10317 12550 11027 12552
rect 10317 12547 10383 12550
rect 10961 12547 11027 12550
rect 15193 12610 15259 12613
rect 19149 12610 19215 12613
rect 15193 12608 19215 12610
rect 15193 12552 15198 12608
rect 15254 12552 19154 12608
rect 19210 12552 19215 12608
rect 15193 12550 19215 12552
rect 15193 12547 15259 12550
rect 19149 12547 19215 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 7557 12474 7623 12477
rect 11094 12474 11100 12476
rect 7557 12472 11100 12474
rect 7557 12416 7562 12472
rect 7618 12416 11100 12472
rect 7557 12414 11100 12416
rect 7557 12411 7623 12414
rect 11094 12412 11100 12414
rect 11164 12412 11170 12476
rect 2957 12338 3023 12341
rect 3325 12338 3391 12341
rect 4245 12340 4311 12341
rect 7373 12340 7439 12341
rect 3918 12338 3924 12340
rect 2957 12336 3924 12338
rect 2957 12280 2962 12336
rect 3018 12280 3330 12336
rect 3386 12280 3924 12336
rect 2957 12278 3924 12280
rect 2957 12275 3023 12278
rect 3325 12275 3391 12278
rect 3918 12276 3924 12278
rect 3988 12276 3994 12340
rect 4245 12338 4292 12340
rect 4200 12336 4292 12338
rect 4200 12280 4250 12336
rect 4200 12278 4292 12280
rect 4245 12276 4292 12278
rect 4356 12276 4362 12340
rect 7373 12338 7420 12340
rect 7328 12336 7420 12338
rect 7328 12280 7378 12336
rect 7328 12278 7420 12280
rect 7373 12276 7420 12278
rect 7484 12276 7490 12340
rect 19609 12338 19675 12341
rect 25037 12338 25103 12341
rect 19609 12336 25103 12338
rect 19609 12280 19614 12336
rect 19670 12280 25042 12336
rect 25098 12280 25103 12336
rect 19609 12278 25103 12280
rect 4245 12275 4311 12276
rect 7373 12275 7439 12276
rect 19609 12275 19675 12278
rect 25037 12275 25103 12278
rect 0 12202 800 12232
rect 1301 12202 1367 12205
rect 0 12200 1367 12202
rect 0 12144 1306 12200
rect 1362 12144 1367 12200
rect 0 12142 1367 12144
rect 0 12112 800 12142
rect 1301 12139 1367 12142
rect 3601 12202 3667 12205
rect 9806 12202 9812 12204
rect 3601 12200 9812 12202
rect 3601 12144 3606 12200
rect 3662 12144 9812 12200
rect 3601 12142 9812 12144
rect 3601 12139 3667 12142
rect 9806 12140 9812 12142
rect 9876 12140 9882 12204
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 6177 11930 6243 11933
rect 7046 11930 7052 11932
rect 6177 11928 7052 11930
rect 6177 11872 6182 11928
rect 6238 11872 7052 11928
rect 6177 11870 7052 11872
rect 6177 11867 6243 11870
rect 7046 11868 7052 11870
rect 7116 11868 7122 11932
rect 12249 11930 12315 11933
rect 17309 11930 17375 11933
rect 12249 11928 17375 11930
rect 12249 11872 12254 11928
rect 12310 11872 17314 11928
rect 17370 11872 17375 11928
rect 12249 11870 17375 11872
rect 12249 11867 12315 11870
rect 17309 11867 17375 11870
rect 0 11794 800 11824
rect 1393 11794 1459 11797
rect 0 11792 1459 11794
rect 0 11736 1398 11792
rect 1454 11736 1459 11792
rect 0 11734 1459 11736
rect 0 11704 800 11734
rect 1393 11731 1459 11734
rect 12433 11794 12499 11797
rect 13077 11794 13143 11797
rect 12433 11792 13143 11794
rect 12433 11736 12438 11792
rect 12494 11736 13082 11792
rect 13138 11736 13143 11792
rect 12433 11734 13143 11736
rect 12433 11731 12499 11734
rect 13077 11731 13143 11734
rect 6729 11658 6795 11661
rect 27705 11658 27771 11661
rect 6729 11656 27771 11658
rect 6729 11600 6734 11656
rect 6790 11600 27710 11656
rect 27766 11600 27771 11656
rect 6729 11598 27771 11600
rect 6729 11595 6795 11598
rect 27705 11595 27771 11598
rect 4102 11460 4108 11524
rect 4172 11522 4178 11524
rect 5349 11522 5415 11525
rect 4172 11520 5415 11522
rect 4172 11464 5354 11520
rect 5410 11464 5415 11520
rect 4172 11462 5415 11464
rect 4172 11460 4178 11462
rect 5349 11459 5415 11462
rect 6913 11522 6979 11525
rect 9489 11522 9555 11525
rect 6913 11520 9555 11522
rect 6913 11464 6918 11520
rect 6974 11464 9494 11520
rect 9550 11464 9555 11520
rect 6913 11462 9555 11464
rect 6913 11459 6979 11462
rect 9489 11459 9555 11462
rect 11421 11524 11487 11525
rect 11421 11520 11468 11524
rect 11532 11522 11538 11524
rect 11421 11464 11426 11520
rect 11421 11460 11468 11464
rect 11532 11462 11578 11522
rect 11532 11460 11538 11462
rect 11421 11459 11487 11460
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 0 11326 2790 11386
rect 0 11296 800 11326
rect 2730 11250 2790 11326
rect 3366 11324 3372 11388
rect 3436 11386 3442 11388
rect 4153 11386 4219 11389
rect 11973 11386 12039 11389
rect 3436 11384 12039 11386
rect 3436 11328 4158 11384
rect 4214 11328 11978 11384
rect 12034 11328 12039 11384
rect 3436 11326 12039 11328
rect 3436 11324 3442 11326
rect 4153 11323 4219 11326
rect 11973 11323 12039 11326
rect 3509 11250 3575 11253
rect 2730 11248 3575 11250
rect 2730 11192 3514 11248
rect 3570 11192 3575 11248
rect 2730 11190 3575 11192
rect 3509 11187 3575 11190
rect 3693 11250 3759 11253
rect 19149 11250 19215 11253
rect 3693 11248 19215 11250
rect 3693 11192 3698 11248
rect 3754 11192 19154 11248
rect 19210 11192 19215 11248
rect 3693 11190 19215 11192
rect 3693 11187 3759 11190
rect 19149 11187 19215 11190
rect 4613 11116 4679 11117
rect 5441 11116 5507 11117
rect 4613 11114 4660 11116
rect 4568 11112 4660 11114
rect 4568 11056 4618 11112
rect 4568 11054 4660 11056
rect 4613 11052 4660 11054
rect 4724 11052 4730 11116
rect 5390 11052 5396 11116
rect 5460 11114 5507 11116
rect 7189 11114 7255 11117
rect 7598 11114 7604 11116
rect 5460 11112 5552 11114
rect 5502 11056 5552 11112
rect 5460 11054 5552 11056
rect 7189 11112 7604 11114
rect 7189 11056 7194 11112
rect 7250 11056 7604 11112
rect 7189 11054 7604 11056
rect 5460 11052 5507 11054
rect 4613 11051 4679 11052
rect 5441 11051 5507 11052
rect 7189 11051 7255 11054
rect 7598 11052 7604 11054
rect 7668 11052 7674 11116
rect 10041 11114 10107 11117
rect 11513 11114 11579 11117
rect 10041 11112 11579 11114
rect 10041 11056 10046 11112
rect 10102 11056 11518 11112
rect 11574 11056 11579 11112
rect 10041 11054 11579 11056
rect 10041 11051 10107 11054
rect 11513 11051 11579 11054
rect 12341 11114 12407 11117
rect 16481 11114 16547 11117
rect 12341 11112 16547 11114
rect 12341 11056 12346 11112
rect 12402 11056 16486 11112
rect 16542 11056 16547 11112
rect 12341 11054 16547 11056
rect 12341 11051 12407 11054
rect 16481 11051 16547 11054
rect 0 10978 800 11008
rect 1669 10978 1735 10981
rect 0 10976 1735 10978
rect 0 10920 1674 10976
rect 1730 10920 1735 10976
rect 0 10918 1735 10920
rect 0 10888 800 10918
rect 1669 10915 1735 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 12249 10842 12315 10845
rect 12893 10842 12959 10845
rect 13813 10842 13879 10845
rect 12249 10840 13879 10842
rect 12249 10784 12254 10840
rect 12310 10784 12898 10840
rect 12954 10784 13818 10840
rect 13874 10784 13879 10840
rect 12249 10782 13879 10784
rect 12249 10779 12315 10782
rect 12893 10779 12959 10782
rect 13813 10779 13879 10782
rect 2773 10706 2839 10709
rect 4429 10706 4495 10709
rect 7005 10706 7071 10709
rect 22134 10706 22140 10708
rect 2773 10704 6930 10706
rect 2773 10648 2778 10704
rect 2834 10648 4434 10704
rect 4490 10648 6930 10704
rect 2773 10646 6930 10648
rect 2773 10643 2839 10646
rect 4429 10643 4495 10646
rect 0 10570 800 10600
rect 2773 10570 2839 10573
rect 0 10568 2839 10570
rect 0 10512 2778 10568
rect 2834 10512 2839 10568
rect 0 10510 2839 10512
rect 6870 10570 6930 10646
rect 7005 10704 22140 10706
rect 7005 10648 7010 10704
rect 7066 10648 22140 10704
rect 7005 10646 22140 10648
rect 7005 10643 7071 10646
rect 22134 10644 22140 10646
rect 22204 10644 22210 10708
rect 11053 10570 11119 10573
rect 11513 10570 11579 10573
rect 6870 10568 11579 10570
rect 6870 10512 11058 10568
rect 11114 10512 11518 10568
rect 11574 10512 11579 10568
rect 6870 10510 11579 10512
rect 0 10480 800 10510
rect 2773 10507 2839 10510
rect 11053 10507 11119 10510
rect 11513 10507 11579 10510
rect 3693 10434 3759 10437
rect 7373 10434 7439 10437
rect 3693 10432 7439 10434
rect 3693 10376 3698 10432
rect 3754 10376 7378 10432
rect 7434 10376 7439 10432
rect 3693 10374 7439 10376
rect 3693 10371 3759 10374
rect 7373 10371 7439 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 42946 10303 43262 10304
rect 15469 10298 15535 10301
rect 16573 10298 16639 10301
rect 15469 10296 16639 10298
rect 15469 10240 15474 10296
rect 15530 10240 16578 10296
rect 16634 10240 16639 10296
rect 15469 10238 16639 10240
rect 15469 10235 15535 10238
rect 16573 10235 16639 10238
rect 0 10162 800 10192
rect 2865 10162 2931 10165
rect 0 10160 2931 10162
rect 0 10104 2870 10160
rect 2926 10104 2931 10160
rect 0 10102 2931 10104
rect 0 10072 800 10102
rect 2865 10099 2931 10102
rect 3417 10162 3483 10165
rect 3693 10164 3759 10165
rect 3550 10162 3556 10164
rect 3417 10160 3556 10162
rect 3417 10104 3422 10160
rect 3478 10104 3556 10160
rect 3417 10102 3556 10104
rect 3417 10099 3483 10102
rect 3550 10100 3556 10102
rect 3620 10100 3626 10164
rect 3693 10160 3740 10164
rect 3804 10162 3810 10164
rect 3693 10104 3698 10160
rect 3693 10100 3740 10104
rect 3804 10102 3850 10162
rect 3804 10100 3810 10102
rect 3693 10099 3759 10100
rect 6913 10026 6979 10029
rect 6913 10024 12450 10026
rect 6913 9968 6918 10024
rect 6974 9968 12450 10024
rect 6913 9966 12450 9968
rect 6913 9963 6979 9966
rect 11421 9892 11487 9893
rect 11421 9890 11468 9892
rect 11376 9888 11468 9890
rect 11376 9832 11426 9888
rect 11376 9830 11468 9832
rect 11421 9828 11468 9830
rect 11532 9828 11538 9892
rect 11421 9827 11487 9828
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 1577 9754 1643 9757
rect 0 9752 1643 9754
rect 0 9696 1582 9752
rect 1638 9696 1643 9752
rect 0 9694 1643 9696
rect 12390 9754 12450 9966
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 13854 9754 13860 9756
rect 12390 9694 13860 9754
rect 0 9664 800 9694
rect 1577 9691 1643 9694
rect 13854 9692 13860 9694
rect 13924 9692 13930 9756
rect 5533 9620 5599 9621
rect 5533 9616 5580 9620
rect 5644 9618 5650 9620
rect 5533 9560 5538 9616
rect 5533 9556 5580 9560
rect 5644 9558 5690 9618
rect 5644 9556 5650 9558
rect 6126 9556 6132 9620
rect 6196 9618 6202 9620
rect 6361 9618 6427 9621
rect 6196 9616 6427 9618
rect 6196 9560 6366 9616
rect 6422 9560 6427 9616
rect 6196 9558 6427 9560
rect 6196 9556 6202 9558
rect 5533 9555 5599 9556
rect 6361 9555 6427 9558
rect 6862 9556 6868 9620
rect 6932 9618 6938 9620
rect 8661 9618 8727 9621
rect 6932 9616 8727 9618
rect 6932 9560 8666 9616
rect 8722 9560 8727 9616
rect 6932 9558 8727 9560
rect 6932 9556 6938 9558
rect 8661 9555 8727 9558
rect 2262 9420 2268 9484
rect 2332 9482 2338 9484
rect 3601 9482 3667 9485
rect 2332 9480 3667 9482
rect 2332 9424 3606 9480
rect 3662 9424 3667 9480
rect 2332 9422 3667 9424
rect 2332 9420 2338 9422
rect 3601 9419 3667 9422
rect 12065 9482 12131 9485
rect 14733 9482 14799 9485
rect 17585 9482 17651 9485
rect 12065 9480 17651 9482
rect 12065 9424 12070 9480
rect 12126 9424 14738 9480
rect 14794 9424 17590 9480
rect 17646 9424 17651 9480
rect 12065 9422 17651 9424
rect 12065 9419 12131 9422
rect 14733 9419 14799 9422
rect 17585 9419 17651 9422
rect 0 9346 800 9376
rect 2773 9346 2839 9349
rect 0 9344 2839 9346
rect 0 9288 2778 9344
rect 2834 9288 2839 9344
rect 0 9286 2839 9288
rect 0 9256 800 9286
rect 2773 9283 2839 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 7741 9074 7807 9077
rect 24301 9074 24367 9077
rect 7741 9072 24367 9074
rect 7741 9016 7746 9072
rect 7802 9016 24306 9072
rect 24362 9016 24367 9072
rect 7741 9014 24367 9016
rect 7741 9011 7807 9014
rect 24301 9011 24367 9014
rect 0 8938 800 8968
rect 1761 8938 1827 8941
rect 0 8936 1827 8938
rect 0 8880 1766 8936
rect 1822 8880 1827 8936
rect 0 8878 1827 8880
rect 0 8848 800 8878
rect 1761 8875 1827 8878
rect 3325 8938 3391 8941
rect 22686 8938 22692 8940
rect 3325 8936 22692 8938
rect 3325 8880 3330 8936
rect 3386 8880 22692 8936
rect 3325 8878 22692 8880
rect 3325 8875 3391 8878
rect 22686 8876 22692 8878
rect 22756 8876 22762 8940
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 6637 8668 6703 8669
rect 6637 8666 6684 8668
rect 6592 8664 6684 8666
rect 6592 8608 6642 8664
rect 6592 8606 6684 8608
rect 6637 8604 6684 8606
rect 6748 8604 6754 8668
rect 6637 8603 6703 8604
rect 0 8530 800 8560
rect 2865 8530 2931 8533
rect 0 8528 2931 8530
rect 0 8472 2870 8528
rect 2926 8472 2931 8528
rect 0 8470 2931 8472
rect 0 8440 800 8470
rect 2865 8467 2931 8470
rect 4245 8530 4311 8533
rect 8334 8530 8340 8532
rect 4245 8528 8340 8530
rect 4245 8472 4250 8528
rect 4306 8472 8340 8528
rect 4245 8470 8340 8472
rect 4245 8467 4311 8470
rect 8334 8468 8340 8470
rect 8404 8468 8410 8532
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 2773 8122 2839 8125
rect 0 8120 2839 8122
rect 0 8064 2778 8120
rect 2834 8064 2839 8120
rect 0 8062 2839 8064
rect 0 8032 800 8062
rect 2773 8059 2839 8062
rect 2221 7850 2287 7853
rect 8518 7850 8524 7852
rect 2221 7848 8524 7850
rect 2221 7792 2226 7848
rect 2282 7792 8524 7848
rect 2221 7790 8524 7792
rect 2221 7787 2287 7790
rect 8518 7788 8524 7790
rect 8588 7788 8594 7852
rect 0 7714 800 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 800 7654
rect 1301 7651 1367 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 0 7306 800 7336
rect 2865 7306 2931 7309
rect 0 7304 2931 7306
rect 0 7248 2870 7304
rect 2926 7248 2931 7304
rect 0 7246 2931 7248
rect 0 7216 800 7246
rect 2865 7243 2931 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 0 6898 800 6928
rect 3601 6898 3667 6901
rect 0 6896 3667 6898
rect 0 6840 3606 6896
rect 3662 6840 3667 6896
rect 0 6838 3667 6840
rect 0 6808 800 6838
rect 3601 6835 3667 6838
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1301 6490 1367 6493
rect 0 6488 1367 6490
rect 0 6432 1306 6488
rect 1362 6432 1367 6488
rect 0 6430 1367 6432
rect 0 6400 800 6430
rect 1301 6427 1367 6430
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 1301 5266 1367 5269
rect 0 5264 1367 5266
rect 0 5208 1306 5264
rect 1362 5208 1367 5264
rect 0 5206 1367 5208
rect 0 5176 800 5206
rect 1301 5203 1367 5206
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 0 4450 800 4480
rect 4153 4450 4219 4453
rect 0 4448 4219 4450
rect 0 4392 4158 4448
rect 4214 4392 4219 4448
rect 0 4390 4219 4392
rect 0 4360 800 4390
rect 4153 4387 4219 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 0 4042 800 4072
rect 4061 4042 4127 4045
rect 0 4040 4127 4042
rect 0 3984 4066 4040
rect 4122 3984 4127 4040
rect 0 3982 4127 3984
rect 0 3952 800 3982
rect 4061 3979 4127 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 2865 3634 2931 3637
rect 0 3632 2931 3634
rect 0 3576 2870 3632
rect 2926 3576 2931 3632
rect 0 3574 2931 3576
rect 0 3544 800 3574
rect 2865 3571 2931 3574
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 1301 3226 1367 3229
rect 0 3224 1367 3226
rect 0 3168 1306 3224
rect 1362 3168 1367 3224
rect 0 3166 1367 3168
rect 0 3136 800 3166
rect 1301 3163 1367 3166
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 0 2410 800 2440
rect 1209 2410 1275 2413
rect 0 2408 1275 2410
rect 0 2352 1214 2408
rect 1270 2352 1275 2408
rect 0 2350 1275 2352
rect 0 2320 800 2350
rect 1209 2347 1275 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 1301 2002 1367 2005
rect 0 2000 1367 2002
rect 0 1944 1306 2000
rect 1362 1944 1367 2000
rect 0 1942 1367 1944
rect 0 1912 800 1942
rect 1301 1939 1367 1942
rect 0 1594 800 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 800 1534
rect 2865 1531 2931 1534
<< via3 >>
rect 16988 24924 17052 24988
rect 14412 24516 14476 24580
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 5580 24108 5644 24172
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 4292 23564 4356 23628
rect 2268 23428 2332 23492
rect 5396 23428 5460 23492
rect 7604 23428 7668 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 5580 23156 5644 23220
rect 22140 23216 22204 23220
rect 22140 23160 22190 23216
rect 22190 23160 22204 23216
rect 22140 23156 22204 23160
rect 4660 22884 4724 22948
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 17172 22748 17236 22812
rect 4108 22536 4172 22540
rect 4108 22480 4158 22536
rect 4158 22480 4172 22536
rect 4108 22476 4172 22480
rect 17172 22476 17236 22540
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 6684 22128 6748 22132
rect 6684 22072 6698 22128
rect 6698 22072 6748 22128
rect 6684 22068 6748 22072
rect 14412 21992 14476 21996
rect 14412 21936 14426 21992
rect 14426 21936 14476 21992
rect 14412 21932 14476 21936
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 3924 21720 3988 21724
rect 3924 21664 3974 21720
rect 3974 21664 3988 21720
rect 3924 21660 3988 21664
rect 22692 21660 22756 21724
rect 5948 21252 6012 21316
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 5764 20768 5828 20772
rect 5764 20712 5778 20768
rect 5778 20712 5828 20768
rect 5764 20708 5828 20712
rect 6868 20768 6932 20772
rect 6868 20712 6918 20768
rect 6918 20712 6932 20768
rect 6868 20708 6932 20712
rect 7052 20708 7116 20772
rect 10548 20708 10612 20772
rect 11100 20708 11164 20772
rect 13860 20768 13924 20772
rect 13860 20712 13910 20768
rect 13910 20712 13924 20768
rect 13860 20708 13924 20712
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 9628 19348 9692 19412
rect 7420 19212 7484 19276
rect 17540 19076 17604 19140
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 3740 18940 3804 19004
rect 3556 18668 3620 18732
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 6132 18456 6196 18460
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 6132 18400 6146 18456
rect 6146 18400 6196 18456
rect 6132 18396 6196 18400
rect 3372 17988 3436 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 5948 17444 6012 17508
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 18460 17172 18524 17236
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 5764 16628 5828 16692
rect 8524 16628 8588 16692
rect 8340 16492 8404 16556
rect 16988 16416 17052 16420
rect 16988 16360 17002 16416
rect 17002 16360 17052 16416
rect 16988 16356 17052 16360
rect 17540 16416 17604 16420
rect 17540 16360 17554 16416
rect 17554 16360 17604 16416
rect 17540 16356 17604 16360
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 9628 16220 9692 16284
rect 17172 16280 17236 16284
rect 17172 16224 17186 16280
rect 17186 16224 17236 16280
rect 17172 16220 17236 16224
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 9812 15812 9876 15876
rect 10548 15812 10612 15876
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 3924 15540 3988 15604
rect 3924 15404 3988 15468
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 6132 13092 6196 13156
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 18460 12684 18524 12748
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 11100 12412 11164 12476
rect 3924 12276 3988 12340
rect 4292 12336 4356 12340
rect 4292 12280 4306 12336
rect 4306 12280 4356 12336
rect 4292 12276 4356 12280
rect 7420 12336 7484 12340
rect 7420 12280 7434 12336
rect 7434 12280 7484 12336
rect 7420 12276 7484 12280
rect 9812 12140 9876 12204
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 7052 11868 7116 11932
rect 4108 11460 4172 11524
rect 11468 11520 11532 11524
rect 11468 11464 11482 11520
rect 11482 11464 11532 11520
rect 11468 11460 11532 11464
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 3372 11324 3436 11388
rect 4660 11112 4724 11116
rect 4660 11056 4674 11112
rect 4674 11056 4724 11112
rect 4660 11052 4724 11056
rect 5396 11112 5460 11116
rect 5396 11056 5446 11112
rect 5446 11056 5460 11112
rect 5396 11052 5460 11056
rect 7604 11052 7668 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 22140 10644 22204 10708
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 3556 10100 3620 10164
rect 3740 10160 3804 10164
rect 3740 10104 3754 10160
rect 3754 10104 3804 10160
rect 3740 10100 3804 10104
rect 11468 9888 11532 9892
rect 11468 9832 11482 9888
rect 11482 9832 11532 9888
rect 11468 9828 11532 9832
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 13860 9692 13924 9756
rect 5580 9616 5644 9620
rect 5580 9560 5594 9616
rect 5594 9560 5644 9616
rect 5580 9556 5644 9560
rect 6132 9556 6196 9620
rect 6868 9556 6932 9620
rect 2268 9420 2332 9484
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 22692 8876 22756 8940
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 6684 8664 6748 8668
rect 6684 8608 6698 8664
rect 6698 8608 6748 8664
rect 6684 8604 6748 8608
rect 8340 8468 8404 8532
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 8524 7788 8588 7852
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 16987 24988 17053 24989
rect 16987 24924 16988 24988
rect 17052 24924 17053 24988
rect 16987 24923 17053 24924
rect 14411 24580 14477 24581
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2267 23492 2333 23493
rect 2267 23428 2268 23492
rect 2332 23428 2333 23492
rect 2267 23427 2333 23428
rect 2270 9485 2330 23427
rect 2944 23424 3264 24448
rect 5579 24172 5645 24173
rect 5579 24108 5580 24172
rect 5644 24108 5645 24172
rect 5579 24107 5645 24108
rect 4291 23628 4357 23629
rect 4291 23564 4292 23628
rect 4356 23564 4357 23628
rect 4291 23563 4357 23564
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 4107 22540 4173 22541
rect 4107 22476 4108 22540
rect 4172 22476 4173 22540
rect 4107 22475 4173 22476
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 3923 21724 3989 21725
rect 3923 21660 3924 21724
rect 3988 21660 3989 21724
rect 3923 21659 3989 21660
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 3739 19004 3805 19005
rect 3739 18940 3740 19004
rect 3804 18940 3805 19004
rect 3739 18939 3805 18940
rect 3555 18732 3621 18733
rect 3555 18668 3556 18732
rect 3620 18668 3621 18732
rect 3555 18667 3621 18668
rect 3371 18052 3437 18053
rect 3371 17988 3372 18052
rect 3436 17988 3437 18052
rect 3371 17987 3437 17988
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 3374 11389 3434 17987
rect 3371 11388 3437 11389
rect 3371 11324 3372 11388
rect 3436 11324 3437 11388
rect 3371 11323 3437 11324
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2267 9484 2333 9485
rect 2267 9420 2268 9484
rect 2332 9420 2333 9484
rect 2267 9419 2333 9420
rect 2944 9280 3264 10304
rect 3558 10165 3618 18667
rect 3742 10165 3802 18939
rect 3926 15605 3986 21659
rect 3923 15604 3989 15605
rect 3923 15540 3924 15604
rect 3988 15540 3989 15604
rect 3923 15539 3989 15540
rect 3923 15468 3989 15469
rect 3923 15404 3924 15468
rect 3988 15404 3989 15468
rect 3923 15403 3989 15404
rect 3926 12341 3986 15403
rect 3923 12340 3989 12341
rect 3923 12276 3924 12340
rect 3988 12276 3989 12340
rect 3923 12275 3989 12276
rect 4110 11525 4170 22475
rect 4294 12341 4354 23563
rect 5395 23492 5461 23493
rect 5395 23428 5396 23492
rect 5460 23428 5461 23492
rect 5395 23427 5461 23428
rect 4659 22948 4725 22949
rect 4659 22884 4660 22948
rect 4724 22884 4725 22948
rect 4659 22883 4725 22884
rect 4291 12340 4357 12341
rect 4291 12276 4292 12340
rect 4356 12276 4357 12340
rect 4291 12275 4357 12276
rect 4107 11524 4173 11525
rect 4107 11460 4108 11524
rect 4172 11460 4173 11524
rect 4107 11459 4173 11460
rect 4662 11117 4722 22883
rect 5398 11117 5458 23427
rect 5582 23221 5642 24107
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7603 23492 7669 23493
rect 7603 23428 7604 23492
rect 7668 23428 7669 23492
rect 7603 23427 7669 23428
rect 5579 23220 5645 23221
rect 5579 23156 5580 23220
rect 5644 23156 5645 23220
rect 5579 23155 5645 23156
rect 4659 11116 4725 11117
rect 4659 11052 4660 11116
rect 4724 11052 4725 11116
rect 4659 11051 4725 11052
rect 5395 11116 5461 11117
rect 5395 11052 5396 11116
rect 5460 11052 5461 11116
rect 5395 11051 5461 11052
rect 3555 10164 3621 10165
rect 3555 10100 3556 10164
rect 3620 10100 3621 10164
rect 3555 10099 3621 10100
rect 3739 10164 3805 10165
rect 3739 10100 3740 10164
rect 3804 10100 3805 10164
rect 3739 10099 3805 10100
rect 5582 9621 5642 23155
rect 6683 22132 6749 22133
rect 6683 22068 6684 22132
rect 6748 22068 6749 22132
rect 6683 22067 6749 22068
rect 5947 21316 6013 21317
rect 5947 21252 5948 21316
rect 6012 21252 6013 21316
rect 5947 21251 6013 21252
rect 5763 20772 5829 20773
rect 5763 20708 5764 20772
rect 5828 20708 5829 20772
rect 5763 20707 5829 20708
rect 5766 16693 5826 20707
rect 5950 17509 6010 21251
rect 6686 19350 6746 22067
rect 6867 20772 6933 20773
rect 6867 20708 6868 20772
rect 6932 20708 6933 20772
rect 6867 20707 6933 20708
rect 7051 20772 7117 20773
rect 7051 20708 7052 20772
rect 7116 20708 7117 20772
rect 7051 20707 7117 20708
rect 6318 19290 6746 19350
rect 6131 18460 6197 18461
rect 6131 18396 6132 18460
rect 6196 18396 6197 18460
rect 6131 18395 6197 18396
rect 5947 17508 6013 17509
rect 5947 17444 5948 17508
rect 6012 17444 6013 17508
rect 5947 17443 6013 17444
rect 5763 16692 5829 16693
rect 5763 16628 5764 16692
rect 5828 16628 5829 16692
rect 5763 16627 5829 16628
rect 6134 13157 6194 18395
rect 6131 13156 6197 13157
rect 6131 13092 6132 13156
rect 6196 13092 6197 13156
rect 6131 13091 6197 13092
rect 6134 9621 6194 13091
rect 6318 9690 6378 19290
rect 6318 9630 6746 9690
rect 5579 9620 5645 9621
rect 5579 9556 5580 9620
rect 5644 9556 5645 9620
rect 5579 9555 5645 9556
rect 6131 9620 6197 9621
rect 6131 9556 6132 9620
rect 6196 9556 6197 9620
rect 6131 9555 6197 9556
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 6686 8669 6746 9630
rect 6870 9621 6930 20707
rect 7054 11933 7114 20707
rect 7419 19276 7485 19277
rect 7419 19212 7420 19276
rect 7484 19212 7485 19276
rect 7419 19211 7485 19212
rect 7422 12341 7482 19211
rect 7419 12340 7485 12341
rect 7419 12276 7420 12340
rect 7484 12276 7485 12340
rect 7419 12275 7485 12276
rect 7051 11932 7117 11933
rect 7051 11868 7052 11932
rect 7116 11868 7117 11932
rect 7051 11867 7117 11868
rect 7606 11117 7666 23427
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 12944 24512 13264 24528
rect 14411 24516 14412 24580
rect 14476 24516 14477 24580
rect 14411 24515 14477 24516
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 14414 21997 14474 24515
rect 14411 21996 14477 21997
rect 14411 21932 14412 21996
rect 14476 21932 14477 21996
rect 14411 21931 14477 21932
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 10547 20772 10613 20773
rect 10547 20708 10548 20772
rect 10612 20708 10613 20772
rect 10547 20707 10613 20708
rect 11099 20772 11165 20773
rect 11099 20708 11100 20772
rect 11164 20708 11165 20772
rect 11099 20707 11165 20708
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 9627 19412 9693 19413
rect 9627 19348 9628 19412
rect 9692 19348 9693 19412
rect 9627 19347 9693 19348
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 8523 16692 8589 16693
rect 8523 16628 8524 16692
rect 8588 16628 8589 16692
rect 8523 16627 8589 16628
rect 8339 16556 8405 16557
rect 8339 16492 8340 16556
rect 8404 16492 8405 16556
rect 8339 16491 8405 16492
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7603 11116 7669 11117
rect 7603 11052 7604 11116
rect 7668 11052 7669 11116
rect 7603 11051 7669 11052
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 6867 9620 6933 9621
rect 6867 9556 6868 9620
rect 6932 9556 6933 9620
rect 6867 9555 6933 9556
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 6683 8668 6749 8669
rect 6683 8604 6684 8668
rect 6748 8604 6749 8668
rect 6683 8603 6749 8604
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 7648 8264 8672
rect 8342 8533 8402 16491
rect 8339 8532 8405 8533
rect 8339 8468 8340 8532
rect 8404 8468 8405 8532
rect 8339 8467 8405 8468
rect 8526 7853 8586 16627
rect 9630 16285 9690 19347
rect 9627 16284 9693 16285
rect 9627 16220 9628 16284
rect 9692 16220 9693 16284
rect 9627 16219 9693 16220
rect 10550 15877 10610 20707
rect 9811 15876 9877 15877
rect 9811 15812 9812 15876
rect 9876 15812 9877 15876
rect 9811 15811 9877 15812
rect 10547 15876 10613 15877
rect 10547 15812 10548 15876
rect 10612 15812 10613 15876
rect 10547 15811 10613 15812
rect 9814 12205 9874 15811
rect 11102 12477 11162 20707
rect 12944 20160 13264 21184
rect 13859 20772 13925 20773
rect 13859 20708 13860 20772
rect 13924 20708 13925 20772
rect 13859 20707 13925 20708
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 11099 12476 11165 12477
rect 11099 12412 11100 12476
rect 11164 12412 11165 12476
rect 11099 12411 11165 12412
rect 9811 12204 9877 12205
rect 9811 12140 9812 12204
rect 9876 12140 9877 12204
rect 9811 12139 9877 12140
rect 11467 11524 11533 11525
rect 11467 11460 11468 11524
rect 11532 11460 11533 11524
rect 11467 11459 11533 11460
rect 11470 9893 11530 11459
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 11467 9892 11533 9893
rect 11467 9828 11468 9892
rect 11532 9828 11533 9892
rect 11467 9827 11533 9828
rect 12944 9280 13264 10304
rect 13862 9757 13922 20707
rect 16990 16421 17050 24923
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22139 23220 22205 23221
rect 22139 23156 22140 23220
rect 22204 23156 22205 23220
rect 22139 23155 22205 23156
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17171 22812 17237 22813
rect 17171 22748 17172 22812
rect 17236 22748 17237 22812
rect 17171 22747 17237 22748
rect 17174 22541 17234 22747
rect 17171 22540 17237 22541
rect 17171 22476 17172 22540
rect 17236 22476 17237 22540
rect 17171 22475 17237 22476
rect 16987 16420 17053 16421
rect 16987 16356 16988 16420
rect 17052 16356 17053 16420
rect 16987 16355 17053 16356
rect 17174 16285 17234 22475
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17539 19140 17605 19141
rect 17539 19076 17540 19140
rect 17604 19076 17605 19140
rect 17539 19075 17605 19076
rect 17542 16421 17602 19075
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17539 16420 17605 16421
rect 17539 16356 17540 16420
rect 17604 16356 17605 16420
rect 17539 16355 17605 16356
rect 17944 16352 18264 17376
rect 18459 17236 18525 17237
rect 18459 17172 18460 17236
rect 18524 17172 18525 17236
rect 18459 17171 18525 17172
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17171 16284 17237 16285
rect 17171 16220 17172 16284
rect 17236 16220 17237 16284
rect 17171 16219 17237 16220
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 18462 12749 18522 17171
rect 18459 12748 18525 12749
rect 18459 12684 18460 12748
rect 18524 12684 18525 12748
rect 18459 12683 18525 12684
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 22142 10709 22202 23155
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22691 21724 22757 21725
rect 22691 21660 22692 21724
rect 22756 21660 22757 21724
rect 22691 21659 22757 21660
rect 22139 10708 22205 10709
rect 22139 10644 22140 10708
rect 22204 10644 22205 10708
rect 22139 10643 22205 10644
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 13859 9756 13925 9757
rect 13859 9692 13860 9756
rect 13924 9692 13925 9756
rect 13859 9691 13925 9692
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 8523 7852 8589 7853
rect 8523 7788 8524 7852
rect 8588 7788 8589 7852
rect 8523 7787 8589 7788
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 8736 18264 9760
rect 22694 8941 22754 21659
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22691 8940 22757 8941
rect 22691 8876 22692 8940
rect 22756 8876 22757 8940
rect 22691 8875 22757 8876
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _096_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22448 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1676037725
transform 1 0 19504 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _099_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _100_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _101_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1676037725
transform 1 0 10672 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1676037725
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 6900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1676037725
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1676037725
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 4140 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 5796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1676037725
transform 1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 8464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1676037725
transform 1 0 3404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform 1 0 6072 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1676037725
transform 1 0 3496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1676037725
transform 1 0 4232 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1676037725
transform 1 0 20884 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _132_
timestamp 1676037725
transform 1 0 8372 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _133_
timestamp 1676037725
transform 1 0 2208 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _134_
timestamp 1676037725
transform 1 0 5888 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _135_
timestamp 1676037725
transform 1 0 3404 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _136_
timestamp 1676037725
transform 1 0 4232 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 33856 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 35328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 33764 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 32292 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 31280 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 34592 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 33028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _146_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _147_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _149_
timestamp 1676037725
transform 1 0 28244 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _150_
timestamp 1676037725
transform 1 0 18584 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _151_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _152_
timestamp 1676037725
transform 1 0 33580 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 11408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1676037725
transform 1 0 14996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1676037725
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 12328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 4508 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 3956 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 5612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 7636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 20700 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 10212 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 3036 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 4876 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1676037725
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1676037725
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1676037725
transform 1 0 3864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1676037725
transform 1 0 3312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1676037725
transform 1 0 1656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1676037725
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1676037725
transform 1 0 7636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1676037725
transform 1 0 4232 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1676037725
transform 1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1676037725
transform 1 0 2852 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1676037725
transform 1 0 11592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1676037725
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1676037725
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1676037725
transform 1 0 1748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1676037725
transform 1 0 9752 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1676037725
transform 1 0 3128 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1676037725
transform 1 0 33672 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform 1 0 33856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 32200 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform 1 0 35052 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1676037725
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1676037725
transform 1 0 22448 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1676037725
transform 1 0 31556 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1676037725
transform 1 0 7452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1676037725
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1676037725
transform 1 0 16008 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1676037725
transform 1 0 11960 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 9016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 6440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 6440 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 9108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 6440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 3312 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 11592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 11132 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 4784 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 4600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 5336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 10028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 9016 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__S
timestamp 1676037725
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 3036 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 5152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 2668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 10580 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 9016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 6440 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 3312 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 11592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 9844 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 6348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 13800 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 20148 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 21620 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR_A
timestamp 1676037725
transform 1 0 22816 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
timestamp 1676037725
transform 1 0 28520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 28336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE_TE_B
timestamp 1676037725
transform 1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 32016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 19320 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 9016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 9752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform 1 0 15916 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 16284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform 1 0 14996 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform 1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 19320 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 22724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 18308 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 21988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform 1 0 23276 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 26496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1676037725
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold10_A
timestamp 1676037725
transform 1 0 47380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold12_A
timestamp 1676037725
transform 1 0 2852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform 1 0 3404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform 1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform 1 0 4140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform 1 0 3312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform 1 0 3956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform 1 0 4416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform 1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform 1 0 4140 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform 1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform 1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform 1 0 4600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 4324 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 2668 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform 1 0 4600 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform 1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform 1 0 4416 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform 1 0 4508 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform 1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform 1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform 1 0 34868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 36984 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform 1 0 33396 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform 1 0 33580 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform 1 0 35328 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform 1 0 34224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform 1 0 36616 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform 1 0 34684 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform 1 0 37904 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform 1 0 36984 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform 1 0 31832 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform 1 0 38548 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 36800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform 1 0 37260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 38180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 38916 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 39836 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 40296 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform 1 0 41768 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform 1 0 5520 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform 1 0 32752 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform 1 0 33396 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform 1 0 25944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform 1 0 28612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform 1 0 31280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform 1 0 33948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform 1 0 46276 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform 1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform 1 0 47564 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform 1 0 44620 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform 1 0 46092 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform 1 0 47932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform 1 0 47748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output81_A
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1676037725
transform 1 0 1748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output114_A
timestamp 1676037725
transform 1 0 6716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output115_A
timestamp 1676037725
transform 1 0 7728 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output116_A
timestamp 1676037725
transform 1 0 3312 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output117_A
timestamp 1676037725
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output118_A
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1676037725
transform 1 0 17020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1676037725
transform 1 0 8464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1676037725
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 1676037725
transform 1 0 10856 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output131_A
timestamp 1676037725
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output142_A
timestamp 1676037725
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23920 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20884 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14904 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 21896 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22080 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26312 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 26496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 27232 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 27876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 25668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 30912 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 30820 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 31740 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31740 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 30728 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 31740 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 31740 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 34316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 31556 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 32844 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 27692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 31740 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 30912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 30728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 37444 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1676037725
transform 1 0 21620 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22908 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22172 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24196 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21896 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20056 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13892 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 5060 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 4140 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 3312 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 1472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15088 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15916 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 30360 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 27600 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15180 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16652 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 12328 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 22264 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23920 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14168 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14168 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 3312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 36800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_15.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 31924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_17.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 30544 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_19.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_29.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 27876 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 9936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_31.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 33028 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_45.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 32016 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_47.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_49.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_51.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 30728 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 31280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 31464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 30912 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 30544 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 19688 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 25576 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 26772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l2_in_0__S
timestamp 1676037725
transform 1 0 26128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l2_in_1__S
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 11592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 25668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26220 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 26404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 15364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24288 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25944 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 14076 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21528 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19504 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22724 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21896 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 11592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 27416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15456 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14168 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 3864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 11592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 30176 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 11592 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 32936 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 31096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 10488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 19872 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_38.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 5704 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16192 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 1472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 32844 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 8280 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 33028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22448 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20792 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9292 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6808 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4140 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 4140 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 4784 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 5336 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 5428 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 7360 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8004 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8464 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6808 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 6624 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 11224 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9200 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9568 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 10304 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__190 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 7820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 10304 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 4048 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 3404 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 9476 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 4232 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6348 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 6808 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__191
timestamp 1676037725
transform 1 0 5796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 5244 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 4048 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10580 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 3956 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 5152 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14260 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__192
timestamp 1676037725
transform 1 0 16468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 8096 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10396 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9384 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7820 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10856 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9384 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__193
timestamp 1676037725
transform 1 0 11868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 6716 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10580 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28612 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8740 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 26956 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22724 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 25760 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 22908 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22172 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 24656 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27508 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17112 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9568 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 14720 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 8464 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 13616 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 12788 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 19504 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 18952 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 23092 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 19596 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 24932 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 25300 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1676037725
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1676037725
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 1676037725
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1676037725
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1676037725
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_268
timestamp 1676037725
transform 1 0 25760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1676037725
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_297
timestamp 1676037725
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1676037725
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1676037725
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1676037725
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1676037725
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1676037725
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1676037725
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_395
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_407
timestamp 1676037725
transform 1 0 38548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1676037725
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1676037725
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1676037725
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1676037725
transform 1 0 48668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_34
timestamp 1676037725
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_67
timestamp 1676037725
transform 1 0 7268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_79
timestamp 1676037725
transform 1 0 8372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_103
timestamp 1676037725
transform 1 0 10580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1676037725
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_128
timestamp 1676037725
transform 1 0 12880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1676037725
transform 1 0 13616 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_142
timestamp 1676037725
transform 1 0 14168 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1676037725
transform 1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1676037725
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_174
timestamp 1676037725
transform 1 0 17112 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_182
timestamp 1676037725
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_188
timestamp 1676037725
transform 1 0 18400 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_200
timestamp 1676037725
transform 1 0 19504 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_208
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_212
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1676037725
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1676037725
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_19
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1676037725
transform 1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_34
timestamp 1676037725
transform 1 0 4232 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_40
timestamp 1676037725
transform 1 0 4784 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_52
timestamp 1676037725
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_64
timestamp 1676037725
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 1676037725
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1676037725
transform 1 0 11776 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_120
timestamp 1676037725
transform 1 0 12144 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1676037725
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1676037725
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_5
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_16
timestamp 1676037725
transform 1 0 2576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_28
timestamp 1676037725
transform 1 0 3680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1676037725
transform 1 0 4324 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_154
timestamp 1676037725
transform 1 0 15272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1676037725
transform 1 0 3128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1676037725
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_205
timestamp 1676037725
transform 1 0 19964 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_258
timestamp 1676037725
transform 1 0 24840 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_266
timestamp 1676037725
transform 1 0 25576 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1676037725
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1676037725
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1676037725
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1676037725
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1676037725
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_157
timestamp 1676037725
transform 1 0 15548 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_177
timestamp 1676037725
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_186
timestamp 1676037725
transform 1 0 18216 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_198
timestamp 1676037725
transform 1 0 19320 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_210
timestamp 1676037725
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_231
timestamp 1676037725
transform 1 0 22356 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_238
timestamp 1676037725
transform 1 0 23000 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_250
timestamp 1676037725
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_262
timestamp 1676037725
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1676037725
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_320
timestamp 1676037725
transform 1 0 30544 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1676037725
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1676037725
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_173
timestamp 1676037725
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_199
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_211
timestamp 1676037725
transform 1 0 20516 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_225
timestamp 1676037725
transform 1 0 21804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_237
timestamp 1676037725
transform 1 0 22908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1676037725
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_302
timestamp 1676037725
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_22
timestamp 1676037725
transform 1 0 3128 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_26
timestamp 1676037725
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_38
timestamp 1676037725
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1676037725
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_234
timestamp 1676037725
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_238
timestamp 1676037725
transform 1 0 23000 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_250
timestamp 1676037725
transform 1 0 24104 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_262
timestamp 1676037725
transform 1 0 25208 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_274
timestamp 1676037725
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1676037725
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_22
timestamp 1676037725
transform 1 0 3128 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_35
timestamp 1676037725
transform 1 0 4324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_47
timestamp 1676037725
transform 1 0 5428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_59
timestamp 1676037725
transform 1 0 6532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_71
timestamp 1676037725
transform 1 0 7636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_106
timestamp 1676037725
transform 1 0 10856 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_118
timestamp 1676037725
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 1676037725
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_243
timestamp 1676037725
transform 1 0 23460 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_247
timestamp 1676037725
transform 1 0 23828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1676037725
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_22
timestamp 1676037725
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_29
timestamp 1676037725
transform 1 0 3772 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 1676037725
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1676037725
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_90
timestamp 1676037725
transform 1 0 9384 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1676037725
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1676037725
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_120
timestamp 1676037725
transform 1 0 12144 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_127
timestamp 1676037725
transform 1 0 12788 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_133
timestamp 1676037725
transform 1 0 13340 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_144
timestamp 1676037725
transform 1 0 14352 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_156
timestamp 1676037725
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1676037725
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1676037725
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1676037725
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1676037725
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1676037725
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_8
timestamp 1676037725
transform 1 0 1840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1676037725
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp 1676037725
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_40
timestamp 1676037725
transform 1 0 4784 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_52
timestamp 1676037725
transform 1 0 5888 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_64
timestamp 1676037725
transform 1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_68
timestamp 1676037725
transform 1 0 7360 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1676037725
transform 1 0 7636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 1676037725
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1676037725
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_101
timestamp 1676037725
transform 1 0 10396 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_120
timestamp 1676037725
transform 1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_128
timestamp 1676037725
transform 1 0 12880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_143
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1676037725
transform 1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_161
timestamp 1676037725
transform 1 0 15916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_173
timestamp 1676037725
transform 1 0 17020 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1676037725
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1676037725
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_22
timestamp 1676037725
transform 1 0 3128 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_28
timestamp 1676037725
transform 1 0 3680 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 1676037725
transform 1 0 4232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1676037725
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_45
timestamp 1676037725
transform 1 0 5244 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_63
timestamp 1676037725
transform 1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1676037725
transform 1 0 8188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_89
timestamp 1676037725
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_96
timestamp 1676037725
transform 1 0 9936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_107
timestamp 1676037725
transform 1 0 10948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp 1676037725
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_129
timestamp 1676037725
transform 1 0 12972 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1676037725
transform 1 0 13524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1676037725
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1676037725
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_156
timestamp 1676037725
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1676037725
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1676037725
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1676037725
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1676037725
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_22
timestamp 1676037725
transform 1 0 3128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_34
timestamp 1676037725
transform 1 0 4232 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_42
timestamp 1676037725
transform 1 0 4968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_50
timestamp 1676037725
transform 1 0 5704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1676037725
transform 1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1676037725
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1676037725
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1676037725
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1676037725
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_107
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_128
timestamp 1676037725
transform 1 0 12880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1676037725
transform 1 0 13432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 1676037725
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_161
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1676037725
transform 1 0 17848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1676037725
transform 1 0 18584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_193
timestamp 1676037725
transform 1 0 18860 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1676037725
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1676037725
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1676037725
transform 1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_19
timestamp 1676037725
transform 1 0 2852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_24
timestamp 1676037725
transform 1 0 3312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_30
timestamp 1676037725
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_44
timestamp 1676037725
transform 1 0 5152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_60
timestamp 1676037725
transform 1 0 6624 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1676037725
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1676037725
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_135
timestamp 1676037725
transform 1 0 13524 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1676037725
transform 1 0 14260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1676037725
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_191
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1676037725
transform 1 0 19872 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_208
timestamp 1676037725
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1676037725
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_294
timestamp 1676037725
transform 1 0 28152 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_300
timestamp 1676037725
transform 1 0 28704 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_312
timestamp 1676037725
transform 1 0 29808 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_324
timestamp 1676037725
transform 1 0 30912 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1676037725
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1676037725
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1676037725
transform 1 0 4048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_44
timestamp 1676037725
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_48
timestamp 1676037725
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_54
timestamp 1676037725
transform 1 0 6072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_60
timestamp 1676037725
transform 1 0 6624 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1676037725
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1676037725
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_106
timestamp 1676037725
transform 1 0 10856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1676037725
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_134
timestamp 1676037725
transform 1 0 13432 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_143
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_172
timestamp 1676037725
transform 1 0 16928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_219
timestamp 1676037725
transform 1 0 21252 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_225
timestamp 1676037725
transform 1 0 21804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_237
timestamp 1676037725
transform 1 0 22908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1676037725
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1676037725
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1676037725
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1676037725
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1676037725
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1676037725
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1676037725
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1676037725
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1676037725
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1676037725
transform 1 0 1932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1676037725
transform 1 0 3036 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_42
timestamp 1676037725
transform 1 0 4968 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_60
timestamp 1676037725
transform 1 0 6624 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 1676037725
transform 1 0 7084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1676037725
transform 1 0 9568 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1676037725
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1676037725
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_116
timestamp 1676037725
transform 1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_139
timestamp 1676037725
transform 1 0 13892 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_143
timestamp 1676037725
transform 1 0 14260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_229
timestamp 1676037725
transform 1 0 22172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_241
timestamp 1676037725
transform 1 0 23276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_253
timestamp 1676037725
transform 1 0 24380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_265
timestamp 1676037725
transform 1 0 25484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1676037725
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1676037725
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1676037725
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1676037725
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1676037725
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1676037725
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1676037725
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1676037725
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1676037725
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1676037725
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_517
timestamp 1676037725
transform 1 0 48668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_8
timestamp 1676037725
transform 1 0 1840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_22
timestamp 1676037725
transform 1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_35
timestamp 1676037725
transform 1 0 4324 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_39
timestamp 1676037725
transform 1 0 4692 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_60
timestamp 1676037725
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_67
timestamp 1676037725
transform 1 0 7268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1676037725
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_96
timestamp 1676037725
transform 1 0 9936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_143
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_168
timestamp 1676037725
transform 1 0 16560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_172
timestamp 1676037725
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_211
timestamp 1676037725
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_235
timestamp 1676037725
transform 1 0 22724 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_239
timestamp 1676037725
transform 1 0 23092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1676037725
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1676037725
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_334
timestamp 1676037725
transform 1 0 31832 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_338
timestamp 1676037725
transform 1 0 32200 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_350
timestamp 1676037725
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1676037725
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1676037725
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1676037725
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1676037725
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1676037725
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1676037725
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1676037725
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1676037725
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1676037725
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_9
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1676037725
transform 1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_28
timestamp 1676037725
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_41
timestamp 1676037725
transform 1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_64
timestamp 1676037725
transform 1 0 6992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1676037725
transform 1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1676037725
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_116
timestamp 1676037725
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1676037725
transform 1 0 15364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_194
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1676037725
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_228
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_251
timestamp 1676037725
transform 1 0 24196 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_255
timestamp 1676037725
transform 1 0 24564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_267
timestamp 1676037725
transform 1 0 25668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1676037725
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1676037725
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1676037725
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1676037725
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1676037725
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1676037725
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1676037725
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_517
timestamp 1676037725
transform 1 0 48668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_23
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_34
timestamp 1676037725
transform 1 0 4232 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_42
timestamp 1676037725
transform 1 0 4968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 1676037725
transform 1 0 7452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1676037725
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_102
timestamp 1676037725
transform 1 0 10488 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_143
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1676037725
transform 1 0 14536 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_159
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_185
timestamp 1676037725
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_191
timestamp 1676037725
transform 1 0 18676 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1676037725
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1676037725
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_255
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_267
timestamp 1676037725
transform 1 0 25668 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_279
timestamp 1676037725
transform 1 0 26772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_291
timestamp 1676037725
transform 1 0 27876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1676037725
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1676037725
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1676037725
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1676037725
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1676037725
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1676037725
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1676037725
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1676037725
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1676037725
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1676037725
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1676037725
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1676037725
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1676037725
transform 1 0 3220 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_29
timestamp 1676037725
transform 1 0 3772 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1676037725
transform 1 0 4508 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1676037725
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1676037725
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_60
timestamp 1676037725
transform 1 0 6624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_71
timestamp 1676037725
transform 1 0 7636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1676037725
transform 1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_120
timestamp 1676037725
transform 1 0 12144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_133
timestamp 1676037725
transform 1 0 13340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1676037725
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_174
timestamp 1676037725
transform 1 0 17112 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_190
timestamp 1676037725
transform 1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_231
timestamp 1676037725
transform 1 0 22356 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_262
timestamp 1676037725
transform 1 0 25208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1676037725
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1676037725
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1676037725
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1676037725
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1676037725
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1676037725
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1676037725
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1676037725
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1676037725
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1676037725
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1676037725
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1676037725
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1676037725
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1676037725
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_21
timestamp 1676037725
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_31
timestamp 1676037725
transform 1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_59
timestamp 1676037725
transform 1 0 6532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1676037725
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1676037725
transform 1 0 16744 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_201
timestamp 1676037725
transform 1 0 19596 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_229
timestamp 1676037725
transform 1 0 22172 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_234
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_266
timestamp 1676037725
transform 1 0 25576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_278
timestamp 1676037725
transform 1 0 26680 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_290
timestamp 1676037725
transform 1 0 27784 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1676037725
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1676037725
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1676037725
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1676037725
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1676037725
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1676037725
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1676037725
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1676037725
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1676037725
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1676037725
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1676037725
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1676037725
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1676037725
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_28
timestamp 1676037725
transform 1 0 3680 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_41
timestamp 1676037725
transform 1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_61
timestamp 1676037725
transform 1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1676037725
transform 1 0 7728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_85
timestamp 1676037725
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 1676037725
transform 1 0 11776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1676037725
transform 1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_171
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1676037725
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1676037725
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_227
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1676037725
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1676037725
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 1676037725
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1676037725
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1676037725
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1676037725
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1676037725
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1676037725
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1676037725
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1676037725
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1676037725
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1676037725
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1676037725
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1676037725
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1676037725
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1676037725
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1676037725
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_21
timestamp 1676037725
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1676037725
transform 1 0 4048 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_43
timestamp 1676037725
transform 1 0 5060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1676037725
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_72
timestamp 1676037725
transform 1 0 7728 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1676037725
transform 1 0 9200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1676037725
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_112
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1676037725
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1676037725
transform 1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_191
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_202
timestamp 1676037725
transform 1 0 19688 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_210
timestamp 1676037725
transform 1 0 20424 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_220
timestamp 1676037725
transform 1 0 21344 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_226
timestamp 1676037725
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_264
timestamp 1676037725
transform 1 0 25392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_277
timestamp 1676037725
transform 1 0 26588 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_283
timestamp 1676037725
transform 1 0 27140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_295
timestamp 1676037725
transform 1 0 28244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1676037725
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1676037725
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1676037725
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1676037725
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1676037725
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1676037725
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1676037725
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1676037725
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1676037725
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1676037725
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1676037725
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1676037725
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1676037725
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1676037725
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1676037725
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_25
timestamp 1676037725
transform 1 0 3404 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_29
timestamp 1676037725
transform 1 0 3772 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1676037725
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_63
timestamp 1676037725
transform 1 0 6900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_76
timestamp 1676037725
transform 1 0 8096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1676037725
transform 1 0 8832 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_97
timestamp 1676037725
transform 1 0 10028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1676037725
transform 1 0 13800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1676037725
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_171
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_194
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_211
timestamp 1676037725
transform 1 0 20516 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_247
timestamp 1676037725
transform 1 0 23828 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_253
timestamp 1676037725
transform 1 0 24380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_257
timestamp 1676037725
transform 1 0 24748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_283
timestamp 1676037725
transform 1 0 27140 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_295
timestamp 1676037725
transform 1 0 28244 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_307
timestamp 1676037725
transform 1 0 29348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_319
timestamp 1676037725
transform 1 0 30452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_331
timestamp 1676037725
transform 1 0 31556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1676037725
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1676037725
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1676037725
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1676037725
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1676037725
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1676037725
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1676037725
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1676037725
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_517
timestamp 1676037725
transform 1 0 48668 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp 1676037725
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_66
timestamp 1676037725
transform 1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1676037725
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_91
timestamp 1676037725
transform 1 0 9476 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1676037725
transform 1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1676037725
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_128
timestamp 1676037725
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1676037725
transform 1 0 15272 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_158
timestamp 1676037725
transform 1 0 15640 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_169
timestamp 1676037725
transform 1 0 16652 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1676037725
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_202
timestamp 1676037725
transform 1 0 19688 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1676037725
transform 1 0 20056 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_228
timestamp 1676037725
transform 1 0 22080 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_234
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_237
timestamp 1676037725
transform 1 0 22908 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_255
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_271
timestamp 1676037725
transform 1 0 26036 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1676037725
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1676037725
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1676037725
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1676037725
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1676037725
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1676037725
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1676037725
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1676037725
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1676037725
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1676037725
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1676037725
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_41
timestamp 1676037725
transform 1 0 4876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_63
timestamp 1676037725
transform 1 0 6900 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_76
timestamp 1676037725
transform 1 0 8096 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1676037725
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1676037725
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_138
timestamp 1676037725
transform 1 0 13800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_142
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1676037725
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1676037725
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1676037725
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1676037725
transform 1 0 19504 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1676037725
transform 1 0 19872 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1676037725
transform 1 0 20884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_250
timestamp 1676037725
transform 1 0 24104 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_256
timestamp 1676037725
transform 1 0 24656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_283
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 1676037725
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_290
timestamp 1676037725
transform 1 0 27784 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_302
timestamp 1676037725
transform 1 0 28888 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_314
timestamp 1676037725
transform 1 0 29992 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_326
timestamp 1676037725
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1676037725
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1676037725
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1676037725
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1676037725
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1676037725
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1676037725
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_517
timestamp 1676037725
transform 1 0 48668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1676037725
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_55
timestamp 1676037725
transform 1 0 6164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_59
timestamp 1676037725
transform 1 0 6532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1676037725
transform 1 0 7452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_91
timestamp 1676037725
transform 1 0 9476 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_95
timestamp 1676037725
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1676037725
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_119
timestamp 1676037725
transform 1 0 12052 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1676037725
transform 1 0 12788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_147
timestamp 1676037725
transform 1 0 14628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_160
timestamp 1676037725
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1676037725
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_173
timestamp 1676037725
transform 1 0 17020 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1676037725
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1676037725
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_222
timestamp 1676037725
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_226
timestamp 1676037725
transform 1 0 21896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1676037725
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1676037725
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_271
timestamp 1676037725
transform 1 0 26036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1676037725
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_299
timestamp 1676037725
transform 1 0 28612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1676037725
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1676037725
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1676037725
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1676037725
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1676037725
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1676037725
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1676037725
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1676037725
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1676037725
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1676037725
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1676037725
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_21
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_60
timestamp 1676037725
transform 1 0 6624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1676037725
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_84
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_89
timestamp 1676037725
transform 1 0 9292 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_100
timestamp 1676037725
transform 1 0 10304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1676037725
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1676037725
transform 1 0 12420 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_133
timestamp 1676037725
transform 1 0 13340 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_154
timestamp 1676037725
transform 1 0 15272 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1676037725
transform 1 0 15732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_180
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1676037725
transform 1 0 18032 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_205
timestamp 1676037725
transform 1 0 19964 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1676037725
transform 1 0 20516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_236
timestamp 1676037725
transform 1 0 22816 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_240
timestamp 1676037725
transform 1 0 23184 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_250
timestamp 1676037725
transform 1 0 24104 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1676037725
transform 1 0 24472 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_276
timestamp 1676037725
transform 1 0 26496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1676037725
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_310
timestamp 1676037725
transform 1 0 29624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_314
timestamp 1676037725
transform 1 0 29992 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_326
timestamp 1676037725
transform 1 0 31096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1676037725
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1676037725
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1676037725
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1676037725
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1676037725
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1676037725
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1676037725
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1676037725
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1676037725
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_21
timestamp 1676037725
transform 1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_31
timestamp 1676037725
transform 1 0 3956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_37
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1676037725
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1676037725
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_102
timestamp 1676037725
transform 1 0 10488 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_112
timestamp 1676037725
transform 1 0 11408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_116
timestamp 1676037725
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_147
timestamp 1676037725
transform 1 0 14628 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_158
timestamp 1676037725
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1676037725
transform 1 0 16100 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_185
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_222
timestamp 1676037725
transform 1 0 21528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_255
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1676037725
transform 1 0 26680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1676037725
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_320
timestamp 1676037725
transform 1 0 30544 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1676037725
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1676037725
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1676037725
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1676037725
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1676037725
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1676037725
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1676037725
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1676037725
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1676037725
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1676037725
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1676037725
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1676037725
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1676037725
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1676037725
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_41
timestamp 1676037725
transform 1 0 4876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1676037725
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_75
timestamp 1676037725
transform 1 0 8004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_79
timestamp 1676037725
transform 1 0 8372 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1676037725
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1676037725
transform 1 0 10212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_116
timestamp 1676037725
transform 1 0 11776 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_127
timestamp 1676037725
transform 1 0 12788 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_134
timestamp 1676037725
transform 1 0 13432 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_147
timestamp 1676037725
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_160
timestamp 1676037725
transform 1 0 15824 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_188
timestamp 1676037725
transform 1 0 18400 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_192
timestamp 1676037725
transform 1 0 18768 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_209
timestamp 1676037725
transform 1 0 20332 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_230
timestamp 1676037725
transform 1 0 22264 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_234
timestamp 1676037725
transform 1 0 22632 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1676037725
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_274
timestamp 1676037725
transform 1 0 26312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_286
timestamp 1676037725
transform 1 0 27416 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_292
timestamp 1676037725
transform 1 0 27968 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1676037725
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_326
timestamp 1676037725
transform 1 0 31096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1676037725
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1676037725
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1676037725
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1676037725
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1676037725
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1676037725
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1676037725
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1676037725
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1676037725
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_517
timestamp 1676037725
transform 1 0 48668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_34
timestamp 1676037725
transform 1 0 4232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1676037725
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1676037725
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_99
timestamp 1676037725
transform 1 0 10212 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_104
timestamp 1676037725
transform 1 0 10672 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_110
timestamp 1676037725
transform 1 0 11224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1676037725
transform 1 0 12420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_143
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1676037725
transform 1 0 14812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_173
timestamp 1676037725
transform 1 0 17020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_199
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1676037725
transform 1 0 20608 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_216
timestamp 1676037725
transform 1 0 20976 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_238
timestamp 1676037725
transform 1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_245
timestamp 1676037725
transform 1 0 23644 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_258
timestamp 1676037725
transform 1 0 24840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_262
timestamp 1676037725
transform 1 0 25208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1676037725
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1676037725
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_320
timestamp 1676037725
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_324
timestamp 1676037725
transform 1 0 30912 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_336
timestamp 1676037725
transform 1 0 32016 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_348
timestamp 1676037725
transform 1 0 33120 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1676037725
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1676037725
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1676037725
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1676037725
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1676037725
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1676037725
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1676037725
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1676037725
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1676037725
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1676037725
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1676037725
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1676037725
transform 1 0 8004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_95
timestamp 1676037725
transform 1 0 9844 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_135
timestamp 1676037725
transform 1 0 13524 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_142
timestamp 1676037725
transform 1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_173
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_178
timestamp 1676037725
transform 1 0 17480 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1676037725
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1676037725
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1676037725
transform 1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_240
timestamp 1676037725
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_243
timestamp 1676037725
transform 1 0 23460 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_254
timestamp 1676037725
transform 1 0 24472 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_258
timestamp 1676037725
transform 1 0 24840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_270
timestamp 1676037725
transform 1 0 25944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_274
timestamp 1676037725
transform 1 0 26312 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_283
timestamp 1676037725
transform 1 0 27140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_288
timestamp 1676037725
transform 1 0 27600 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_315
timestamp 1676037725
transform 1 0 30084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_322
timestamp 1676037725
transform 1 0 30728 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1676037725
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1676037725
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1676037725
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1676037725
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1676037725
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1676037725
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1676037725
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1676037725
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_517
timestamp 1676037725
transform 1 0 48668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_35
timestamp 1676037725
transform 1 0 4324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1676037725
transform 1 0 6348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_107
timestamp 1676037725
transform 1 0 10948 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_114
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1676037725
transform 1 0 12604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1676037725
transform 1 0 14352 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_166
timestamp 1676037725
transform 1 0 16376 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1676037725
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_184
timestamp 1676037725
transform 1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_204
timestamp 1676037725
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1676037725
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_236
timestamp 1676037725
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_240
timestamp 1676037725
transform 1 0 23184 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_293
timestamp 1676037725
transform 1 0 28060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_314
timestamp 1676037725
transform 1 0 29992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_320
timestamp 1676037725
transform 1 0 30544 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_331
timestamp 1676037725
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_343
timestamp 1676037725
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1676037725
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1676037725
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1676037725
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1676037725
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1676037725
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1676037725
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1676037725
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1676037725
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1676037725
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1676037725
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1676037725
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1676037725
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_80
timestamp 1676037725
transform 1 0 8464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_86
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_133
timestamp 1676037725
transform 1 0 13340 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1676037725
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_182
timestamp 1676037725
transform 1 0 17848 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_187
timestamp 1676037725
transform 1 0 18308 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1676037725
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_238
timestamp 1676037725
transform 1 0 23000 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_245
timestamp 1676037725
transform 1 0 23644 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_250
timestamp 1676037725
transform 1 0 24104 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_272
timestamp 1676037725
transform 1 0 26128 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1676037725
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 1676037725
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_329
timestamp 1676037725
transform 1 0 31372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1676037725
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_339
timestamp 1676037725
transform 1 0 32292 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_351
timestamp 1676037725
transform 1 0 33396 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_363
timestamp 1676037725
transform 1 0 34500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_375
timestamp 1676037725
transform 1 0 35604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_387
timestamp 1676037725
transform 1 0 36708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1676037725
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1676037725
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1676037725
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1676037725
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_517
timestamp 1676037725
transform 1 0 48668 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_21
timestamp 1676037725
transform 1 0 3036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_45
timestamp 1676037725
transform 1 0 5244 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_103
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_108
timestamp 1676037725
transform 1 0 11040 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_114
timestamp 1676037725
transform 1 0 11592 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_134
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_144
timestamp 1676037725
transform 1 0 14352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1676037725
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_168
timestamp 1676037725
transform 1 0 16560 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1676037725
transform 1 0 17756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_219
timestamp 1676037725
transform 1 0 21252 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_226
timestamp 1676037725
transform 1 0 21896 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1676037725
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_269
timestamp 1676037725
transform 1 0 25852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_291
timestamp 1676037725
transform 1 0 27876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_321
timestamp 1676037725
transform 1 0 30636 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_329
timestamp 1676037725
transform 1 0 31372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_337
timestamp 1676037725
transform 1 0 32108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_344
timestamp 1676037725
transform 1 0 32752 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_348
timestamp 1676037725
transform 1 0 33120 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1676037725
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1676037725
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1676037725
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1676037725
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1676037725
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1676037725
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1676037725
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1676037725
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1676037725
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_61
timestamp 1676037725
transform 1 0 6716 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_67
timestamp 1676037725
transform 1 0 7268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_91
timestamp 1676037725
transform 1 0 9476 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_104
timestamp 1676037725
transform 1 0 10672 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_129
timestamp 1676037725
transform 1 0 12972 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_150
timestamp 1676037725
transform 1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_155
timestamp 1676037725
transform 1 0 15364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1676037725
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_211
timestamp 1676037725
transform 1 0 20516 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_217
timestamp 1676037725
transform 1 0 21068 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_275
timestamp 1676037725
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_293
timestamp 1676037725
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_317
timestamp 1676037725
transform 1 0 30268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_330
timestamp 1676037725
transform 1 0 31464 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_343
timestamp 1676037725
transform 1 0 32660 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_355
timestamp 1676037725
transform 1 0 33764 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_367
timestamp 1676037725
transform 1 0 34868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_379
timestamp 1676037725
transform 1 0 35972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1676037725
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1676037725
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1676037725
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1676037725
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1676037725
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_507
timestamp 1676037725
transform 1 0 47748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_21
timestamp 1676037725
transform 1 0 3036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_47
timestamp 1676037725
transform 1 0 5428 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_52
timestamp 1676037725
transform 1 0 5888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_57
timestamp 1676037725
transform 1 0 6348 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_61
timestamp 1676037725
transform 1 0 6716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_78
timestamp 1676037725
transform 1 0 8280 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_87
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_98
timestamp 1676037725
transform 1 0 10120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_147
timestamp 1676037725
transform 1 0 14628 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_151
timestamp 1676037725
transform 1 0 14996 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_169
timestamp 1676037725
transform 1 0 16652 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_173
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1676037725
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_207
timestamp 1676037725
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_225
timestamp 1676037725
transform 1 0 21804 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_229
timestamp 1676037725
transform 1 0 22172 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_232
timestamp 1676037725
transform 1 0 22448 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 1676037725
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1676037725
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1676037725
transform 1 0 28244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_302
timestamp 1676037725
transform 1 0 28888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_313
timestamp 1676037725
transform 1 0 29900 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_324
timestamp 1676037725
transform 1 0 30912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_332
timestamp 1676037725
transform 1 0 31648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_340
timestamp 1676037725
transform 1 0 32384 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_352
timestamp 1676037725
transform 1 0 33488 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1676037725
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1676037725
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1676037725
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1676037725
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1676037725
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1676037725
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1676037725
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_513
timestamp 1676037725
transform 1 0 48300 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_517
timestamp 1676037725
transform 1 0 48668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1676037725
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1676037725
transform 1 0 6532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_70
timestamp 1676037725
transform 1 0 7544 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_90
timestamp 1676037725
transform 1 0 9384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_119
timestamp 1676037725
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_143
timestamp 1676037725
transform 1 0 14260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_148
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1676037725
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_230
timestamp 1676037725
transform 1 0 22264 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_235
timestamp 1676037725
transform 1 0 22724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1676037725
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_272
timestamp 1676037725
transform 1 0 26128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1676037725
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_316
timestamp 1676037725
transform 1 0 30176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_329
timestamp 1676037725
transform 1 0 31372 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1676037725
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_343
timestamp 1676037725
transform 1 0 32660 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_351
timestamp 1676037725
transform 1 0 33396 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_363
timestamp 1676037725
transform 1 0 34500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_371
timestamp 1676037725
transform 1 0 35236 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_374
timestamp 1676037725
transform 1 0 35512 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_386
timestamp 1676037725
transform 1 0 36616 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_397
timestamp 1676037725
transform 1 0 37628 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_419
timestamp 1676037725
transform 1 0 39652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_423
timestamp 1676037725
transform 1 0 40020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_435
timestamp 1676037725
transform 1 0 41124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1676037725
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1676037725
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_511
timestamp 1676037725
transform 1 0 48116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_87
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_133
timestamp 1676037725
transform 1 0 13340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_147
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_152
timestamp 1676037725
transform 1 0 15088 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1676037725
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1676037725
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1676037725
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_277
timestamp 1676037725
transform 1 0 26588 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_281
timestamp 1676037725
transform 1 0 26956 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_304
timestamp 1676037725
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_331
timestamp 1676037725
transform 1 0 31556 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_337
timestamp 1676037725
transform 1 0 32108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_343
timestamp 1676037725
transform 1 0 32660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_351
timestamp 1676037725
transform 1 0 33396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_359
timestamp 1676037725
transform 1 0 34132 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_370
timestamp 1676037725
transform 1 0 35144 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_384
timestamp 1676037725
transform 1 0 36432 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_392
timestamp 1676037725
transform 1 0 37168 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_395
timestamp 1676037725
transform 1 0 37444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_407
timestamp 1676037725
transform 1 0 38548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_433
timestamp 1676037725
transform 1 0 40940 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_455
timestamp 1676037725
transform 1 0 42964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_467
timestamp 1676037725
transform 1 0 44068 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1676037725
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_507
timestamp 1676037725
transform 1 0 47748 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_513
timestamp 1676037725
transform 1 0 48300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_8
timestamp 1676037725
transform 1 0 1840 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1676037725
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1676037725
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_115
timestamp 1676037725
transform 1 0 11684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1676037725
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_187
timestamp 1676037725
transform 1 0 18308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_211
timestamp 1676037725
transform 1 0 20516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_219
timestamp 1676037725
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1676037725
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1676037725
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_303
timestamp 1676037725
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_310
timestamp 1676037725
transform 1 0 29624 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_318
timestamp 1676037725
transform 1 0 30360 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_326
timestamp 1676037725
transform 1 0 31096 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_331
timestamp 1676037725
transform 1 0 31556 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_342
timestamp 1676037725
transform 1 0 32568 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_349
timestamp 1676037725
transform 1 0 33212 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_353
timestamp 1676037725
transform 1 0 33580 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_360
timestamp 1676037725
transform 1 0 34224 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_368
timestamp 1676037725
transform 1 0 34960 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_376
timestamp 1676037725
transform 1 0 35696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_383
timestamp 1676037725
transform 1 0 36340 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1676037725
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_395
timestamp 1676037725
transform 1 0 37444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_401
timestamp 1676037725
transform 1 0 37996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_409
timestamp 1676037725
transform 1 0 38732 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_413
timestamp 1676037725
transform 1 0 39100 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_423
timestamp 1676037725
transform 1 0 40020 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_428
timestamp 1676037725
transform 1 0 40480 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_433
timestamp 1676037725
transform 1 0 40940 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_440
timestamp 1676037725
transform 1 0 41584 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1676037725
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_459
timestamp 1676037725
transform 1 0 43332 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_471
timestamp 1676037725
transform 1 0 44436 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_479
timestamp 1676037725
transform 1 0 45172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_487
timestamp 1676037725
transform 1 0 45908 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_493
timestamp 1676037725
transform 1 0 46460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_500
timestamp 1676037725
transform 1 0 47104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_507
timestamp 1676037725
transform 1 0 47748 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_513
timestamp 1676037725
transform 1 0 48300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_525
timestamp 1676037725
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_8
timestamp 1676037725
transform 1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1676037725
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_191
timestamp 1676037725
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1676037725
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1676037725
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1676037725
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_299
timestamp 1676037725
transform 1 0 28612 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1676037725
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_325
timestamp 1676037725
transform 1 0 31004 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_331
timestamp 1676037725
transform 1 0 31556 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_335
timestamp 1676037725
transform 1 0 31924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1676037725
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_342
timestamp 1676037725
transform 1 0 32568 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_346
timestamp 1676037725
transform 1 0 32936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_353
timestamp 1676037725
transform 1 0 33580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1676037725
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_371
timestamp 1676037725
transform 1 0 35236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_379
timestamp 1676037725
transform 1 0 35972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_386
timestamp 1676037725
transform 1 0 36616 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1676037725
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_398
timestamp 1676037725
transform 1 0 37720 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_402
timestamp 1676037725
transform 1 0 38088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_409
timestamp 1676037725
transform 1 0 38732 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_417
timestamp 1676037725
transform 1 0 39468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_433
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_437
timestamp 1676037725
transform 1 0 41308 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_446
timestamp 1676037725
transform 1 0 42136 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_451
timestamp 1676037725
transform 1 0 42596 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_463
timestamp 1676037725
transform 1 0 43700 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_467
timestamp 1676037725
transform 1 0 44068 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_471
timestamp 1676037725
transform 1 0 44436 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_483
timestamp 1676037725
transform 1 0 45540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_491
timestamp 1676037725
transform 1 0 46276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_499
timestamp 1676037725
transform 1 0 47012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1676037725
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1676037725
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_511
timestamp 1676037725
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_515
timestamp 1676037725
transform 1 0 48484 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_524
timestamp 1676037725
transform 1 0 49312 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42596 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold2
timestamp 1676037725
transform 1 0 41124 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1676037725
transform 1 0 41400 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1676037725
transform 1 0 43332 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold5 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1676037725
transform 1 0 48576 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1676037725
transform 1 0 43884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1676037725
transform 1 0 2944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1676037725
transform 1 0 6532 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1676037725
transform 1 0 48668 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1676037725
transform 1 0 48668 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1676037725
transform 1 0 1840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1676037725
transform 1 0 2852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 48392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 2944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1676037725
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 2852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1676037725
transform 1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1676037725
transform 1 0 29992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 31280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 35512 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 32292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 36064 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1676037725
transform 1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1676037725
transform 1 0 33948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 34868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 28612 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 35604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 36340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 36708 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 37444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 37720 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1676037725
transform 1 0 38364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1676037725
transform 1 0 39100 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 40020 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 40664 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1676037725
transform 1 0 41308 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1676037725
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 28980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 28336 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 29348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1676037725
transform 1 0 31280 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 33488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1676037725
transform 1 0 36064 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1676037725
transform 1 0 44160 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1676037725
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 46644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1676037725
transform 1 0 46736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1676037725
transform 1 0 47748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1676037725
transform 1 0 47932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1676037725
transform 1 0 44804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 45540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 49036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 49036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1676037725
transform 1 0 48300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1676037725
transform 1 0 47932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 3404 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 3404 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 3404 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 3956 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 6532 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 3404 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 10488 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 11960 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 12328 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 15272 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 14904 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 6808 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 7912 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 9476 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 12144 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18676 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21160 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18676 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20056 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24288 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25852 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26036 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25760 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27232 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28428 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28244 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27048 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24656 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37812 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27784 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 24840 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24840 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22356 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20884 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20240 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23000 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17480 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16008 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14720 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14628 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12052 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11224 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11500 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 4600 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7636 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9292 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11500 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12420 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13064 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18124 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30728 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27784 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_1.mux_l1_in_1__194
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17204 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_3.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_5.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11224 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_7.mux_l1_in_1__162
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18492 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_9.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6808 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25760 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_11.mux_l2_in_0__195
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_13.mux_l2_in_0__196
timestamp 1676037725
transform 1 0 36156 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14536 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_15.mux_l2_in_0__197
timestamp 1676037725
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28336 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25760 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15732 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_17.mux_l2_in_0__198
timestamp 1676037725
transform 1 0 17480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_19.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 21252 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_29.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 23368 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27232 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_31.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_33.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 22448 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30544 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_35.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 24196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30084 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_45.mux_l2_in_0__157
timestamp 1676037725
transform 1 0 27968 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25576 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30636 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_47.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 26404 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30544 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_49.mux_l2_in_0__159
timestamp 1676037725
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30912 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_51.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_0.mux_l2_in_1__164
timestamp 1676037725
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23644 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23368 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25760 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_2.mux_l2_in_1__170
timestamp 1676037725
transform 1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19044 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23184 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22172 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_4.mux_l2_in_1__181
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12144 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_6.mux_l2_in_1__188
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19688 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_8.mux_l2_in_1__189
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17204 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23368 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_10.mux_l2_in_1__165
timestamp 1676037725
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_12.mux_l1_in_1__166
timestamp 1676037725
transform 1 0 13616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10120 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_14.mux_l1_in_1__167
timestamp 1676037725
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10120 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_16.mux_l1_in_1__168
timestamp 1676037725
transform 1 0 11868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13156 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_18.mux_l1_in_1__169
timestamp 1676037725
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15824 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_20.mux_l2_in_0__171
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14352 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_22.mux_l2_in_0__172
timestamp 1676037725
transform 1 0 15364 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_24.mux_l2_in_0__173
timestamp 1676037725
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14444 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_26.mux_l2_in_0__174
timestamp 1676037725
transform 1 0 6716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10304 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_28.mux_l2_in_0__175
timestamp 1676037725
transform 1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11316 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_30.mux_l2_in_0__176
timestamp 1676037725
transform 1 0 6624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12052 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11960 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_32.mux_l2_in_0__177
timestamp 1676037725
transform 1 0 9384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32476 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_34.mux_l2_in_0__178
timestamp 1676037725
transform 1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 30452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11592 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9292 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_36.mux_l2_in_0__179
timestamp 1676037725
transform 1 0 3404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 7268 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 4140 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_38.mux_l2_in_0__180
timestamp 1676037725
transform 1 0 4692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 8004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 6716 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_40.mux_l2_in_0__182
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_42.mux_l2_in_0__183
timestamp 1676037725
transform 1 0 32936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17848 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_44.mux_l1_in_1__184
timestamp 1676037725
transform 1 0 4692 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32292 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_46.mux_l1_in_1__185
timestamp 1676037725
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32568 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_48.mux_l1_in_1__186
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27600 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_50.mux_l1_in_1__187
timestamp 1676037725
transform 1 0 10212 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 66 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 67 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 68 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 69 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 70 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 71 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 72 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 73 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 74 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 75 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 76 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 77 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 78 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 79 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 80 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 81 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 82 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 83 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 84 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 85 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 86 nsew signal input
flabel metal2 s 40866 26200 40922 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 87 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 88 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 89 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 90 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 91 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 92 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 93 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 94 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 95 nsew signal input
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 96 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 97 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 98 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 99 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 100 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 101 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 102 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 103 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 104 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 105 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 106 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 107 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 108 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 109 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 110 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 111 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 112 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 113 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 114 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 115 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 116 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 117 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 41510 26200 41566 27000 0 FreeSans 224 90 0 0 prog_reset
port 140 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 reset
port 141 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 test_enable
port 142 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 143 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 144 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 145 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 146 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 147 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 148 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 149 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 150 nsew signal input
flabel metal3 s 50200 21904 51000 22024 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 151 nsew signal input
flabel metal3 s 50200 22856 51000 22976 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 152 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 50200 24760 51000 24880 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 154 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 155 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 156 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 158 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal2 17526 6188 17526 6188 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 15686 6222 15686 6222 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 14812 5746 14812 5746 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal2 13662 8738 13662 8738 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20838 17714 20838 17714 0 cbx_8__0_.cbx_8__0_.ccff_head
rlabel metal1 9798 10166 9798 10166 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 14582 16116 14582 16116 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 10948 13838 10948 13838 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal2 8510 9180 8510 9180 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 5704 12138 5704 12138 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal1 10948 14450 10948 14450 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 5980 12750 5980 12750 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 5520 11662 5520 11662 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 8740 11526 8740 11526 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal1 6256 16014 6256 16014 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal2 13662 15708 13662 15708 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 10994 13328 10994 13328 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal2 5934 17289 5934 17289 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 7544 17102 7544 17102 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 8602 18768 8602 18768 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal1 8050 14450 8050 14450 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8786 9146 8786 9146 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 14306 7344 14306 7344 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 8234 14382 8234 14382 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 8878 14977 8878 14977 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10442 15130 10442 15130 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11592 14042 11592 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8096 11186 8096 11186 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9062 14790 9062 14790 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8970 8058 8970 8058 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 8234 9282 8234 9282 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10718 9622 10718 9622 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 4416 14042 4416 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 4876 11866 4876 11866 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 10120 7378 10120 7378 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 2622 18360 2622 18360 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6808 15538 6808 15538 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7360 15402 7360 15402 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8970 12954 8970 12954 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 5198 13974 5198 13974 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6026 14042 6026 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 6302 11798 6302 11798 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 5382 12614 5382 12614 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 4922 11730 4922 11730 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 5428 15538 5428 15538 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10120 13158 10120 13158 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 12581 7378 12581 7378 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 4784 15402 4784 15402 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6348 13906 6348 13906 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7314 14416 7314 14416 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10534 14450 10534 14450 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 8602 14501 8602 14501 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6946 14008 6946 14008 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 10902 12886 10902 12886 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 13662 14076 13662 14076 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8694 14042 8694 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 8878 17578 8878 17578 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10488 17850 10488 17850 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 4968 13124 4968 13124 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 7682 17646 7682 17646 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6302 17034 6302 17034 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7544 15674 7544 15674 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10396 14382 10396 14382 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7544 22610 7544 22610 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6992 22610 6992 22610 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9476 14586 9476 14586 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 14398 19040 14398 19040 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 5888 19482 5888 19482 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 17434 4284 17434 4284 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal2 17710 4114 17710 4114 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal2 20562 4012 20562 4012 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 26795 4794 26795 4794 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 19964 5882 19964 5882 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 15686 5134 15686 5134 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 18124 3026 18124 3026 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 25047 5338 25047 5338 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 25806 7514 25806 7514 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 16468 5678 16468 5678 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 17066 4284 17066 4284 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal2 25990 4760 25990 4760 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 15456 7854 15456 7854 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 15226 6052 15226 6052 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 23828 5746 23828 5746 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 1656 4114 1656 4114 0 ccff_head
rlabel metal1 48622 23086 48622 23086 0 ccff_head_1
rlabel metal2 49174 21233 49174 21233 0 ccff_tail
rlabel metal2 2254 24218 2254 24218 0 ccff_tail_0
rlabel metal3 1786 1564 1786 1564 0 chanx_left_in[0]
rlabel metal1 1472 5678 1472 5678 0 chanx_left_in[10]
rlabel metal1 1472 6222 1472 6222 0 chanx_left_in[11]
rlabel metal3 1004 6460 1004 6460 0 chanx_left_in[12]
rlabel metal1 3358 7378 3358 7378 0 chanx_left_in[13]
rlabel metal1 2990 6290 2990 6290 0 chanx_left_in[14]
rlabel metal3 1004 7684 1004 7684 0 chanx_left_in[15]
rlabel via1 2622 6749 2622 6749 0 chanx_left_in[16]
rlabel metal1 2990 7854 2990 7854 0 chanx_left_in[17]
rlabel metal2 1794 7837 1794 7837 0 chanx_left_in[18]
rlabel metal1 2530 7378 2530 7378 0 chanx_left_in[19]
rlabel metal1 3082 2380 3082 2380 0 chanx_left_in[1]
rlabel metal2 1610 9367 1610 9367 0 chanx_left_in[20]
rlabel metal1 2990 8942 2990 8942 0 chanx_left_in[21]
rlabel metal2 2622 8687 2622 8687 0 chanx_left_in[22]
rlabel metal1 1656 8466 1656 8466 0 chanx_left_in[23]
rlabel metal3 1717 11356 1717 11356 0 chanx_left_in[24]
rlabel metal1 1518 10098 1518 10098 0 chanx_left_in[25]
rlabel metal1 1564 12206 1564 12206 0 chanx_left_in[26]
rlabel metal3 1372 12580 1372 12580 0 chanx_left_in[27]
rlabel metal1 1794 7956 1794 7956 0 chanx_left_in[28]
rlabel metal3 958 13396 958 13396 0 chanx_left_in[29]
rlabel metal1 2714 2482 2714 2482 0 chanx_left_in[2]
rlabel metal1 3174 2550 3174 2550 0 chanx_left_in[3]
rlabel metal1 1472 3502 1472 3502 0 chanx_left_in[4]
rlabel metal1 2990 4590 2990 4590 0 chanx_left_in[5]
rlabel metal1 4140 3502 4140 3502 0 chanx_left_in[6]
rlabel metal1 4232 4114 4232 4114 0 chanx_left_in[7]
rlabel metal1 1472 4658 1472 4658 0 chanx_left_in[8]
rlabel metal1 1472 5202 1472 5202 0 chanx_left_in[9]
rlabel metal3 1372 13804 1372 13804 0 chanx_left_out[0]
rlabel metal2 2806 18275 2806 18275 0 chanx_left_out[10]
rlabel metal2 2898 18819 2898 18819 0 chanx_left_out[11]
rlabel metal2 3358 19295 3358 19295 0 chanx_left_out[12]
rlabel metal3 1717 19108 1717 19108 0 chanx_left_out[13]
rlabel metal2 2806 20179 2806 20179 0 chanx_left_out[14]
rlabel metal3 1372 19924 1372 19924 0 chanx_left_out[15]
rlabel via2 3910 20349 3910 20349 0 chanx_left_out[16]
rlabel metal3 1004 20740 1004 20740 0 chanx_left_out[17]
rlabel metal2 2852 21148 2852 21148 0 chanx_left_out[18]
rlabel metal3 1832 21556 1832 21556 0 chanx_left_out[19]
rlabel metal3 1004 14212 1004 14212 0 chanx_left_out[1]
rlabel metal3 2660 21964 2660 21964 0 chanx_left_out[20]
rlabel metal3 1418 22372 1418 22372 0 chanx_left_out[21]
rlabel metal3 2844 22780 2844 22780 0 chanx_left_out[22]
rlabel metal3 2200 23188 2200 23188 0 chanx_left_out[23]
rlabel metal1 8786 20910 8786 20910 0 chanx_left_out[24]
rlabel metal2 4324 21148 4324 21148 0 chanx_left_out[25]
rlabel metal2 4554 19353 4554 19353 0 chanx_left_out[26]
rlabel metal2 3082 24735 3082 24735 0 chanx_left_out[27]
rlabel metal2 7544 21828 7544 21828 0 chanx_left_out[28]
rlabel metal1 4094 20502 4094 20502 0 chanx_left_out[29]
rlabel metal3 1004 14620 1004 14620 0 chanx_left_out[2]
rlabel metal3 1004 15028 1004 15028 0 chanx_left_out[3]
rlabel metal3 1004 15436 1004 15436 0 chanx_left_out[4]
rlabel metal3 1004 15844 1004 15844 0 chanx_left_out[5]
rlabel metal3 1004 16252 1004 16252 0 chanx_left_out[6]
rlabel metal3 1004 16660 1004 16660 0 chanx_left_out[7]
rlabel metal3 958 17068 958 17068 0 chanx_left_out[8]
rlabel metal3 1372 17476 1372 17476 0 chanx_left_out[9]
rlabel metal2 5198 8704 5198 8704 0 chany_top_in[0]
rlabel metal1 28842 23086 28842 23086 0 chany_top_in[10]
rlabel metal1 29532 24242 29532 24242 0 chany_top_in[11]
rlabel metal2 33442 21182 33442 21182 0 chany_top_in[12]
rlabel metal1 32614 21454 32614 21454 0 chany_top_in[13]
rlabel metal1 34362 22406 34362 22406 0 chany_top_in[14]
rlabel metal1 33534 22066 33534 22066 0 chany_top_in[15]
rlabel metal2 36294 24174 36294 24174 0 chany_top_in[16]
rlabel metal2 33350 24429 33350 24429 0 chany_top_in[17]
rlabel metal2 34086 25245 34086 25245 0 chany_top_in[18]
rlabel metal1 34776 24106 34776 24106 0 chany_top_in[19]
rlabel metal1 30429 21998 30429 21998 0 chany_top_in[1]
rlabel metal1 35466 24106 35466 24106 0 chany_top_in[20]
rlabel metal1 36248 24174 36248 24174 0 chany_top_in[21]
rlabel metal1 36662 23698 36662 23698 0 chany_top_in[22]
rlabel metal1 37490 24174 37490 24174 0 chany_top_in[23]
rlabel metal1 37812 23698 37812 23698 0 chany_top_in[24]
rlabel metal2 38502 25245 38502 25245 0 chany_top_in[25]
rlabel metal2 39238 25245 39238 25245 0 chany_top_in[26]
rlabel metal1 39836 24242 39836 24242 0 chany_top_in[27]
rlabel metal2 40342 25075 40342 25075 0 chany_top_in[28]
rlabel metal1 41676 23698 41676 23698 0 chany_top_in[29]
rlabel metal2 19274 22253 19274 22253 0 chany_top_in[2]
rlabel metal3 18676 23120 18676 23120 0 chany_top_in[3]
rlabel metal3 22724 23528 22724 23528 0 chany_top_in[4]
rlabel metal3 18492 22984 18492 22984 0 chany_top_in[5]
rlabel metal2 33074 23018 33074 23018 0 chany_top_in[6]
rlabel metal1 28520 24174 28520 24174 0 chany_top_in[7]
rlabel metal2 29578 24208 29578 24208 0 chany_top_in[8]
rlabel metal2 28750 24174 28750 24174 0 chany_top_in[9]
rlabel metal1 3634 23154 3634 23154 0 chany_top_out[0]
rlabel metal1 8740 24242 8740 24242 0 chany_top_out[10]
rlabel metal1 9568 23766 9568 23766 0 chany_top_out[11]
rlabel metal2 10718 24497 10718 24497 0 chany_top_out[12]
rlabel metal2 11270 24184 11270 24184 0 chany_top_out[13]
rlabel metal2 12558 21862 12558 21862 0 chany_top_out[14]
rlabel metal2 12558 25034 12558 25034 0 chany_top_out[15]
rlabel metal2 13301 26316 13301 26316 0 chany_top_out[16]
rlabel metal2 13846 25204 13846 25204 0 chany_top_out[17]
rlabel metal1 13570 24276 13570 24276 0 chany_top_out[18]
rlabel metal1 15410 22066 15410 22066 0 chany_top_out[19]
rlabel metal1 3404 24242 3404 24242 0 chany_top_out[1]
rlabel metal1 15042 23766 15042 23766 0 chany_top_out[20]
rlabel metal2 16146 24497 16146 24497 0 chany_top_out[21]
rlabel metal2 17211 26316 17211 26316 0 chany_top_out[22]
rlabel metal1 16974 23154 16974 23154 0 chany_top_out[23]
rlabel metal1 17250 23766 17250 23766 0 chany_top_out[24]
rlabel metal1 16192 24242 16192 24242 0 chany_top_out[25]
rlabel metal2 17894 23460 17894 23460 0 chany_top_out[26]
rlabel metal1 20792 21930 20792 21930 0 chany_top_out[27]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[28]
rlabel metal2 21574 25272 21574 25272 0 chany_top_out[29]
rlabel metal1 4094 23766 4094 23766 0 chany_top_out[2]
rlabel metal2 5106 24429 5106 24429 0 chany_top_out[3]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[4]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[5]
rlabel metal1 7360 22678 7360 22678 0 chany_top_out[6]
rlabel metal1 6348 24242 6348 24242 0 chany_top_out[7]
rlabel metal2 7866 24735 7866 24735 0 chany_top_out[8]
rlabel metal2 8694 24422 8694 24422 0 chany_top_out[9]
rlabel metal1 20930 18666 20930 18666 0 clknet_0_prog_clk
rlabel metal1 8004 9486 8004 9486 0 clknet_4_0_0_prog_clk
rlabel metal1 26496 13226 26496 13226 0 clknet_4_10_0_prog_clk
rlabel metal2 22034 16320 22034 16320 0 clknet_4_11_0_prog_clk
rlabel metal2 16330 18496 16330 18496 0 clknet_4_12_0_prog_clk
rlabel metal1 19734 20502 19734 20502 0 clknet_4_13_0_prog_clk
rlabel metal1 27968 18258 27968 18258 0 clknet_4_14_0_prog_clk
rlabel metal2 21942 22236 21942 22236 0 clknet_4_15_0_prog_clk
rlabel metal2 9338 13056 9338 13056 0 clknet_4_1_0_prog_clk
rlabel metal1 14536 10030 14536 10030 0 clknet_4_2_0_prog_clk
rlabel metal2 14306 13090 14306 13090 0 clknet_4_3_0_prog_clk
rlabel metal1 4554 17646 4554 17646 0 clknet_4_4_0_prog_clk
rlabel metal1 9430 20298 9430 20298 0 clknet_4_5_0_prog_clk
rlabel metal2 14582 19652 14582 19652 0 clknet_4_6_0_prog_clk
rlabel metal1 12788 21522 12788 21522 0 clknet_4_7_0_prog_clk
rlabel metal2 16882 7616 16882 7616 0 clknet_4_8_0_prog_clk
rlabel metal1 19964 12750 19964 12750 0 clknet_4_9_0_prog_clk
rlabel metal2 4094 1622 4094 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 6762 1622 6762 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 9430 1622 9430 1622 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 12098 1622 12098 1622 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 25576 2414 25576 2414 0 gfpga_pad_io_soc_in[0]
rlabel metal2 28382 1581 28382 1581 0 gfpga_pad_io_soc_in[1]
rlabel metal1 30912 2414 30912 2414 0 gfpga_pad_io_soc_in[2]
rlabel metal1 33580 2414 33580 2414 0 gfpga_pad_io_soc_in[3]
rlabel metal2 14766 1622 14766 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 17434 1622 17434 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 20102 959 20102 959 0 gfpga_pad_io_soc_out[2]
rlabel metal2 22770 1622 22770 1622 0 gfpga_pad_io_soc_out[3]
rlabel metal2 36110 1588 36110 1588 0 isol_n
rlabel metal1 6578 2992 6578 2992 0 net1
rlabel metal2 2300 12716 2300 12716 0 net10
rlabel metal1 5888 17170 5888 17170 0 net100
rlabel metal2 4002 16388 4002 16388 0 net101
rlabel metal2 19320 19380 19320 19380 0 net102
rlabel metal1 8648 19346 8648 19346 0 net103
rlabel metal2 3542 15606 3542 15606 0 net104
rlabel metal1 5106 14314 5106 14314 0 net105
rlabel metal1 1794 15028 1794 15028 0 net106
rlabel metal2 3450 14756 3450 14756 0 net107
rlabel metal1 2277 16082 2277 16082 0 net108
rlabel metal1 2277 16558 2277 16558 0 net109
rlabel metal1 11684 16626 11684 16626 0 net11
rlabel metal2 1794 16966 1794 16966 0 net110
rlabel metal1 1794 17680 1794 17680 0 net111
rlabel metal1 1794 18292 1794 18292 0 net112
rlabel metal1 2254 12682 2254 12682 0 net113
rlabel metal2 8372 16524 8372 16524 0 net114
rlabel metal3 7429 11084 7429 11084 0 net115
rlabel metal2 33626 24684 33626 24684 0 net116
rlabel metal2 35650 24616 35650 24616 0 net117
rlabel metal2 33718 24480 33718 24480 0 net118
rlabel via2 17158 16235 17158 16235 0 net119
rlabel metal1 1610 6664 1610 6664 0 net12
rlabel metal2 12880 22542 12880 22542 0 net120
rlabel metal1 27140 21522 27140 21522 0 net121
rlabel metal1 12696 24174 12696 24174 0 net122
rlabel metal2 15226 21556 15226 21556 0 net123
rlabel metal1 2346 24174 2346 24174 0 net124
rlabel metal2 13524 21420 13524 21420 0 net125
rlabel metal2 15042 23800 15042 23800 0 net126
rlabel metal2 14674 21284 14674 21284 0 net127
rlabel metal2 15502 24072 15502 24072 0 net128
rlabel metal3 18032 17884 18032 17884 0 net129
rlabel metal2 2254 7667 2254 7667 0 net13
rlabel metal1 19688 17714 19688 17714 0 net130
rlabel metal2 16882 23443 16882 23443 0 net131
rlabel metal1 19918 24038 19918 24038 0 net132
rlabel metal1 19274 20026 19274 20026 0 net133
rlabel metal1 21114 24174 21114 24174 0 net134
rlabel metal1 2760 23698 2760 23698 0 net135
rlabel metal2 16146 21386 16146 21386 0 net136
rlabel metal2 21206 24225 21206 24225 0 net137
rlabel metal1 1564 22542 1564 22542 0 net138
rlabel via3 6923 20740 6923 20740 0 net139
rlabel metal1 5336 2618 5336 2618 0 net14
rlabel metal2 1518 23195 1518 23195 0 net140
rlabel metal3 7153 20740 7153 20740 0 net141
rlabel metal1 7636 8262 7636 8262 0 net142
rlabel metal1 4600 2414 4600 2414 0 net143
rlabel metal1 7682 2414 7682 2414 0 net144
rlabel metal1 9706 2414 9706 2414 0 net145
rlabel metal1 12420 2414 12420 2414 0 net146
rlabel metal2 15042 3162 15042 3162 0 net147
rlabel metal1 17204 2822 17204 2822 0 net148
rlabel metal1 19136 2822 19136 2822 0 net149
rlabel metal1 4646 20842 4646 20842 0 net15
rlabel metal1 22356 2414 22356 2414 0 net150
rlabel metal1 21850 21522 21850 21522 0 net151
rlabel metal1 22954 20570 22954 20570 0 net152
rlabel metal1 19136 19754 19136 19754 0 net153
rlabel metal1 23828 21930 23828 21930 0 net154
rlabel metal1 23092 22678 23092 22678 0 net155
rlabel metal1 24610 23834 24610 23834 0 net156
rlabel metal2 25990 21760 25990 21760 0 net157
rlabel metal1 26358 19482 26358 19482 0 net158
rlabel metal1 28658 18394 28658 18394 0 net159
rlabel metal1 6256 21590 6256 21590 0 net16
rlabel metal1 16054 20366 16054 20366 0 net160
rlabel metal1 20240 17646 20240 17646 0 net161
rlabel metal1 24150 18802 24150 18802 0 net162
rlabel metal1 12512 20366 12512 20366 0 net163
rlabel metal2 20470 16796 20470 16796 0 net164
rlabel metal1 14122 8874 14122 8874 0 net165
rlabel metal1 14168 8466 14168 8466 0 net166
rlabel metal1 10580 6834 10580 6834 0 net167
rlabel metal1 11454 7514 11454 7514 0 net168
rlabel metal2 13570 12002 13570 12002 0 net169
rlabel metal1 5934 18258 5934 18258 0 net17
rlabel metal1 13432 7514 13432 7514 0 net170
rlabel metal1 17020 16626 17020 16626 0 net171
rlabel metal2 15410 17034 15410 17034 0 net172
rlabel metal2 14858 15572 14858 15572 0 net173
rlabel metal1 8234 11866 8234 11866 0 net174
rlabel metal2 9430 10030 9430 10030 0 net175
rlabel metal1 9522 15436 9522 15436 0 net176
rlabel metal2 11454 10506 11454 10506 0 net177
rlabel metal1 20102 14790 20102 14790 0 net178
rlabel metal1 16146 15640 16146 15640 0 net179
rlabel metal1 13524 17238 13524 17238 0 net18
rlabel metal2 4646 10115 4646 10115 0 net180
rlabel metal1 12420 8602 12420 8602 0 net181
rlabel metal1 5566 9622 5566 9622 0 net182
rlabel metal2 15916 18564 15916 18564 0 net183
rlabel metal1 9660 21318 9660 21318 0 net184
rlabel metal1 10534 18258 10534 18258 0 net185
rlabel metal1 14030 17170 14030 17170 0 net186
rlabel metal2 12834 16082 12834 16082 0 net187
rlabel metal1 13570 12138 13570 12138 0 net188
rlabel metal1 16146 8602 16146 8602 0 net189
rlabel metal1 13110 16626 13110 16626 0 net19
rlabel metal1 7452 10778 7452 10778 0 net190
rlabel metal1 5750 10098 5750 10098 0 net191
rlabel metal2 16514 14756 16514 14756 0 net192
rlabel metal2 13708 12886 13708 12886 0 net193
rlabel metal1 27922 16558 27922 16558 0 net194
rlabel metal1 32292 23630 32292 23630 0 net195
rlabel via2 15962 21573 15962 21573 0 net196
rlabel metal1 18676 16422 18676 16422 0 net197
rlabel metal1 17112 18802 17112 18802 0 net198
rlabel metal2 43378 23290 43378 23290 0 net199
rlabel metal2 44758 22236 44758 22236 0 net2
rlabel metal1 14352 18870 14352 18870 0 net20
rlabel metal1 31924 11322 31924 11322 0 net200
rlabel metal1 42366 23698 42366 23698 0 net201
rlabel metal1 44206 23290 44206 23290 0 net202
rlabel metal2 41446 23324 41446 23324 0 net203
rlabel metal2 48714 23868 48714 23868 0 net204
rlabel metal1 41354 22542 41354 22542 0 net205
rlabel metal1 3128 3026 3128 3026 0 net206
rlabel metal1 8142 2958 8142 2958 0 net207
rlabel metal1 48990 23290 48990 23290 0 net208
rlabel metal1 48668 21998 48668 21998 0 net209
rlabel metal1 6440 16626 6440 16626 0 net21
rlabel metal1 2760 4114 2760 4114 0 net210
rlabel metal1 3864 3026 3864 3026 0 net211
rlabel metal1 1840 10438 1840 10438 0 net22
rlabel metal1 1978 9588 1978 9588 0 net23
rlabel metal2 2346 14722 2346 14722 0 net24
rlabel metal1 3381 2278 3381 2278 0 net25
rlabel metal2 2438 6698 2438 6698 0 net26
rlabel metal1 2208 3502 2208 3502 0 net27
rlabel metal2 7590 6290 7590 6290 0 net28
rlabel metal1 7314 3706 7314 3706 0 net29
rlabel metal2 13478 5678 13478 5678 0 net3
rlabel metal1 6900 3978 6900 3978 0 net30
rlabel metal1 12558 13906 12558 13906 0 net31
rlabel metal2 15502 15232 15502 15232 0 net32
rlabel via2 13938 20757 13938 20757 0 net33
rlabel metal2 14398 23205 14398 23205 0 net34
rlabel metal2 14766 23392 14766 23392 0 net35
rlabel metal2 9890 16847 9890 16847 0 net36
rlabel metal1 27462 20570 27462 20570 0 net37
rlabel metal1 33074 21556 33074 21556 0 net38
rlabel metal1 27462 22542 27462 22542 0 net39
rlabel metal1 14490 14042 14490 14042 0 net4
rlabel metal2 31970 22814 31970 22814 0 net40
rlabel metal2 33442 23885 33442 23885 0 net41
rlabel metal1 15916 18054 15916 18054 0 net42
rlabel metal2 35098 24089 35098 24089 0 net43
rlabel via2 17434 20893 17434 20893 0 net44
rlabel metal2 12558 17204 12558 17204 0 net45
rlabel metal1 32706 21998 32706 21998 0 net46
rlabel metal1 33166 21624 33166 21624 0 net47
rlabel metal1 37214 24310 37214 24310 0 net48
rlabel metal1 37582 23494 37582 23494 0 net49
rlabel metal1 13800 12818 13800 12818 0 net5
rlabel metal2 16974 16303 16974 16303 0 net50
rlabel metal1 14306 19278 14306 19278 0 net51
rlabel metal1 20056 19754 20056 19754 0 net52
rlabel metal2 40710 24072 40710 24072 0 net53
rlabel metal1 39284 23562 39284 23562 0 net54
rlabel metal3 14812 24344 14812 24344 0 net55
rlabel metal1 15962 20026 15962 20026 0 net56
rlabel metal2 14306 24378 14306 24378 0 net57
rlabel metal1 27048 24242 27048 24242 0 net58
rlabel metal1 25070 22984 25070 22984 0 net59
rlabel metal1 6348 6630 6348 6630 0 net6
rlabel metal1 26588 23018 26588 23018 0 net60
rlabel metal2 25806 23188 25806 23188 0 net61
rlabel via3 14421 21964 14421 21964 0 net62
rlabel metal1 25116 5610 25116 5610 0 net63
rlabel metal1 28014 2618 28014 2618 0 net64
rlabel metal1 29808 2618 29808 2618 0 net65
rlabel metal2 33534 3842 33534 3842 0 net66
rlabel metal2 36386 5814 36386 5814 0 net67
rlabel metal2 43746 23868 43746 23868 0 net68
rlabel metal2 45402 21369 45402 21369 0 net69
rlabel metal1 2944 7174 2944 7174 0 net7
rlabel metal1 45540 24072 45540 24072 0 net70
rlabel metal2 46874 20621 46874 20621 0 net71
rlabel metal2 46966 21148 46966 21148 0 net72
rlabel metal2 47150 20502 47150 20502 0 net73
rlabel metal2 44850 18224 44850 18224 0 net74
rlabel metal1 45034 23596 45034 23596 0 net75
rlabel metal2 45770 21165 45770 21165 0 net76
rlabel metal2 49266 20944 49266 20944 0 net77
rlabel metal2 47426 19754 47426 19754 0 net78
rlabel metal2 48530 19822 48530 19822 0 net79
rlabel metal1 3634 15402 3634 15402 0 net8
rlabel metal2 47058 21216 47058 21216 0 net80
rlabel metal1 47794 21318 47794 21318 0 net81
rlabel metal2 5934 20026 5934 20026 0 net82
rlabel via2 1794 13277 1794 13277 0 net83
rlabel metal1 13110 19176 13110 19176 0 net84
rlabel metal1 1794 19380 1794 19380 0 net85
rlabel metal2 4094 20349 4094 20349 0 net86
rlabel metal1 2024 23494 2024 23494 0 net87
rlabel metal1 1840 20910 1840 20910 0 net88
rlabel metal1 1794 21556 1794 21556 0 net89
rlabel metal2 13386 14790 13386 14790 0 net9
rlabel metal2 3404 16252 3404 16252 0 net90
rlabel metal1 1886 21998 1886 21998 0 net91
rlabel metal1 1840 22610 1840 22610 0 net92
rlabel metal1 13570 21862 13570 21862 0 net93
rlabel via2 1794 13923 1794 13923 0 net94
rlabel metal2 4002 21845 4002 21845 0 net95
rlabel metal2 3634 16150 3634 16150 0 net96
rlabel metal2 6118 21148 6118 21148 0 net97
rlabel metal1 4784 14518 4784 14518 0 net98
rlabel metal1 4922 12750 4922 12750 0 net99
rlabel metal2 38778 2098 38778 2098 0 prog_clk
rlabel metal1 41492 24174 41492 24174 0 prog_reset
rlabel metal1 18722 16966 18722 16966 0 sb_8__0_.mem_left_track_1.ccff_head
rlabel metal2 25254 19516 25254 19516 0 sb_8__0_.mem_left_track_1.ccff_tail
rlabel metal1 28612 16626 28612 16626 0 sb_8__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 16698 20570 16698 20570 0 sb_8__0_.mem_left_track_11.ccff_head
rlabel metal1 17250 23018 17250 23018 0 sb_8__0_.mem_left_track_11.ccff_tail
rlabel metal1 18722 22746 18722 22746 0 sb_8__0_.mem_left_track_11.mem_out\[0\]
rlabel metal1 16744 21454 16744 21454 0 sb_8__0_.mem_left_track_13.ccff_tail
rlabel metal1 18998 23800 18998 23800 0 sb_8__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 15318 20978 15318 20978 0 sb_8__0_.mem_left_track_15.ccff_tail
rlabel metal2 21482 23018 21482 23018 0 sb_8__0_.mem_left_track_15.mem_out\[0\]
rlabel metal1 17434 22202 17434 22202 0 sb_8__0_.mem_left_track_17.ccff_tail
rlabel metal2 23782 23358 23782 23358 0 sb_8__0_.mem_left_track_17.mem_out\[0\]
rlabel metal1 23920 21454 23920 21454 0 sb_8__0_.mem_left_track_19.ccff_tail
rlabel metal1 23828 21590 23828 21590 0 sb_8__0_.mem_left_track_19.mem_out\[0\]
rlabel metal1 26680 18938 26680 18938 0 sb_8__0_.mem_left_track_29.ccff_tail
rlabel metal1 26910 20366 26910 20366 0 sb_8__0_.mem_left_track_29.mem_out\[0\]
rlabel metal1 17894 19924 17894 19924 0 sb_8__0_.mem_left_track_3.ccff_tail
rlabel metal1 20509 19142 20509 19142 0 sb_8__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 26949 22202 26949 22202 0 sb_8__0_.mem_left_track_31.ccff_tail
rlabel metal1 27784 19686 27784 19686 0 sb_8__0_.mem_left_track_31.mem_out\[0\]
rlabel metal2 26634 23052 26634 23052 0 sb_8__0_.mem_left_track_33.ccff_tail
rlabel metal1 27738 22508 27738 22508 0 sb_8__0_.mem_left_track_33.mem_out\[0\]
rlabel metal1 29072 23290 29072 23290 0 sb_8__0_.mem_left_track_35.ccff_tail
rlabel metal1 28888 23494 28888 23494 0 sb_8__0_.mem_left_track_35.mem_out\[0\]
rlabel metal1 29578 22406 29578 22406 0 sb_8__0_.mem_left_track_45.ccff_tail
rlabel via1 30774 22073 30774 22073 0 sb_8__0_.mem_left_track_45.mem_out\[0\]
rlabel metal2 27738 20672 27738 20672 0 sb_8__0_.mem_left_track_47.ccff_tail
rlabel metal2 30222 20842 30222 20842 0 sb_8__0_.mem_left_track_47.mem_out\[0\]
rlabel metal1 28612 18054 28612 18054 0 sb_8__0_.mem_left_track_49.ccff_tail
rlabel metal1 29348 19142 29348 19142 0 sb_8__0_.mem_left_track_49.mem_out\[0\]
rlabel metal1 19688 19890 19688 19890 0 sb_8__0_.mem_left_track_5.ccff_tail
rlabel metal2 19734 21148 19734 21148 0 sb_8__0_.mem_left_track_5.mem_out\[0\]
rlabel metal1 28842 17680 28842 17680 0 sb_8__0_.mem_left_track_51.mem_out\[0\]
rlabel metal2 20654 19822 20654 19822 0 sb_8__0_.mem_left_track_7.ccff_tail
rlabel metal1 21758 19686 21758 19686 0 sb_8__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 19090 20332 19090 20332 0 sb_8__0_.mem_left_track_9.mem_out\[0\]
rlabel metal1 25070 15062 25070 15062 0 sb_8__0_.mem_top_track_0.ccff_tail
rlabel metal1 38686 22406 38686 22406 0 sb_8__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 24748 16014 24748 16014 0 sb_8__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 21298 12410 21298 12410 0 sb_8__0_.mem_top_track_10.ccff_head
rlabel metal1 17250 9962 17250 9962 0 sb_8__0_.mem_top_track_10.ccff_tail
rlabel metal2 24058 14926 24058 14926 0 sb_8__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 21436 12750 21436 12750 0 sb_8__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 16284 8874 16284 8874 0 sb_8__0_.mem_top_track_12.ccff_tail
rlabel metal1 20654 14450 20654 14450 0 sb_8__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 15548 10098 15548 10098 0 sb_8__0_.mem_top_track_14.ccff_tail
rlabel via2 14766 9469 14766 9469 0 sb_8__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 14628 12682 14628 12682 0 sb_8__0_.mem_top_track_16.ccff_tail
rlabel metal2 15042 10064 15042 10064 0 sb_8__0_.mem_top_track_16.mem_out\[0\]
rlabel via1 17427 13702 17427 13702 0 sb_8__0_.mem_top_track_18.ccff_tail
rlabel metal1 16790 13226 16790 13226 0 sb_8__0_.mem_top_track_18.mem_out\[0\]
rlabel metal2 21206 9690 21206 9690 0 sb_8__0_.mem_top_track_2.ccff_tail
rlabel metal1 25162 14416 25162 14416 0 sb_8__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 13892 7922 13892 7922 0 sb_8__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 18124 15334 18124 15334 0 sb_8__0_.mem_top_track_20.ccff_tail
rlabel metal2 17342 14722 17342 14722 0 sb_8__0_.mem_top_track_20.mem_out\[0\]
rlabel metal2 16330 14620 16330 14620 0 sb_8__0_.mem_top_track_22.ccff_tail
rlabel metal1 14904 14926 14904 14926 0 sb_8__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 15548 13498 15548 13498 0 sb_8__0_.mem_top_track_24.ccff_tail
rlabel metal1 15502 13362 15502 13362 0 sb_8__0_.mem_top_track_24.mem_out\[0\]
rlabel metal1 12558 11730 12558 11730 0 sb_8__0_.mem_top_track_26.ccff_tail
rlabel metal2 12098 11900 12098 11900 0 sb_8__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 13432 9418 13432 9418 0 sb_8__0_.mem_top_track_28.ccff_tail
rlabel metal1 11960 9622 11960 9622 0 sb_8__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 13754 13940 13754 13940 0 sb_8__0_.mem_top_track_30.ccff_tail
rlabel metal1 12328 13226 12328 13226 0 sb_8__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 12972 17714 12972 17714 0 sb_8__0_.mem_top_track_32.ccff_tail
rlabel metal1 13432 14926 13432 14926 0 sb_8__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 13478 19312 13478 19312 0 sb_8__0_.mem_top_track_34.ccff_tail
rlabel metal1 13110 17068 13110 17068 0 sb_8__0_.mem_top_track_34.mem_out\[0\]
rlabel metal2 9890 21046 9890 21046 0 sb_8__0_.mem_top_track_36.ccff_tail
rlabel metal2 11178 19516 11178 19516 0 sb_8__0_.mem_top_track_36.mem_out\[0\]
rlabel metal1 4876 18666 4876 18666 0 sb_8__0_.mem_top_track_38.ccff_tail
rlabel metal2 7958 16065 7958 16065 0 sb_8__0_.mem_top_track_38.mem_out\[0\]
rlabel metal1 19688 13226 19688 13226 0 sb_8__0_.mem_top_track_4.ccff_tail
rlabel metal1 22862 13804 22862 13804 0 sb_8__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 16974 11050 16974 11050 0 sb_8__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 7774 21590 7774 21590 0 sb_8__0_.mem_top_track_40.ccff_tail
rlabel metal1 7590 18598 7590 18598 0 sb_8__0_.mem_top_track_40.mem_out\[0\]
rlabel metal1 8694 20978 8694 20978 0 sb_8__0_.mem_top_track_42.ccff_tail
rlabel metal1 9430 21624 9430 21624 0 sb_8__0_.mem_top_track_42.mem_out\[0\]
rlabel metal2 13386 20672 13386 20672 0 sb_8__0_.mem_top_track_44.ccff_tail
rlabel via1 13570 21301 13570 21301 0 sb_8__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 15180 19890 15180 19890 0 sb_8__0_.mem_top_track_46.ccff_tail
rlabel metal1 14582 20366 14582 20366 0 sb_8__0_.mem_top_track_46.mem_out\[0\]
rlabel metal1 16790 17714 16790 17714 0 sb_8__0_.mem_top_track_48.ccff_tail
rlabel metal1 15502 18632 15502 18632 0 sb_8__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 18308 17238 18308 17238 0 sb_8__0_.mem_top_track_50.mem_out\[0\]
rlabel metal2 21942 14824 21942 14824 0 sb_8__0_.mem_top_track_6.ccff_tail
rlabel metal1 21390 17068 21390 17068 0 sb_8__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 19872 15402 19872 15402 0 sb_8__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 23828 14518 23828 14518 0 sb_8__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 21022 13498 21022 13498 0 sb_8__0_.mem_top_track_8.mem_out\[1\]
rlabel metal1 3864 18666 3864 18666 0 sb_8__0_.mux_left_track_1.out
rlabel metal1 25162 19958 25162 19958 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27278 16422 27278 16422 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23782 19958 23782 19958 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 4324 12886 4324 12886 0 sb_8__0_.mux_left_track_11.out
rlabel metal2 15962 24208 15962 24208 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 4232 12206 4232 12206 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 18354 17680 18354 17680 0 sb_8__0_.mux_left_track_13.out
rlabel metal3 17273 23732 17273 23732 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 15594 21403 15594 21403 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6394 21998 6394 21998 0 sb_8__0_.mux_left_track_15.out
rlabel metal1 16882 20842 16882 20842 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14582 20808 14582 20808 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3634 12886 3634 12886 0 sb_8__0_.mux_left_track_17.out
rlabel metal1 16238 21046 16238 21046 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 14076 18904 14076 18904 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19412 15334 19412 15334 0 sb_8__0_.mux_left_track_19.out
rlabel metal1 22494 21386 22494 21386 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19918 15470 19918 15470 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7820 15130 7820 15130 0 sb_8__0_.mux_left_track_29.out
rlabel metal1 26404 20298 26404 20298 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21114 14773 21114 14773 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21390 16592 21390 16592 0 sb_8__0_.mux_left_track_3.out
rlabel metal2 17710 20332 17710 20332 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 17250 19941 17250 19941 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15226 17306 15226 17306 0 sb_8__0_.mux_left_track_31.out
rlabel metal1 26818 21658 26818 21658 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18952 17850 18952 17850 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 2231 23460 2231 23460 0 sb_8__0_.mux_left_track_33.out
rlabel metal1 24288 21998 24288 21998 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 3358 8925 3358 8925 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 9361 12444 9361 12444 0 sb_8__0_.mux_left_track_35.out
rlabel metal2 30590 22967 30590 22967 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7912 8602 7912 8602 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20309 15878 20309 15878 0 sb_8__0_.mux_left_track_45.out
rlabel metal2 30130 21590 30130 21590 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24472 20910 24472 20910 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13570 16082 13570 16082 0 sb_8__0_.mux_left_track_47.out
rlabel metal1 27922 20774 27922 20774 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13754 15436 13754 15436 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12926 14297 12926 14297 0 sb_8__0_.mux_left_track_49.out
rlabel metal2 30222 19516 30222 19516 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21574 15640 21574 15640 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 14950 21947 14950 21947 0 sb_8__0_.mux_left_track_5.out
rlabel metal1 17250 20570 17250 20570 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16928 20298 16928 20298 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel via1 5750 13770 5750 13770 0 sb_8__0_.mux_left_track_51.out
rlabel metal1 21643 17578 21643 17578 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16974 16082 16974 16082 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13662 18632 13662 18632 0 sb_8__0_.mux_left_track_7.out
rlabel metal1 22586 19414 22586 19414 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 19482 22862 19482 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22034 19040 22034 19040 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 1058 22413 1058 22413 0 sb_8__0_.mux_left_track_9.out
rlabel metal1 18538 20536 18538 20536 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12788 15572 12788 15572 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19550 18972 19550 18972 0 sb_8__0_.mux_top_track_0.out
rlabel metal2 27094 17408 27094 17408 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27738 16490 27738 16490 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26634 16456 26634 16456 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23414 16507 23414 16507 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23598 19108 23598 19108 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18676 16082 18676 16082 0 sb_8__0_.mux_top_track_10.out
rlabel metal1 21643 12818 21643 12818 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21160 12954 21160 12954 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20838 12614 20838 12614 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15134 9146 15134 9146 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal3 17204 14756 17204 14756 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 14398 16473 14398 16473 0 sb_8__0_.mux_top_track_12.out
rlabel metal1 16054 10540 16054 10540 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14582 8602 14582 8602 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14628 16558 14628 16558 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 13478 14348 13478 14348 0 sb_8__0_.mux_top_track_14.out
rlabel metal1 15916 10778 15916 10778 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13662 10438 13662 10438 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15042 10438 15042 10438 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 10994 15963 10994 15963 0 sb_8__0_.mux_top_track_16.out
rlabel metal1 15686 12614 15686 12614 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12673 12818 12673 12818 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12512 12954 12512 12954 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 14950 23936 14950 23936 0 sb_8__0_.mux_top_track_18.out
rlabel metal2 17894 16762 17894 16762 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13662 14042 13662 14042 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17756 19788 17756 19788 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19090 19652 19090 19652 0 sb_8__0_.mux_top_track_2.out
rlabel metal1 24840 13974 24840 13974 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25392 14042 25392 14042 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22080 9622 22080 9622 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15272 8058 15272 8058 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19182 19346 19182 19346 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33718 21998 33718 21998 0 sb_8__0_.mux_top_track_20.out
rlabel metal2 15870 16388 15870 16388 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16882 16864 16882 16864 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34914 22746 34914 22746 0 sb_8__0_.mux_top_track_22.out
rlabel metal1 14398 13804 14398 13804 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19642 14654 19642 14654 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31970 21964 31970 21964 0 sb_8__0_.mux_top_track_24.out
rlabel metal1 14168 12954 14168 12954 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14398 14416 14398 14416 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32430 22576 32430 22576 0 sb_8__0_.mux_top_track_26.out
rlabel metal2 10626 11968 10626 11968 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 3703 18020 3703 18020 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32430 10511 32430 10511 0 sb_8__0_.mux_top_track_28.out
rlabel metal1 10442 10234 10442 10234 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11132 9010 11132 9010 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33718 23018 33718 23018 0 sb_8__0_.mux_top_track_30.out
rlabel metal2 12558 13872 12558 13872 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12098 15385 12098 15385 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32568 21114 32568 21114 0 sb_8__0_.mux_top_track_32.out
rlabel metal1 12834 14858 12834 14858 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32706 19533 32706 19533 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33028 23698 33028 23698 0 sb_8__0_.mux_top_track_34.out
rlabel metal1 12512 17306 12512 17306 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 11454 19397 11454 19397 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4094 11186 4094 11186 0 sb_8__0_.mux_top_track_36.out
rlabel metal1 10718 18938 10718 18938 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 1794 10370 1794 10370 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 4278 10064 4278 10064 0 sb_8__0_.mux_top_track_38.out
rlabel metal1 7176 16218 7176 16218 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 4761 11492 4761 11492 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18216 16422 18216 16422 0 sb_8__0_.mux_top_track_4.out
rlabel metal1 20194 12852 20194 12852 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18492 12954 18492 12954 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17388 12954 17388 12954 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 15962 13163 15962 13163 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16100 14042 16100 14042 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 5888 8602 5888 8602 0 sb_8__0_.mux_top_track_40.out
rlabel metal1 7912 17306 7912 17306 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 1794 23562 1794 23562 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9154 8194 9154 8194 0 sb_8__0_.mux_top_track_42.out
rlabel metal1 8326 21012 8326 21012 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7774 21046 7774 21046 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19734 13770 19734 13770 0 sb_8__0_.mux_top_track_44.out
rlabel metal1 17710 19482 17710 19482 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11638 19822 11638 19822 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32338 21522 32338 21522 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32890 15164 32890 15164 0 sb_8__0_.mux_top_track_46.out
rlabel metal1 18262 18870 18262 18870 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11178 18394 11178 18394 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13432 20026 13432 20026 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 2024 10574 2024 10574 0 sb_8__0_.mux_top_track_48.out
rlabel metal1 17526 18122 17526 18122 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13754 17850 13754 17850 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15042 18479 15042 18479 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19458 14008 19458 14008 0 sb_8__0_.mux_top_track_50.out
rlabel metal2 20746 18632 20746 18632 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 13018 16677 13018 16677 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19136 13906 19136 13906 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20654 22593 20654 22593 0 sb_8__0_.mux_top_track_6.out
rlabel metal2 20746 16796 20746 16796 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 16558 22862 16558 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20240 14926 20240 14926 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19780 14994 19780 14994 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19872 14858 19872 14858 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19228 17714 19228 17714 0 sb_8__0_.mux_top_track_8.out
rlabel metal1 23552 13226 23552 13226 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23184 13226 23184 13226 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22862 13192 22862 13192 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15686 8602 15686 8602 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20102 14246 20102 14246 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 44758 25340 44758 25340 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal2 45494 25296 45494 25296 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 46368 24174 46368 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 46736 23698 46736 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 47564 24174 47564 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 47932 23086 47932 23086 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 44344 23698 44344 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel via1 44206 23749 44206 23749 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel via2 49082 21981 49082 21981 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 49082 22763 49082 22763 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 48346 22831 48346 22831 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 48162 23698 48162 23698 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 41446 2948 41446 2948 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 44114 2200 44114 2200 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 46782 2166 46782 2166 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 49450 2132 49450 2132 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
