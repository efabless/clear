magic
tech sky130A
magscale 1 2
timestamp 1656943510
<< viali >>
rect 6561 14025 6595 14059
rect 6837 14025 6871 14059
rect 7757 14025 7791 14059
rect 8217 14025 8251 14059
rect 8585 14025 8619 14059
rect 8861 14025 8895 14059
rect 9137 14025 9171 14059
rect 9965 14025 9999 14059
rect 11161 14025 11195 14059
rect 12633 14025 12667 14059
rect 13369 14025 13403 14059
rect 13737 14025 13771 14059
rect 14105 14025 14139 14059
rect 11897 13957 11931 13991
rect 6377 13889 6411 13923
rect 7021 13889 7055 13923
rect 7113 13889 7147 13923
rect 7573 13889 7607 13923
rect 8401 13889 8435 13923
rect 8769 13889 8803 13923
rect 10149 13889 10183 13923
rect 11345 13889 11379 13923
rect 12817 13889 12851 13923
rect 13553 13889 13587 13923
rect 13921 13889 13955 13923
rect 15209 13889 15243 13923
rect 6101 13821 6135 13855
rect 10333 13821 10367 13855
rect 7389 13753 7423 13787
rect 11621 13685 11655 13719
rect 15025 13685 15059 13719
rect 5825 13345 5859 13379
rect 6469 13345 6503 13379
rect 6653 13345 6687 13379
rect 7481 13345 7515 13379
rect 9781 13345 9815 13379
rect 11621 13345 11655 13379
rect 12265 13345 12299 13379
rect 12449 13345 12483 13379
rect 7297 13277 7331 13311
rect 7757 13277 7791 13311
rect 12173 13277 12207 13311
rect 13001 13277 13035 13311
rect 5549 13209 5583 13243
rect 9689 13209 9723 13243
rect 10057 13209 10091 13243
rect 5181 13141 5215 13175
rect 5641 13141 5675 13175
rect 6009 13141 6043 13175
rect 6377 13141 6411 13175
rect 6837 13141 6871 13175
rect 7205 13141 7239 13175
rect 9229 13141 9263 13175
rect 9597 13141 9631 13175
rect 10977 13141 11011 13175
rect 11345 13141 11379 13175
rect 11437 13141 11471 13175
rect 11805 13141 11839 13175
rect 12633 13141 12667 13175
rect 13829 13141 13863 13175
rect 2789 12937 2823 12971
rect 3341 12937 3375 12971
rect 3893 12937 3927 12971
rect 3985 12937 4019 12971
rect 4445 12937 4479 12971
rect 5181 12937 5215 12971
rect 5825 12937 5859 12971
rect 6561 12937 6595 12971
rect 9229 12937 9263 12971
rect 9597 12937 9631 12971
rect 11621 12937 11655 12971
rect 11989 12937 12023 12971
rect 13553 12937 13587 12971
rect 13921 12937 13955 12971
rect 6837 12869 6871 12903
rect 8677 12869 8711 12903
rect 10057 12869 10091 12903
rect 12081 12869 12115 12903
rect 12541 12869 12575 12903
rect 14381 12869 14415 12903
rect 2053 12801 2087 12835
rect 2421 12801 2455 12835
rect 5273 12801 5307 12835
rect 9137 12801 9171 12835
rect 9965 12801 9999 12835
rect 13461 12801 13495 12835
rect 14289 12801 14323 12835
rect 2605 12733 2639 12767
rect 4077 12733 4111 12767
rect 5365 12733 5399 12767
rect 6929 12733 6963 12767
rect 9321 12733 9355 12767
rect 10241 12733 10275 12767
rect 12265 12733 12299 12767
rect 13645 12733 13679 12767
rect 14473 12733 14507 12767
rect 1869 12665 1903 12699
rect 8769 12665 8803 12699
rect 10517 12665 10551 12699
rect 2237 12597 2271 12631
rect 3525 12597 3559 12631
rect 4813 12597 4847 12631
rect 12633 12597 12667 12631
rect 13093 12597 13127 12631
rect 14841 12597 14875 12631
rect 2237 12393 2271 12427
rect 9689 12393 9723 12427
rect 13829 12393 13863 12427
rect 14105 12393 14139 12427
rect 4169 12325 4203 12359
rect 3065 12257 3099 12291
rect 4997 12257 5031 12291
rect 6653 12257 6687 12291
rect 7481 12257 7515 12291
rect 8309 12257 8343 12291
rect 9597 12257 9631 12291
rect 10241 12257 10275 12291
rect 11529 12257 11563 12291
rect 12541 12257 12575 12291
rect 13369 12257 13403 12291
rect 14657 12257 14691 12291
rect 15209 12257 15243 12291
rect 2053 12189 2087 12223
rect 7297 12189 7331 12223
rect 8217 12189 8251 12223
rect 9229 12189 9263 12223
rect 10149 12189 10183 12223
rect 11253 12189 11287 12223
rect 12449 12189 12483 12223
rect 13185 12189 13219 12223
rect 14565 12189 14599 12223
rect 17693 12189 17727 12223
rect 17785 12189 17819 12223
rect 3157 12121 3191 12155
rect 3249 12121 3283 12155
rect 3801 12121 3835 12155
rect 4261 12121 4295 12155
rect 4813 12121 4847 12155
rect 6469 12121 6503 12155
rect 12357 12121 12391 12155
rect 1869 12053 1903 12087
rect 3617 12053 3651 12087
rect 4445 12053 4479 12087
rect 4905 12053 4939 12087
rect 6101 12053 6135 12087
rect 6561 12053 6595 12087
rect 6929 12053 6963 12087
rect 7389 12053 7423 12087
rect 7757 12053 7791 12087
rect 8125 12053 8159 12087
rect 8585 12053 8619 12087
rect 10057 12053 10091 12087
rect 10517 12053 10551 12087
rect 10885 12053 10919 12087
rect 11345 12053 11379 12087
rect 11989 12053 12023 12087
rect 12817 12053 12851 12087
rect 13277 12053 13311 12087
rect 14473 12053 14507 12087
rect 15393 12053 15427 12087
rect 17969 12053 18003 12087
rect 2697 11849 2731 11883
rect 2973 11849 3007 11883
rect 3341 11849 3375 11883
rect 3433 11849 3467 11883
rect 4353 11849 4387 11883
rect 5457 11849 5491 11883
rect 5825 11849 5859 11883
rect 6653 11849 6687 11883
rect 7113 11849 7147 11883
rect 8309 11849 8343 11883
rect 12633 11849 12667 11883
rect 13093 11849 13127 11883
rect 15945 11849 15979 11883
rect 16773 11849 16807 11883
rect 4445 11781 4479 11815
rect 12173 11781 12207 11815
rect 17693 11781 17727 11815
rect 2053 11713 2087 11747
rect 2421 11713 2455 11747
rect 2513 11713 2547 11747
rect 5273 11713 5307 11747
rect 7021 11713 7055 11747
rect 9137 11713 9171 11747
rect 9965 11713 9999 11747
rect 10425 11713 10459 11747
rect 12725 11713 12759 11747
rect 13185 11713 13219 11747
rect 15025 11713 15059 11747
rect 15117 11713 15151 11747
rect 16405 11713 16439 11747
rect 17877 11713 17911 11747
rect 3617 11645 3651 11679
rect 4537 11645 4571 11679
rect 5917 11645 5951 11679
rect 6101 11645 6135 11679
rect 7205 11645 7239 11679
rect 7757 11645 7791 11679
rect 8125 11645 8159 11679
rect 8217 11645 8251 11679
rect 9229 11645 9263 11679
rect 9413 11645 9447 11679
rect 10057 11645 10091 11679
rect 10241 11645 10275 11679
rect 12541 11645 12575 11679
rect 14933 11645 14967 11679
rect 16037 11645 16071 11679
rect 16129 11645 16163 11679
rect 1869 11577 1903 11611
rect 8769 11577 8803 11611
rect 2237 11509 2271 11543
rect 3985 11509 4019 11543
rect 6469 11509 6503 11543
rect 7573 11509 7607 11543
rect 8677 11509 8711 11543
rect 9597 11509 9631 11543
rect 14565 11509 14599 11543
rect 15485 11509 15519 11543
rect 15577 11509 15611 11543
rect 16957 11509 16991 11543
rect 18061 11509 18095 11543
rect 7757 11305 7791 11339
rect 8953 11305 8987 11339
rect 9781 11305 9815 11339
rect 4537 11237 4571 11271
rect 13093 11237 13127 11271
rect 16129 11237 16163 11271
rect 16957 11237 16991 11271
rect 18061 11237 18095 11271
rect 3065 11169 3099 11203
rect 3249 11169 3283 11203
rect 8217 11169 8251 11203
rect 8309 11169 8343 11203
rect 8585 11169 8619 11203
rect 9597 11169 9631 11203
rect 14565 11169 14599 11203
rect 14749 11169 14783 11203
rect 15393 11169 15427 11203
rect 15485 11169 15519 11203
rect 16681 11169 16715 11203
rect 17417 11169 17451 11203
rect 17509 11169 17543 11203
rect 2973 11101 3007 11135
rect 5650 11101 5684 11135
rect 5917 11101 5951 11135
rect 7665 11101 7699 11135
rect 8125 11101 8159 11135
rect 9321 11101 9355 11135
rect 9413 11101 9447 11135
rect 11713 11101 11747 11135
rect 15301 11101 15335 11135
rect 16497 11101 16531 11135
rect 17877 11101 17911 11135
rect 18245 11101 18279 11135
rect 9965 11033 9999 11067
rect 11958 11033 11992 11067
rect 14473 11033 14507 11067
rect 18521 11033 18555 11067
rect 2605 10965 2639 10999
rect 14105 10965 14139 10999
rect 14933 10965 14967 10999
rect 16589 10965 16623 10999
rect 17325 10965 17359 10999
rect 2329 10761 2363 10795
rect 2789 10761 2823 10795
rect 8217 10761 8251 10795
rect 11529 10761 11563 10795
rect 14381 10761 14415 10795
rect 14657 10761 14691 10795
rect 15117 10761 15151 10795
rect 16681 10761 16715 10795
rect 2145 10693 2179 10727
rect 3709 10693 3743 10727
rect 5926 10693 5960 10727
rect 13268 10693 13302 10727
rect 17049 10693 17083 10727
rect 17509 10693 17543 10727
rect 3617 10625 3651 10659
rect 7104 10625 7138 10659
rect 9422 10625 9456 10659
rect 10140 10625 10174 10659
rect 12642 10625 12676 10659
rect 15025 10625 15059 10659
rect 17877 10625 17911 10659
rect 2881 10557 2915 10591
rect 2973 10557 3007 10591
rect 3893 10557 3927 10591
rect 6193 10557 6227 10591
rect 6837 10557 6871 10591
rect 9689 10557 9723 10591
rect 9873 10557 9907 10591
rect 12909 10557 12943 10591
rect 13001 10557 13035 10591
rect 14473 10557 14507 10591
rect 15301 10557 15335 10591
rect 17141 10557 17175 10591
rect 17233 10557 17267 10591
rect 8309 10489 8343 10523
rect 16405 10489 16439 10523
rect 17693 10489 17727 10523
rect 2421 10421 2455 10455
rect 3249 10421 3283 10455
rect 4169 10421 4203 10455
rect 4813 10421 4847 10455
rect 11253 10421 11287 10455
rect 18061 10421 18095 10455
rect 6561 10217 6595 10251
rect 9045 10217 9079 10251
rect 11437 10217 11471 10251
rect 16405 10217 16439 10251
rect 16589 10217 16623 10251
rect 17693 10217 17727 10251
rect 2513 10081 2547 10115
rect 2605 10081 2639 10115
rect 3065 10081 3099 10115
rect 17049 10081 17083 10115
rect 17233 10081 17267 10115
rect 1961 10013 1995 10047
rect 2421 10013 2455 10047
rect 4537 10013 4571 10047
rect 4804 10013 4838 10047
rect 7941 10013 7975 10047
rect 10158 10013 10192 10047
rect 10425 10013 10459 10047
rect 12817 10013 12851 10047
rect 17877 10013 17911 10047
rect 7674 9945 7708 9979
rect 12572 9945 12606 9979
rect 1777 9877 1811 9911
rect 2053 9877 2087 9911
rect 3341 9877 3375 9911
rect 5917 9877 5951 9911
rect 16957 9877 16991 9911
rect 17509 9877 17543 9911
rect 18061 9877 18095 9911
rect 5580 9605 5614 9639
rect 13032 9605 13066 9639
rect 2053 9537 2087 9571
rect 2605 9537 2639 9571
rect 7297 9537 7331 9571
rect 8401 9537 8435 9571
rect 8841 9537 8875 9571
rect 17693 9537 17727 9571
rect 17877 9537 17911 9571
rect 18245 9537 18279 9571
rect 2697 9469 2731 9503
rect 2789 9469 2823 9503
rect 5825 9469 5859 9503
rect 7665 9469 7699 9503
rect 8585 9469 8619 9503
rect 13277 9469 13311 9503
rect 1869 9401 1903 9435
rect 4445 9401 4479 9435
rect 2237 9333 2271 9367
rect 9965 9333 9999 9367
rect 11897 9333 11931 9367
rect 15393 9333 15427 9367
rect 18061 9333 18095 9367
rect 18429 9333 18463 9367
rect 2145 9129 2179 9163
rect 2513 9129 2547 9163
rect 6837 9129 6871 9163
rect 10149 9129 10183 9163
rect 11989 9129 12023 9163
rect 15301 9129 15335 9163
rect 16405 9129 16439 9163
rect 18061 9129 18095 9163
rect 2421 9061 2455 9095
rect 8769 9061 8803 9095
rect 3065 8993 3099 9027
rect 11529 8993 11563 9027
rect 14565 8993 14599 9027
rect 16037 8993 16071 9027
rect 5365 8925 5399 8959
rect 5457 8925 5491 8959
rect 7389 8925 7423 8959
rect 11262 8925 11296 8959
rect 13369 8925 13403 8959
rect 14749 8925 14783 8959
rect 15945 8925 15979 8959
rect 17509 8925 17543 8959
rect 2881 8857 2915 8891
rect 3341 8857 3375 8891
rect 5098 8857 5132 8891
rect 5724 8857 5758 8891
rect 7634 8857 7668 8891
rect 13124 8857 13158 8891
rect 17325 8857 17359 8891
rect 2973 8789 3007 8823
rect 3801 8789 3835 8823
rect 3985 8789 4019 8823
rect 14289 8789 14323 8823
rect 14657 8789 14691 8823
rect 15117 8789 15151 8823
rect 15485 8789 15519 8823
rect 15853 8789 15887 8823
rect 17693 8789 17727 8823
rect 1869 8585 1903 8619
rect 2329 8585 2363 8619
rect 12909 8585 12943 8619
rect 14381 8585 14415 8619
rect 15761 8585 15795 8619
rect 16313 8585 16347 8619
rect 17509 8585 17543 8619
rect 2789 8517 2823 8551
rect 4077 8517 4111 8551
rect 9312 8517 9346 8551
rect 13268 8517 13302 8551
rect 2697 8449 2731 8483
rect 3525 8449 3559 8483
rect 4988 8449 5022 8483
rect 7490 8449 7524 8483
rect 7757 8449 7791 8483
rect 9045 8449 9079 8483
rect 11529 8449 11563 8483
rect 11785 8449 11819 8483
rect 13001 8449 13035 8483
rect 17693 8449 17727 8483
rect 1961 8381 1995 8415
rect 2145 8381 2179 8415
rect 2973 8381 3007 8415
rect 3617 8381 3651 8415
rect 3801 8381 3835 8415
rect 4721 8381 4755 8415
rect 15853 8381 15887 8415
rect 16037 8381 16071 8415
rect 1501 8313 1535 8347
rect 6101 8313 6135 8347
rect 15209 8313 15243 8347
rect 17877 8313 17911 8347
rect 3157 8245 3191 8279
rect 6377 8245 6411 8279
rect 10425 8245 10459 8279
rect 15393 8245 15427 8279
rect 1501 8041 1535 8075
rect 1777 8041 1811 8075
rect 2145 8041 2179 8075
rect 2053 7973 2087 8007
rect 16957 7973 16991 8007
rect 2697 7905 2731 7939
rect 14933 7905 14967 7939
rect 15117 7905 15151 7939
rect 2605 7837 2639 7871
rect 4537 7837 4571 7871
rect 6929 7837 6963 7871
rect 8953 7837 8987 7871
rect 10517 7837 10551 7871
rect 12081 7837 12115 7871
rect 15209 7837 15243 7871
rect 17049 7837 17083 7871
rect 4782 7769 4816 7803
rect 7196 7769 7230 7803
rect 9198 7769 9232 7803
rect 10762 7769 10796 7803
rect 12348 7769 12382 7803
rect 2513 7701 2547 7735
rect 3157 7701 3191 7735
rect 5917 7701 5951 7735
rect 8309 7701 8343 7735
rect 10333 7701 10367 7735
rect 11897 7701 11931 7735
rect 13461 7701 13495 7735
rect 15577 7701 15611 7735
rect 17233 7701 17267 7735
rect 1777 7497 1811 7531
rect 2145 7497 2179 7531
rect 2605 7497 2639 7531
rect 2973 7497 3007 7531
rect 14565 7497 14599 7531
rect 14933 7497 14967 7531
rect 15393 7497 15427 7531
rect 17141 7497 17175 7531
rect 17509 7497 17543 7531
rect 2513 7429 2547 7463
rect 12326 7429 12360 7463
rect 4189 7361 4223 7395
rect 5650 7361 5684 7395
rect 5917 7361 5951 7395
rect 7869 7361 7903 7395
rect 10342 7361 10376 7395
rect 10609 7361 10643 7395
rect 12081 7361 12115 7395
rect 14473 7361 14507 7395
rect 15301 7361 15335 7395
rect 17049 7361 17083 7395
rect 17693 7361 17727 7395
rect 17877 7361 17911 7395
rect 18245 7361 18279 7395
rect 1501 7293 1535 7327
rect 1685 7293 1719 7327
rect 2421 7293 2455 7327
rect 4445 7293 4479 7327
rect 8125 7293 8159 7327
rect 14657 7293 14691 7327
rect 15577 7293 15611 7327
rect 16405 7293 16439 7327
rect 17233 7293 17267 7327
rect 13461 7225 13495 7259
rect 16681 7225 16715 7259
rect 3065 7157 3099 7191
rect 4537 7157 4571 7191
rect 6009 7157 6043 7191
rect 6745 7157 6779 7191
rect 9229 7157 9263 7191
rect 14105 7157 14139 7191
rect 18061 7157 18095 7191
rect 18429 7157 18463 7191
rect 1961 6953 1995 6987
rect 5825 6953 5859 6987
rect 15393 6953 15427 6987
rect 18153 6953 18187 6987
rect 12449 6885 12483 6919
rect 2421 6817 2455 6851
rect 2605 6817 2639 6851
rect 2881 6817 2915 6851
rect 12357 6817 12391 6851
rect 14749 6817 14783 6851
rect 14933 6817 14967 6851
rect 16221 6817 16255 6851
rect 16313 6817 16347 6851
rect 17141 6817 17175 6851
rect 1501 6749 1535 6783
rect 1869 6749 1903 6783
rect 3157 6749 3191 6783
rect 3893 6749 3927 6783
rect 4445 6749 4479 6783
rect 8493 6749 8527 6783
rect 9321 6749 9355 6783
rect 9577 6749 9611 6783
rect 13829 6749 13863 6783
rect 17049 6749 17083 6783
rect 17417 6749 17451 6783
rect 4690 6681 4724 6715
rect 8248 6681 8282 6715
rect 12090 6681 12124 6715
rect 13562 6681 13596 6715
rect 16129 6681 16163 6715
rect 1685 6613 1719 6647
rect 2329 6613 2363 6647
rect 3065 6613 3099 6647
rect 3525 6613 3559 6647
rect 3985 6613 4019 6647
rect 4261 6613 4295 6647
rect 7113 6613 7147 6647
rect 10701 6613 10735 6647
rect 10977 6613 11011 6647
rect 14473 6613 14507 6647
rect 15025 6613 15059 6647
rect 15761 6613 15795 6647
rect 16589 6613 16623 6647
rect 16957 6613 16991 6647
rect 1593 6409 1627 6443
rect 2329 6409 2363 6443
rect 3065 6409 3099 6443
rect 3433 6409 3467 6443
rect 3893 6409 3927 6443
rect 4261 6409 4295 6443
rect 13277 6409 13311 6443
rect 14013 6409 14047 6443
rect 14381 6409 14415 6443
rect 14841 6409 14875 6443
rect 15209 6409 15243 6443
rect 16221 6409 16255 6443
rect 16957 6409 16991 6443
rect 12164 6341 12198 6375
rect 13921 6341 13955 6375
rect 1777 6273 1811 6307
rect 2237 6273 2271 6307
rect 2973 6273 3007 6307
rect 5926 6273 5960 6307
rect 6193 6273 6227 6307
rect 7685 6273 7719 6307
rect 7941 6273 7975 6307
rect 9985 6273 10019 6307
rect 10241 6273 10275 6307
rect 11897 6273 11931 6307
rect 14749 6273 14783 6307
rect 15577 6273 15611 6307
rect 2513 6205 2547 6239
rect 3525 6205 3559 6239
rect 3617 6205 3651 6239
rect 4353 6205 4387 6239
rect 4537 6205 4571 6239
rect 6469 6205 6503 6239
rect 14105 6205 14139 6239
rect 14933 6205 14967 6239
rect 15669 6205 15703 6239
rect 15761 6205 15795 6239
rect 13553 6137 13587 6171
rect 18061 6137 18095 6171
rect 1869 6069 1903 6103
rect 2789 6069 2823 6103
rect 4813 6069 4847 6103
rect 6561 6069 6595 6103
rect 8861 6069 8895 6103
rect 16037 6069 16071 6103
rect 2789 5865 2823 5899
rect 3617 5865 3651 5899
rect 4077 5865 4111 5899
rect 5917 5865 5951 5899
rect 14197 5865 14231 5899
rect 15117 5865 15151 5899
rect 15577 5865 15611 5899
rect 16405 5865 16439 5899
rect 17509 5865 17543 5899
rect 18061 5865 18095 5899
rect 2605 5797 2639 5831
rect 7849 5797 7883 5831
rect 7941 5797 7975 5831
rect 8677 5797 8711 5831
rect 9689 5797 9723 5831
rect 10149 5797 10183 5831
rect 10333 5797 10367 5831
rect 17233 5797 17267 5831
rect 1961 5729 1995 5763
rect 2145 5729 2179 5763
rect 3065 5729 3099 5763
rect 4537 5729 4571 5763
rect 6745 5729 6779 5763
rect 12541 5729 12575 5763
rect 13645 5729 13679 5763
rect 14473 5729 14507 5763
rect 14657 5729 14691 5763
rect 16129 5729 16163 5763
rect 16957 5729 16991 5763
rect 1869 5661 1903 5695
rect 6653 5661 6687 5695
rect 7481 5661 7515 5695
rect 9321 5661 9355 5695
rect 10701 5661 10735 5695
rect 14749 5661 14783 5695
rect 16037 5661 16071 5695
rect 16865 5661 16899 5695
rect 17877 5661 17911 5695
rect 18245 5661 18279 5695
rect 3157 5593 3191 5627
rect 4782 5593 4816 5627
rect 6009 5593 6043 5627
rect 8217 5593 8251 5627
rect 11069 5593 11103 5627
rect 12633 5593 12667 5627
rect 13553 5593 13587 5627
rect 15945 5593 15979 5627
rect 16773 5593 16807 5627
rect 1501 5525 1535 5559
rect 2421 5525 2455 5559
rect 3249 5525 3283 5559
rect 3893 5525 3927 5559
rect 6193 5525 6227 5559
rect 6561 5525 6595 5559
rect 7389 5525 7423 5559
rect 9229 5525 9263 5559
rect 15209 5525 15243 5559
rect 17693 5525 17727 5559
rect 18429 5525 18463 5559
rect 1777 5321 1811 5355
rect 2605 5321 2639 5355
rect 3065 5321 3099 5355
rect 3525 5321 3559 5355
rect 3985 5321 4019 5355
rect 4905 5321 4939 5355
rect 5365 5321 5399 5355
rect 5733 5321 5767 5355
rect 6929 5321 6963 5355
rect 7665 5321 7699 5355
rect 11069 5321 11103 5355
rect 11299 5321 11333 5355
rect 13277 5321 13311 5355
rect 13645 5321 13679 5355
rect 14013 5321 14047 5355
rect 14105 5321 14139 5355
rect 14473 5321 14507 5355
rect 14841 5321 14875 5355
rect 15301 5321 15335 5355
rect 17601 5321 17635 5355
rect 4813 5253 4847 5287
rect 11621 5253 11655 5287
rect 11713 5253 11747 5287
rect 13185 5253 13219 5287
rect 15669 5253 15703 5287
rect 2145 5185 2179 5219
rect 2237 5185 2271 5219
rect 2513 5185 2547 5219
rect 2973 5185 3007 5219
rect 3893 5185 3927 5219
rect 6837 5185 6871 5219
rect 8125 5185 8159 5219
rect 8493 5185 8527 5219
rect 9413 5185 9447 5219
rect 10425 5185 10459 5219
rect 11196 5185 11230 5219
rect 15761 5185 15795 5219
rect 16129 5185 16163 5219
rect 16681 5185 16715 5219
rect 17049 5185 17083 5219
rect 17785 5185 17819 5219
rect 3249 5117 3283 5151
rect 4077 5117 4111 5151
rect 4721 5117 4755 5151
rect 5825 5117 5859 5151
rect 5917 5117 5951 5151
rect 7021 5117 7055 5151
rect 7757 5117 7791 5151
rect 7849 5117 7883 5151
rect 8861 5117 8895 5151
rect 9689 5117 9723 5151
rect 10793 5117 10827 5151
rect 12633 5117 12667 5151
rect 13369 5117 13403 5151
rect 14197 5117 14231 5151
rect 14933 5117 14967 5151
rect 15025 5117 15059 5151
rect 15853 5117 15887 5151
rect 9045 5049 9079 5083
rect 9873 5049 9907 5083
rect 10057 5049 10091 5083
rect 12817 5049 12851 5083
rect 1961 4981 1995 5015
rect 4445 4981 4479 5015
rect 5273 4981 5307 5015
rect 6469 4981 6503 5015
rect 7297 4981 7331 5015
rect 16313 4981 16347 5015
rect 16865 4981 16899 5015
rect 17969 4981 18003 5015
rect 2605 4777 2639 4811
rect 5273 4777 5307 4811
rect 6193 4777 6227 4811
rect 14289 4777 14323 4811
rect 14565 4777 14599 4811
rect 16129 4777 16163 4811
rect 16313 4777 16347 4811
rect 2237 4709 2271 4743
rect 2789 4709 2823 4743
rect 16497 4709 16531 4743
rect 3157 4641 3191 4675
rect 5549 4641 5583 4675
rect 5733 4641 5767 4675
rect 6745 4641 6779 4675
rect 6837 4641 6871 4675
rect 7389 4641 7423 4675
rect 9689 4641 9723 4675
rect 9873 4641 9907 4675
rect 10057 4641 10091 4675
rect 10977 4641 11011 4675
rect 12265 4641 12299 4675
rect 13277 4641 13311 4675
rect 1685 4573 1719 4607
rect 2053 4573 2087 4607
rect 2421 4573 2455 4607
rect 2973 4573 3007 4607
rect 3433 4573 3467 4607
rect 9321 4573 9355 4607
rect 10425 4573 10459 4607
rect 13645 4573 13679 4607
rect 15945 4573 15979 4607
rect 17509 4573 17543 4607
rect 17693 4573 17727 4607
rect 5825 4505 5859 4539
rect 8033 4505 8067 4539
rect 8493 4505 8527 4539
rect 8677 4505 8711 4539
rect 10793 4505 10827 4539
rect 11069 4505 11103 4539
rect 11989 4505 12023 4539
rect 12357 4505 12391 4539
rect 14841 4505 14875 4539
rect 14933 4505 14967 4539
rect 15853 4505 15887 4539
rect 1501 4437 1535 4471
rect 1869 4437 1903 4471
rect 3617 4437 3651 4471
rect 6285 4437 6319 4471
rect 6653 4437 6687 4471
rect 7205 4437 7239 4471
rect 9229 4437 9263 4471
rect 13553 4437 13587 4471
rect 17877 4437 17911 4471
rect 6101 4233 6135 4267
rect 6469 4233 6503 4267
rect 8033 4233 8067 4267
rect 9137 4165 9171 4199
rect 10333 4165 10367 4199
rect 11253 4165 11287 4199
rect 12541 4165 12575 4199
rect 14795 4165 14829 4199
rect 15117 4165 15151 4199
rect 1685 4097 1719 4131
rect 2513 4097 2547 4131
rect 2881 4097 2915 4131
rect 3065 4097 3099 4131
rect 3249 4097 3283 4131
rect 8493 4097 8527 4131
rect 14692 4096 14726 4130
rect 17693 4097 17727 4131
rect 17785 4097 17819 4131
rect 1869 4029 1903 4063
rect 8125 4029 8159 4063
rect 9045 4029 9079 4063
rect 10057 4029 10091 4063
rect 10241 4029 10275 4063
rect 11897 4029 11931 4063
rect 12081 4029 12115 4063
rect 12449 4029 12483 4063
rect 13461 4029 13495 4063
rect 15025 4029 15059 4063
rect 15577 4029 15611 4063
rect 2329 3961 2363 3995
rect 8861 3961 8895 3995
rect 2697 3893 2731 3927
rect 11529 3893 11563 3927
rect 14565 3893 14599 3927
rect 17969 3893 18003 3927
rect 8953 3689 8987 3723
rect 10149 3689 10183 3723
rect 15761 3689 15795 3723
rect 2789 3553 2823 3587
rect 7757 3553 7791 3587
rect 8769 3553 8803 3587
rect 14197 3553 14231 3587
rect 15025 3553 15059 3587
rect 16037 3553 16071 3587
rect 2145 3485 2179 3519
rect 2513 3485 2547 3519
rect 2697 3485 2731 3519
rect 5825 3485 5859 3519
rect 7456 3485 7490 3519
rect 9172 3485 9206 3519
rect 10920 3485 10954 3519
rect 13128 3485 13162 3519
rect 1869 3417 1903 3451
rect 5549 3417 5583 3451
rect 7849 3417 7883 3451
rect 12725 3417 12759 3451
rect 13231 3417 13265 3451
rect 14289 3417 14323 3451
rect 16129 3417 16163 3451
rect 17049 3417 17083 3451
rect 2329 3349 2363 3383
rect 7527 3349 7561 3383
rect 9275 3349 9309 3383
rect 11023 3349 11057 3383
rect 13829 3349 13863 3383
rect 5549 3077 5583 3111
rect 7849 3077 7883 3111
rect 8769 3077 8803 3111
rect 9321 3077 9355 3111
rect 10241 3077 10275 3111
rect 11713 3077 11747 3111
rect 12633 3077 12667 3111
rect 12955 3077 12989 3111
rect 13277 3077 13311 3111
rect 14381 3077 14415 3111
rect 14473 3077 14507 3111
rect 1685 3009 1719 3043
rect 2513 3009 2547 3043
rect 3341 3009 3375 3043
rect 3433 3009 3467 3043
rect 4813 3009 4847 3043
rect 5181 3009 5215 3043
rect 5825 3009 5859 3043
rect 6653 3009 6687 3043
rect 7205 3009 7239 3043
rect 7297 3009 7331 3043
rect 9229 3009 9263 3043
rect 10793 3009 10827 3043
rect 11161 3009 11195 3043
rect 12852 3009 12886 3043
rect 15485 3009 15519 3043
rect 16037 3009 16071 3043
rect 16681 3009 16715 3043
rect 17049 3009 17083 3043
rect 17417 3009 17451 3043
rect 17877 3009 17911 3043
rect 18245 3009 18279 3043
rect 1869 2941 1903 2975
rect 2697 2941 2731 2975
rect 4629 2941 4663 2975
rect 6929 2941 6963 2975
rect 7757 2941 7791 2975
rect 10333 2941 10367 2975
rect 11253 2941 11287 2975
rect 11621 2941 11655 2975
rect 13185 2941 13219 2975
rect 14013 2941 14047 2975
rect 14657 2941 14691 2975
rect 10977 2873 11011 2907
rect 15853 2873 15887 2907
rect 18061 2873 18095 2907
rect 3157 2805 3191 2839
rect 4997 2805 5031 2839
rect 5917 2805 5951 2839
rect 6469 2805 6503 2839
rect 7481 2805 7515 2839
rect 9045 2805 9079 2839
rect 10609 2805 10643 2839
rect 15669 2805 15703 2839
rect 16221 2805 16255 2839
rect 16865 2805 16899 2839
rect 17233 2805 17267 2839
rect 17601 2805 17635 2839
rect 18429 2805 18463 2839
rect 11207 2601 11241 2635
rect 14335 2601 14369 2635
rect 15485 2601 15519 2635
rect 17693 2601 17727 2635
rect 10517 2533 10551 2567
rect 14657 2533 14691 2567
rect 12909 2465 12943 2499
rect 2145 2397 2179 2431
rect 7021 2397 7055 2431
rect 7849 2397 7883 2431
rect 9229 2397 9263 2431
rect 10241 2397 10275 2431
rect 10701 2397 10735 2431
rect 11136 2397 11170 2431
rect 14232 2397 14266 2431
rect 14473 2397 14507 2431
rect 14841 2397 14875 2431
rect 17877 2397 17911 2431
rect 1869 2329 1903 2363
rect 6745 2329 6779 2363
rect 9413 2329 9447 2363
rect 11897 2329 11931 2363
rect 11989 2329 12023 2363
rect 7665 2261 7699 2295
rect 9045 2261 9079 2295
rect 10057 2261 10091 2295
rect 13001 2261 13035 2295
rect 15025 2261 15059 2295
rect 18061 2261 18095 2295
<< metal1 >>
rect 11698 15172 11704 15224
rect 11756 15212 11762 15224
rect 15470 15212 15476 15224
rect 11756 15184 15476 15212
rect 11756 15172 11762 15184
rect 15470 15172 15476 15184
rect 15528 15172 15534 15224
rect 4430 14900 4436 14952
rect 4488 14940 4494 14952
rect 11238 14940 11244 14952
rect 4488 14912 11244 14940
rect 4488 14900 4494 14912
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 8846 14832 8852 14884
rect 8904 14872 8910 14884
rect 17034 14872 17040 14884
rect 8904 14844 17040 14872
rect 8904 14832 8910 14844
rect 17034 14832 17040 14844
rect 17092 14832 17098 14884
rect 3510 14764 3516 14816
rect 3568 14804 3574 14816
rect 13354 14804 13360 14816
rect 3568 14776 13360 14804
rect 3568 14764 3574 14776
rect 13354 14764 13360 14776
rect 13412 14764 13418 14816
rect 1104 14714 18860 14736
rect 1104 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 3302 14714
rect 3354 14662 3366 14714
rect 3418 14662 3430 14714
rect 3482 14662 7622 14714
rect 7674 14662 7686 14714
rect 7738 14662 7750 14714
rect 7802 14662 7814 14714
rect 7866 14662 7878 14714
rect 7930 14662 12070 14714
rect 12122 14662 12134 14714
rect 12186 14662 12198 14714
rect 12250 14662 12262 14714
rect 12314 14662 12326 14714
rect 12378 14662 16518 14714
rect 16570 14662 16582 14714
rect 16634 14662 16646 14714
rect 16698 14662 16710 14714
rect 16762 14662 16774 14714
rect 16826 14662 18860 14714
rect 1104 14640 18860 14662
rect 2958 14560 2964 14612
rect 3016 14600 3022 14612
rect 13630 14600 13636 14612
rect 3016 14572 13636 14600
rect 3016 14560 3022 14572
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 11146 14532 11152 14544
rect 2746 14504 11152 14532
rect 2222 14424 2228 14476
rect 2280 14464 2286 14476
rect 2746 14464 2774 14504
rect 11146 14492 11152 14504
rect 11204 14492 11210 14544
rect 11238 14492 11244 14544
rect 11296 14532 11302 14544
rect 15838 14532 15844 14544
rect 11296 14504 15844 14532
rect 11296 14492 11302 14504
rect 15838 14492 15844 14504
rect 15896 14492 15902 14544
rect 2280 14436 2774 14464
rect 2280 14424 2286 14436
rect 7742 14424 7748 14476
rect 7800 14464 7806 14476
rect 17310 14464 17316 14476
rect 7800 14436 17316 14464
rect 7800 14424 7806 14436
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 1210 14356 1216 14408
rect 1268 14396 1274 14408
rect 8570 14396 8576 14408
rect 1268 14368 8576 14396
rect 1268 14356 1274 14368
rect 8570 14356 8576 14368
rect 8628 14356 8634 14408
rect 9122 14356 9128 14408
rect 9180 14396 9186 14408
rect 16390 14396 16396 14408
rect 9180 14368 16396 14396
rect 9180 14356 9186 14368
rect 16390 14356 16396 14368
rect 16448 14356 16454 14408
rect 2866 14288 2872 14340
rect 2924 14328 2930 14340
rect 9766 14328 9772 14340
rect 2924 14300 9772 14328
rect 2924 14288 2930 14300
rect 9766 14288 9772 14300
rect 9824 14288 9830 14340
rect 12434 14288 12440 14340
rect 12492 14328 12498 14340
rect 12986 14328 12992 14340
rect 12492 14300 12992 14328
rect 12492 14288 12498 14300
rect 12986 14288 12992 14300
rect 13044 14328 13050 14340
rect 18322 14328 18328 14340
rect 13044 14300 18328 14328
rect 13044 14288 13050 14300
rect 18322 14288 18328 14300
rect 18380 14288 18386 14340
rect 4798 14220 4804 14272
rect 4856 14260 4862 14272
rect 13722 14260 13728 14272
rect 4856 14232 13728 14260
rect 4856 14220 4862 14232
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 1104 14170 18860 14192
rect 1104 14118 5398 14170
rect 5450 14118 5462 14170
rect 5514 14118 5526 14170
rect 5578 14118 5590 14170
rect 5642 14118 5654 14170
rect 5706 14118 9846 14170
rect 9898 14118 9910 14170
rect 9962 14118 9974 14170
rect 10026 14118 10038 14170
rect 10090 14118 10102 14170
rect 10154 14118 14294 14170
rect 14346 14118 14358 14170
rect 14410 14118 14422 14170
rect 14474 14118 14486 14170
rect 14538 14118 14550 14170
rect 14602 14118 18860 14170
rect 1104 14096 18860 14118
rect 6546 14056 6552 14068
rect 6507 14028 6552 14056
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 6788 14028 6837 14056
rect 6788 14016 6794 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 7742 14056 7748 14068
rect 7703 14028 7748 14056
rect 6825 14019 6883 14025
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 8205 14059 8263 14065
rect 8205 14025 8217 14059
rect 8251 14025 8263 14059
rect 8570 14056 8576 14068
rect 8531 14028 8576 14056
rect 8205 14019 8263 14025
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 8220 13988 8248 14019
rect 8570 14016 8576 14028
rect 8628 14016 8634 14068
rect 8846 14056 8852 14068
rect 8807 14028 8852 14056
rect 8846 14016 8852 14028
rect 8904 14016 8910 14068
rect 9122 14056 9128 14068
rect 9083 14028 9128 14056
rect 9122 14016 9128 14028
rect 9180 14016 9186 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 9953 14059 10011 14065
rect 9953 14056 9965 14059
rect 9824 14028 9965 14056
rect 9824 14016 9830 14028
rect 9953 14025 9965 14028
rect 9999 14025 10011 14059
rect 11146 14056 11152 14068
rect 11107 14028 11152 14056
rect 9953 14019 10011 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 12618 14056 12624 14068
rect 12579 14028 12624 14056
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 13354 14056 13360 14068
rect 13315 14028 13360 14056
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 13722 14056 13728 14068
rect 13683 14028 13728 14056
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 14090 14056 14096 14068
rect 14003 14028 14096 14056
rect 14090 14016 14096 14028
rect 14148 14056 14154 14068
rect 14918 14056 14924 14068
rect 14148 14028 14924 14056
rect 14148 14016 14154 14028
rect 14918 14016 14924 14028
rect 14976 14056 14982 14068
rect 19610 14056 19616 14068
rect 14976 14028 19616 14056
rect 14976 14016 14982 14028
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 9140 13988 9168 14016
rect 11885 13991 11943 13997
rect 11885 13988 11897 13991
rect 5592 13960 8248 13988
rect 8404 13960 9168 13988
rect 11348 13960 11897 13988
rect 5592 13948 5598 13960
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 5994 13812 6000 13864
rect 6052 13852 6058 13864
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 6052 13824 6101 13852
rect 6052 13812 6058 13824
rect 6089 13821 6101 13824
rect 6135 13852 6147 13855
rect 6380 13852 6408 13883
rect 6454 13880 6460 13932
rect 6512 13920 6518 13932
rect 7009 13923 7067 13929
rect 7009 13920 7021 13923
rect 6512 13892 7021 13920
rect 6512 13880 6518 13892
rect 7009 13889 7021 13892
rect 7055 13920 7067 13923
rect 7101 13923 7159 13929
rect 7101 13920 7113 13923
rect 7055 13892 7113 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 7101 13889 7113 13892
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 7742 13920 7748 13932
rect 7607 13892 7748 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 8404 13929 8432 13960
rect 8389 13923 8447 13929
rect 8389 13889 8401 13923
rect 8435 13889 8447 13923
rect 8389 13883 8447 13889
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13920 8815 13923
rect 8846 13920 8852 13932
rect 8803 13892 8852 13920
rect 8803 13889 8815 13892
rect 8757 13883 8815 13889
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 11348 13929 11376 13960
rect 11885 13957 11897 13960
rect 11931 13988 11943 13991
rect 12434 13988 12440 14000
rect 11931 13960 12440 13988
rect 11931 13957 11943 13960
rect 11885 13951 11943 13957
rect 12434 13948 12440 13960
rect 12492 13948 12498 14000
rect 13998 13988 14004 14000
rect 12820 13960 14004 13988
rect 12820 13929 12848 13960
rect 13998 13948 14004 13960
rect 14056 13948 14062 14000
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13920 10195 13923
rect 11333 13923 11391 13929
rect 10183 13892 10364 13920
rect 10183 13889 10195 13892
rect 10137 13883 10195 13889
rect 10336 13861 10364 13892
rect 11333 13889 11345 13923
rect 11379 13889 11391 13923
rect 11333 13883 11391 13889
rect 12805 13923 12863 13929
rect 12805 13889 12817 13923
rect 12851 13889 12863 13923
rect 12805 13883 12863 13889
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13889 13599 13923
rect 13906 13920 13912 13932
rect 13819 13892 13912 13920
rect 13541 13883 13599 13889
rect 6135 13824 6408 13852
rect 10321 13855 10379 13861
rect 6135 13821 6147 13824
rect 6089 13815 6147 13821
rect 10321 13821 10333 13855
rect 10367 13852 10379 13855
rect 13170 13852 13176 13864
rect 10367 13824 13176 13852
rect 10367 13821 10379 13824
rect 10321 13815 10379 13821
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 13556 13852 13584 13883
rect 13906 13880 13912 13892
rect 13964 13920 13970 13932
rect 15102 13920 15108 13932
rect 13964 13892 15108 13920
rect 13964 13880 13970 13892
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15197 13923 15255 13929
rect 15197 13889 15209 13923
rect 15243 13920 15255 13923
rect 15470 13920 15476 13932
rect 15243 13892 15476 13920
rect 15243 13889 15255 13892
rect 15197 13883 15255 13889
rect 15470 13880 15476 13892
rect 15528 13920 15534 13932
rect 15746 13920 15752 13932
rect 15528 13892 15752 13920
rect 15528 13880 15534 13892
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 14090 13852 14096 13864
rect 13556 13824 14096 13852
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 1578 13744 1584 13796
rect 1636 13784 1642 13796
rect 7377 13787 7435 13793
rect 7377 13784 7389 13787
rect 1636 13756 7389 13784
rect 1636 13744 1642 13756
rect 7377 13753 7389 13756
rect 7423 13753 7435 13787
rect 7377 13747 7435 13753
rect 290 13676 296 13728
rect 348 13716 354 13728
rect 5534 13716 5540 13728
rect 348 13688 5540 13716
rect 348 13676 354 13688
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 11606 13716 11612 13728
rect 6420 13688 11612 13716
rect 6420 13676 6426 13688
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 15010 13716 15016 13728
rect 14971 13688 15016 13716
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 1104 13626 18860 13648
rect 1104 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 3302 13626
rect 3354 13574 3366 13626
rect 3418 13574 3430 13626
rect 3482 13574 7622 13626
rect 7674 13574 7686 13626
rect 7738 13574 7750 13626
rect 7802 13574 7814 13626
rect 7866 13574 7878 13626
rect 7930 13574 12070 13626
rect 12122 13574 12134 13626
rect 12186 13574 12198 13626
rect 12250 13574 12262 13626
rect 12314 13574 12326 13626
rect 12378 13574 16518 13626
rect 16570 13574 16582 13626
rect 16634 13574 16646 13626
rect 16698 13574 16710 13626
rect 16762 13574 16774 13626
rect 16826 13574 18860 13626
rect 1104 13552 18860 13574
rect 11606 13472 11612 13524
rect 11664 13512 11670 13524
rect 12158 13512 12164 13524
rect 11664 13484 12164 13512
rect 11664 13472 11670 13484
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 6822 13444 6828 13456
rect 6472 13416 6828 13444
rect 5813 13379 5871 13385
rect 5813 13345 5825 13379
rect 5859 13376 5871 13379
rect 5902 13376 5908 13388
rect 5859 13348 5908 13376
rect 5859 13345 5871 13348
rect 5813 13339 5871 13345
rect 5902 13336 5908 13348
rect 5960 13336 5966 13388
rect 6472 13385 6500 13416
rect 6822 13404 6828 13416
rect 6880 13444 6886 13456
rect 6880 13416 13032 13444
rect 6880 13404 6886 13416
rect 6457 13379 6515 13385
rect 6457 13345 6469 13379
rect 6503 13345 6515 13379
rect 6457 13339 6515 13345
rect 6641 13379 6699 13385
rect 6641 13345 6653 13379
rect 6687 13376 6699 13379
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 6687 13348 7481 13376
rect 6687 13345 6699 13348
rect 6641 13339 6699 13345
rect 7469 13345 7481 13348
rect 7515 13376 7527 13379
rect 8202 13376 8208 13388
rect 7515 13348 8208 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 9769 13379 9827 13385
rect 9769 13376 9781 13379
rect 9456 13348 9781 13376
rect 9456 13336 9462 13348
rect 9769 13345 9781 13348
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 11609 13379 11667 13385
rect 11609 13345 11621 13379
rect 11655 13376 11667 13379
rect 11974 13376 11980 13388
rect 11655 13348 11980 13376
rect 11655 13345 11667 13348
rect 11609 13339 11667 13345
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 12268 13385 12296 13416
rect 12253 13379 12311 13385
rect 12253 13345 12265 13379
rect 12299 13345 12311 13379
rect 12253 13339 12311 13345
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 12492 13348 12537 13376
rect 12492 13336 12498 13348
rect 2866 13268 2872 13320
rect 2924 13308 2930 13320
rect 7285 13311 7343 13317
rect 7285 13308 7297 13311
rect 2924 13280 7297 13308
rect 2924 13268 2930 13280
rect 7285 13277 7297 13280
rect 7331 13308 7343 13311
rect 7745 13311 7803 13317
rect 7745 13308 7757 13311
rect 7331 13280 7757 13308
rect 7331 13277 7343 13280
rect 7285 13271 7343 13277
rect 7745 13277 7757 13280
rect 7791 13308 7803 13311
rect 12066 13308 12072 13320
rect 7791 13280 12072 13308
rect 7791 13277 7803 13280
rect 7745 13271 7803 13277
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 13004 13317 13032 13416
rect 13262 13336 13268 13388
rect 13320 13376 13326 13388
rect 15286 13376 15292 13388
rect 13320 13348 15292 13376
rect 13320 13336 13326 13348
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 12989 13311 13047 13317
rect 12216 13280 12261 13308
rect 12216 13268 12222 13280
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 15194 13308 15200 13320
rect 13035 13280 15200 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 15194 13268 15200 13280
rect 15252 13268 15258 13320
rect 3970 13200 3976 13252
rect 4028 13240 4034 13252
rect 5258 13240 5264 13252
rect 4028 13212 5264 13240
rect 4028 13200 4034 13212
rect 5258 13200 5264 13212
rect 5316 13200 5322 13252
rect 5537 13243 5595 13249
rect 5537 13209 5549 13243
rect 5583 13240 5595 13243
rect 5583 13212 6868 13240
rect 5583 13209 5595 13212
rect 5537 13203 5595 13209
rect 5166 13172 5172 13184
rect 5127 13144 5172 13172
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 5629 13175 5687 13181
rect 5629 13141 5641 13175
rect 5675 13172 5687 13175
rect 5997 13175 6055 13181
rect 5997 13172 6009 13175
rect 5675 13144 6009 13172
rect 5675 13141 5687 13144
rect 5629 13135 5687 13141
rect 5997 13141 6009 13144
rect 6043 13141 6055 13175
rect 6362 13172 6368 13184
rect 6323 13144 6368 13172
rect 5997 13135 6055 13141
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 6840 13181 6868 13212
rect 7006 13200 7012 13252
rect 7064 13240 7070 13252
rect 9677 13243 9735 13249
rect 9677 13240 9689 13243
rect 7064 13212 9689 13240
rect 7064 13200 7070 13212
rect 9677 13209 9689 13212
rect 9723 13240 9735 13243
rect 10045 13243 10103 13249
rect 10045 13240 10057 13243
rect 9723 13212 10057 13240
rect 9723 13209 9735 13212
rect 9677 13203 9735 13209
rect 10045 13209 10057 13212
rect 10091 13240 10103 13243
rect 16022 13240 16028 13252
rect 10091 13212 16028 13240
rect 10091 13209 10103 13212
rect 10045 13203 10103 13209
rect 16022 13200 16028 13212
rect 16080 13200 16086 13252
rect 6825 13175 6883 13181
rect 6825 13141 6837 13175
rect 6871 13141 6883 13175
rect 7190 13172 7196 13184
rect 7151 13144 7196 13172
rect 6825 13135 6883 13141
rect 7190 13132 7196 13144
rect 7248 13132 7254 13184
rect 8294 13132 8300 13184
rect 8352 13172 8358 13184
rect 9217 13175 9275 13181
rect 9217 13172 9229 13175
rect 8352 13144 9229 13172
rect 8352 13132 8358 13144
rect 9217 13141 9229 13144
rect 9263 13141 9275 13175
rect 9582 13172 9588 13184
rect 9543 13144 9588 13172
rect 9217 13135 9275 13141
rect 9582 13132 9588 13144
rect 9640 13132 9646 13184
rect 10965 13175 11023 13181
rect 10965 13141 10977 13175
rect 11011 13172 11023 13175
rect 11146 13172 11152 13184
rect 11011 13144 11152 13172
rect 11011 13141 11023 13144
rect 10965 13135 11023 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 11330 13172 11336 13184
rect 11291 13144 11336 13172
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 11425 13175 11483 13181
rect 11425 13141 11437 13175
rect 11471 13172 11483 13175
rect 11793 13175 11851 13181
rect 11793 13172 11805 13175
rect 11471 13144 11805 13172
rect 11471 13141 11483 13144
rect 11425 13135 11483 13141
rect 11793 13141 11805 13144
rect 11839 13141 11851 13175
rect 12618 13172 12624 13184
rect 12579 13144 12624 13172
rect 11793 13135 11851 13141
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 13814 13172 13820 13184
rect 13775 13144 13820 13172
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 1104 13082 18860 13104
rect 1104 13030 5398 13082
rect 5450 13030 5462 13082
rect 5514 13030 5526 13082
rect 5578 13030 5590 13082
rect 5642 13030 5654 13082
rect 5706 13030 9846 13082
rect 9898 13030 9910 13082
rect 9962 13030 9974 13082
rect 10026 13030 10038 13082
rect 10090 13030 10102 13082
rect 10154 13030 14294 13082
rect 14346 13030 14358 13082
rect 14410 13030 14422 13082
rect 14474 13030 14486 13082
rect 14538 13030 14550 13082
rect 14602 13030 18860 13082
rect 1104 13008 18860 13030
rect 2777 12971 2835 12977
rect 2777 12937 2789 12971
rect 2823 12968 2835 12971
rect 2866 12968 2872 12980
rect 2823 12940 2872 12968
rect 2823 12937 2835 12940
rect 2777 12931 2835 12937
rect 2792 12900 2820 12931
rect 2866 12928 2872 12940
rect 2924 12928 2930 12980
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 3329 12971 3387 12977
rect 3329 12968 3341 12971
rect 3108 12940 3341 12968
rect 3108 12928 3114 12940
rect 3329 12937 3341 12940
rect 3375 12968 3387 12971
rect 3878 12968 3884 12980
rect 3375 12940 3884 12968
rect 3375 12937 3387 12940
rect 3329 12931 3387 12937
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 3973 12971 4031 12977
rect 3973 12937 3985 12971
rect 4019 12968 4031 12971
rect 4430 12968 4436 12980
rect 4019 12940 4436 12968
rect 4019 12937 4031 12940
rect 3973 12931 4031 12937
rect 2056 12872 2820 12900
rect 2056 12841 2084 12872
rect 2958 12860 2964 12912
rect 3016 12900 3022 12912
rect 3988 12900 4016 12931
rect 4430 12928 4436 12940
rect 4488 12928 4494 12980
rect 5166 12968 5172 12980
rect 5127 12940 5172 12968
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 5258 12928 5264 12980
rect 5316 12968 5322 12980
rect 5813 12971 5871 12977
rect 5813 12968 5825 12971
rect 5316 12940 5825 12968
rect 5316 12928 5322 12940
rect 5813 12937 5825 12940
rect 5859 12968 5871 12971
rect 6362 12968 6368 12980
rect 5859 12940 6368 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 6362 12928 6368 12940
rect 6420 12928 6426 12980
rect 6549 12971 6607 12977
rect 6549 12937 6561 12971
rect 6595 12968 6607 12971
rect 7190 12968 7196 12980
rect 6595 12940 7196 12968
rect 6595 12937 6607 12940
rect 6549 12931 6607 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 9217 12971 9275 12977
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 9585 12971 9643 12977
rect 9585 12968 9597 12971
rect 9263 12940 9597 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 9585 12937 9597 12940
rect 9631 12937 9643 12971
rect 9585 12931 9643 12937
rect 10226 12928 10232 12980
rect 10284 12968 10290 12980
rect 11146 12968 11152 12980
rect 10284 12940 11152 12968
rect 10284 12928 10290 12940
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 11609 12971 11667 12977
rect 11609 12968 11621 12971
rect 11388 12940 11621 12968
rect 11388 12928 11394 12940
rect 11609 12937 11621 12940
rect 11655 12937 11667 12971
rect 11609 12931 11667 12937
rect 11977 12971 12035 12977
rect 11977 12937 11989 12971
rect 12023 12968 12035 12971
rect 12618 12968 12624 12980
rect 12023 12940 12624 12968
rect 12023 12937 12035 12940
rect 11977 12931 12035 12937
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 13541 12971 13599 12977
rect 13541 12937 13553 12971
rect 13587 12968 13599 12971
rect 13909 12971 13967 12977
rect 13909 12968 13921 12971
rect 13587 12940 13921 12968
rect 13587 12937 13599 12940
rect 13541 12931 13599 12937
rect 13909 12937 13921 12940
rect 13955 12937 13967 12971
rect 13909 12931 13967 12937
rect 3016 12872 4016 12900
rect 3016 12860 3022 12872
rect 4062 12860 4068 12912
rect 4120 12900 4126 12912
rect 6270 12900 6276 12912
rect 4120 12872 6276 12900
rect 4120 12860 4126 12872
rect 6270 12860 6276 12872
rect 6328 12860 6334 12912
rect 6825 12903 6883 12909
rect 6825 12869 6837 12903
rect 6871 12900 6883 12903
rect 8665 12903 8723 12909
rect 8665 12900 8677 12903
rect 6871 12872 8677 12900
rect 6871 12869 6883 12872
rect 6825 12863 6883 12869
rect 7208 12844 7236 12872
rect 8665 12869 8677 12872
rect 8711 12900 8723 12903
rect 10045 12903 10103 12909
rect 10045 12900 10057 12903
rect 8711 12872 10057 12900
rect 8711 12869 8723 12872
rect 8665 12863 8723 12869
rect 10045 12869 10057 12872
rect 10091 12900 10103 12903
rect 12066 12900 12072 12912
rect 10091 12872 10640 12900
rect 11979 12872 12072 12900
rect 10091 12869 10103 12872
rect 10045 12863 10103 12869
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12801 2099 12835
rect 2041 12795 2099 12801
rect 2409 12835 2467 12841
rect 2409 12801 2421 12835
rect 2455 12801 2467 12835
rect 2409 12795 2467 12801
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12832 5319 12835
rect 6638 12832 6644 12844
rect 5307 12804 6644 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 2424 12764 2452 12795
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 7190 12792 7196 12844
rect 7248 12792 7254 12844
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12832 9183 12835
rect 9674 12832 9680 12844
rect 9171 12804 9680 12832
rect 9171 12801 9183 12804
rect 9125 12795 9183 12801
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 9953 12835 10011 12841
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10612 12832 10640 12872
rect 12066 12860 12072 12872
rect 12124 12900 12130 12912
rect 12529 12903 12587 12909
rect 12529 12900 12541 12903
rect 12124 12872 12541 12900
rect 12124 12860 12130 12872
rect 12529 12869 12541 12872
rect 12575 12900 12587 12903
rect 13262 12900 13268 12912
rect 12575 12872 13268 12900
rect 12575 12869 12587 12872
rect 12529 12863 12587 12869
rect 13262 12860 13268 12872
rect 13320 12860 13326 12912
rect 13814 12900 13820 12912
rect 13372 12872 13820 12900
rect 13372 12832 13400 12872
rect 13814 12860 13820 12872
rect 13872 12900 13878 12912
rect 14369 12903 14427 12909
rect 14369 12900 14381 12903
rect 13872 12872 14381 12900
rect 13872 12860 13878 12872
rect 14369 12869 14381 12872
rect 14415 12900 14427 12903
rect 15654 12900 15660 12912
rect 14415 12872 15660 12900
rect 14415 12869 14427 12872
rect 14369 12863 14427 12869
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 9999 12804 10548 12832
rect 10612 12804 13400 12832
rect 13449 12835 13507 12841
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 2424 12736 2605 12764
rect 2593 12733 2605 12736
rect 2639 12764 2651 12767
rect 2639 12736 4016 12764
rect 2639 12733 2651 12736
rect 2593 12727 2651 12733
rect 1857 12699 1915 12705
rect 1857 12665 1869 12699
rect 1903 12696 1915 12699
rect 2866 12696 2872 12708
rect 1903 12668 2872 12696
rect 1903 12665 1915 12668
rect 1857 12659 1915 12665
rect 2866 12656 2872 12668
rect 2924 12656 2930 12708
rect 3988 12696 4016 12736
rect 4062 12724 4068 12776
rect 4120 12764 4126 12776
rect 4120 12736 4165 12764
rect 4908 12736 5304 12764
rect 4120 12724 4126 12736
rect 4908 12696 4936 12736
rect 3988 12668 4936 12696
rect 5276 12696 5304 12736
rect 5350 12724 5356 12776
rect 5408 12764 5414 12776
rect 5408 12736 5453 12764
rect 5408 12724 5414 12736
rect 6362 12724 6368 12776
rect 6420 12764 6426 12776
rect 6822 12764 6828 12776
rect 6420 12736 6828 12764
rect 6420 12724 6426 12736
rect 6822 12724 6828 12736
rect 6880 12764 6886 12776
rect 6917 12767 6975 12773
rect 6917 12764 6929 12767
rect 6880 12736 6929 12764
rect 6880 12724 6886 12736
rect 6917 12733 6929 12736
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 8202 12724 8208 12776
rect 8260 12764 8266 12776
rect 9309 12767 9367 12773
rect 9309 12764 9321 12767
rect 8260 12736 9321 12764
rect 8260 12724 8266 12736
rect 9309 12733 9321 12736
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 9490 12724 9496 12776
rect 9548 12764 9554 12776
rect 9968 12764 9996 12795
rect 10226 12764 10232 12776
rect 9548 12736 9996 12764
rect 10187 12736 10232 12764
rect 9548 12724 9554 12736
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 10520 12708 10548 12804
rect 13449 12801 13461 12835
rect 13495 12832 13507 12835
rect 14090 12832 14096 12844
rect 13495 12804 14096 12832
rect 13495 12801 13507 12804
rect 13449 12795 13507 12801
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 14274 12832 14280 12844
rect 14235 12804 14280 12832
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12764 12311 12767
rect 12434 12764 12440 12776
rect 12299 12736 12440 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12434 12724 12440 12736
rect 12492 12764 12498 12776
rect 13354 12764 13360 12776
rect 12492 12736 13360 12764
rect 12492 12724 12498 12736
rect 13354 12724 13360 12736
rect 13412 12764 13418 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 13412 12736 13645 12764
rect 13412 12724 13418 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 14458 12724 14464 12776
rect 14516 12764 14522 12776
rect 14516 12736 14561 12764
rect 14516 12724 14522 12736
rect 7006 12696 7012 12708
rect 5276 12668 7012 12696
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 7098 12656 7104 12708
rect 7156 12696 7162 12708
rect 8757 12699 8815 12705
rect 8757 12696 8769 12699
rect 7156 12668 8769 12696
rect 7156 12656 7162 12668
rect 8757 12665 8769 12668
rect 8803 12665 8815 12699
rect 10502 12696 10508 12708
rect 10463 12668 10508 12696
rect 8757 12659 8815 12665
rect 10502 12656 10508 12668
rect 10560 12656 10566 12708
rect 12158 12656 12164 12708
rect 12216 12696 12222 12708
rect 17862 12696 17868 12708
rect 12216 12668 17868 12696
rect 12216 12656 12222 12668
rect 17862 12656 17868 12668
rect 17920 12656 17926 12708
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 2225 12631 2283 12637
rect 2225 12628 2237 12631
rect 2096 12600 2237 12628
rect 2096 12588 2102 12600
rect 2225 12597 2237 12600
rect 2271 12597 2283 12631
rect 3510 12628 3516 12640
rect 3471 12600 3516 12628
rect 2225 12591 2283 12597
rect 3510 12588 3516 12600
rect 3568 12588 3574 12640
rect 4798 12628 4804 12640
rect 4759 12600 4804 12628
rect 4798 12588 4804 12600
rect 4856 12588 4862 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12618 12628 12624 12640
rect 11848 12600 12624 12628
rect 11848 12588 11854 12600
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 13078 12628 13084 12640
rect 13039 12600 13084 12628
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 14274 12588 14280 12640
rect 14332 12628 14338 12640
rect 14829 12631 14887 12637
rect 14829 12628 14841 12631
rect 14332 12600 14841 12628
rect 14332 12588 14338 12600
rect 14829 12597 14841 12600
rect 14875 12628 14887 12631
rect 16390 12628 16396 12640
rect 14875 12600 16396 12628
rect 14875 12597 14887 12600
rect 14829 12591 14887 12597
rect 16390 12588 16396 12600
rect 16448 12588 16454 12640
rect 1104 12538 18860 12560
rect 1104 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 3302 12538
rect 3354 12486 3366 12538
rect 3418 12486 3430 12538
rect 3482 12486 7622 12538
rect 7674 12486 7686 12538
rect 7738 12486 7750 12538
rect 7802 12486 7814 12538
rect 7866 12486 7878 12538
rect 7930 12486 12070 12538
rect 12122 12486 12134 12538
rect 12186 12486 12198 12538
rect 12250 12486 12262 12538
rect 12314 12486 12326 12538
rect 12378 12486 16518 12538
rect 16570 12486 16582 12538
rect 16634 12486 16646 12538
rect 16698 12486 16710 12538
rect 16762 12486 16774 12538
rect 16826 12486 18860 12538
rect 1104 12464 18860 12486
rect 2225 12427 2283 12433
rect 2225 12393 2237 12427
rect 2271 12424 2283 12427
rect 2958 12424 2964 12436
rect 2271 12396 2964 12424
rect 2271 12393 2283 12396
rect 2225 12387 2283 12393
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12220 2099 12223
rect 2240 12220 2268 12387
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 9490 12424 9496 12436
rect 7340 12396 9496 12424
rect 7340 12384 7346 12396
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 11698 12384 11704 12436
rect 11756 12384 11762 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 13817 12427 13875 12433
rect 13817 12424 13829 12427
rect 12492 12396 13829 12424
rect 12492 12384 12498 12396
rect 13817 12393 13829 12396
rect 13863 12393 13875 12427
rect 14090 12424 14096 12436
rect 14051 12396 14096 12424
rect 13817 12387 13875 12393
rect 2682 12316 2688 12368
rect 2740 12356 2746 12368
rect 3142 12356 3148 12368
rect 2740 12328 3148 12356
rect 2740 12316 2746 12328
rect 3142 12316 3148 12328
rect 3200 12356 3206 12368
rect 4157 12359 4215 12365
rect 4157 12356 4169 12359
rect 3200 12328 4169 12356
rect 3200 12316 3206 12328
rect 4157 12325 4169 12328
rect 4203 12356 4215 12359
rect 11716 12356 11744 12384
rect 4203 12328 11744 12356
rect 4203 12325 4215 12328
rect 4157 12319 4215 12325
rect 12710 12316 12716 12368
rect 12768 12356 12774 12368
rect 13630 12356 13636 12368
rect 12768 12328 13636 12356
rect 12768 12316 12774 12328
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 3053 12291 3111 12297
rect 3053 12257 3065 12291
rect 3099 12288 3111 12291
rect 4062 12288 4068 12300
rect 3099 12260 4068 12288
rect 3099 12257 3111 12260
rect 3053 12251 3111 12257
rect 4062 12248 4068 12260
rect 4120 12288 4126 12300
rect 4985 12291 5043 12297
rect 4985 12288 4997 12291
rect 4120 12260 4997 12288
rect 4120 12248 4126 12260
rect 4985 12257 4997 12260
rect 5031 12288 5043 12291
rect 6546 12288 6552 12300
rect 5031 12260 6552 12288
rect 5031 12257 5043 12260
rect 4985 12251 5043 12257
rect 6546 12248 6552 12260
rect 6604 12288 6610 12300
rect 6641 12291 6699 12297
rect 6641 12288 6653 12291
rect 6604 12260 6653 12288
rect 6604 12248 6610 12260
rect 6641 12257 6653 12260
rect 6687 12257 6699 12291
rect 6641 12251 6699 12257
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 7432 12260 7481 12288
rect 7432 12248 7438 12260
rect 7469 12257 7481 12260
rect 7515 12288 7527 12291
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 7515 12260 8309 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 8297 12257 8309 12260
rect 8343 12257 8355 12291
rect 9582 12288 9588 12300
rect 9543 12260 9588 12288
rect 8297 12251 8355 12257
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 10226 12288 10232 12300
rect 10187 12260 10232 12288
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 11517 12291 11575 12297
rect 11517 12257 11529 12291
rect 11563 12288 11575 12291
rect 11606 12288 11612 12300
rect 11563 12260 11612 12288
rect 11563 12257 11575 12260
rect 11517 12251 11575 12257
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 11974 12288 11980 12300
rect 11756 12260 11980 12288
rect 11756 12248 11762 12260
rect 11974 12248 11980 12260
rect 12032 12288 12038 12300
rect 12529 12291 12587 12297
rect 12529 12288 12541 12291
rect 12032 12260 12541 12288
rect 12032 12248 12038 12260
rect 12529 12257 12541 12260
rect 12575 12257 12587 12291
rect 12529 12251 12587 12257
rect 12618 12248 12624 12300
rect 12676 12288 12682 12300
rect 13354 12288 13360 12300
rect 12676 12260 13216 12288
rect 13315 12260 13360 12288
rect 12676 12248 12682 12260
rect 3694 12220 3700 12232
rect 2087 12192 2268 12220
rect 2746 12192 3700 12220
rect 2087 12189 2099 12192
rect 2041 12183 2099 12189
rect 1857 12087 1915 12093
rect 1857 12053 1869 12087
rect 1903 12084 1915 12087
rect 2746 12084 2774 12192
rect 3694 12180 3700 12192
rect 3752 12180 3758 12232
rect 7282 12220 7288 12232
rect 7243 12192 7288 12220
rect 7282 12180 7288 12192
rect 7340 12180 7346 12232
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 8205 12223 8263 12229
rect 8205 12220 8217 12223
rect 7616 12192 8217 12220
rect 7616 12180 7622 12192
rect 8205 12189 8217 12192
rect 8251 12220 8263 12223
rect 9217 12223 9275 12229
rect 9217 12220 9229 12223
rect 8251 12192 9229 12220
rect 8251 12189 8263 12192
rect 8205 12183 8263 12189
rect 9217 12189 9229 12192
rect 9263 12220 9275 12223
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9263 12192 10149 12220
rect 9263 12189 9275 12192
rect 9217 12183 9275 12189
rect 10137 12189 10149 12192
rect 10183 12220 10195 12223
rect 10410 12220 10416 12232
rect 10183 12192 10416 12220
rect 10183 12189 10195 12192
rect 10137 12183 10195 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 11238 12220 11244 12232
rect 11199 12192 11244 12220
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12220 12495 12223
rect 13078 12220 13084 12232
rect 12483 12192 13084 12220
rect 12483 12189 12495 12192
rect 12437 12183 12495 12189
rect 13078 12180 13084 12192
rect 13136 12180 13142 12232
rect 13188 12229 13216 12260
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12220 13231 12223
rect 13538 12220 13544 12232
rect 13219 12192 13544 12220
rect 13219 12189 13231 12192
rect 13173 12183 13231 12189
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 13832 12220 13860 12387
rect 14090 12384 14096 12396
rect 14148 12384 14154 12436
rect 14642 12288 14648 12300
rect 14603 12260 14648 12288
rect 14642 12248 14648 12260
rect 14700 12248 14706 12300
rect 15194 12288 15200 12300
rect 15155 12260 15200 12288
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 15838 12248 15844 12300
rect 15896 12288 15902 12300
rect 16114 12288 16120 12300
rect 15896 12260 16120 12288
rect 15896 12248 15902 12260
rect 16114 12248 16120 12260
rect 16172 12248 16178 12300
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 13832 12192 14565 12220
rect 14553 12189 14565 12192
rect 14599 12220 14611 12223
rect 16758 12220 16764 12232
rect 14599 12192 16764 12220
rect 14599 12189 14611 12192
rect 14553 12183 14611 12189
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12220 17739 12223
rect 17773 12223 17831 12229
rect 17773 12220 17785 12223
rect 17727 12192 17785 12220
rect 17727 12189 17739 12192
rect 17681 12183 17739 12189
rect 17773 12189 17785 12192
rect 17819 12189 17831 12223
rect 17773 12183 17831 12189
rect 3142 12152 3148 12164
rect 3103 12124 3148 12152
rect 3142 12112 3148 12124
rect 3200 12112 3206 12164
rect 3237 12155 3295 12161
rect 3237 12121 3249 12155
rect 3283 12152 3295 12155
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 3283 12124 3801 12152
rect 3283 12121 3295 12124
rect 3237 12115 3295 12121
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 3789 12115 3847 12121
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 4249 12155 4307 12161
rect 4249 12152 4261 12155
rect 4212 12124 4261 12152
rect 4212 12112 4218 12124
rect 4249 12121 4261 12124
rect 4295 12152 4307 12155
rect 4801 12155 4859 12161
rect 4801 12152 4813 12155
rect 4295 12124 4813 12152
rect 4295 12121 4307 12124
rect 4249 12115 4307 12121
rect 4801 12121 4813 12124
rect 4847 12152 4859 12155
rect 5166 12152 5172 12164
rect 4847 12124 5172 12152
rect 4847 12121 4859 12124
rect 4801 12115 4859 12121
rect 5166 12112 5172 12124
rect 5224 12112 5230 12164
rect 6457 12155 6515 12161
rect 6457 12121 6469 12155
rect 6503 12152 6515 12155
rect 6503 12124 7788 12152
rect 6503 12121 6515 12124
rect 6457 12115 6515 12121
rect 1903 12056 2774 12084
rect 1903 12053 1915 12056
rect 1857 12047 1915 12053
rect 3326 12044 3332 12096
rect 3384 12084 3390 12096
rect 3605 12087 3663 12093
rect 3605 12084 3617 12087
rect 3384 12056 3617 12084
rect 3384 12044 3390 12056
rect 3605 12053 3617 12056
rect 3651 12053 3663 12087
rect 3605 12047 3663 12053
rect 4338 12044 4344 12096
rect 4396 12084 4402 12096
rect 4433 12087 4491 12093
rect 4433 12084 4445 12087
rect 4396 12056 4445 12084
rect 4396 12044 4402 12056
rect 4433 12053 4445 12056
rect 4479 12053 4491 12087
rect 4433 12047 4491 12053
rect 4890 12044 4896 12096
rect 4948 12084 4954 12096
rect 6086 12084 6092 12096
rect 4948 12056 4993 12084
rect 6047 12056 6092 12084
rect 4948 12044 4954 12056
rect 6086 12044 6092 12056
rect 6144 12044 6150 12096
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 6595 12056 6929 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 6917 12053 6929 12056
rect 6963 12053 6975 12087
rect 6917 12047 6975 12053
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 7760 12093 7788 12124
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 12345 12155 12403 12161
rect 9456 12124 12112 12152
rect 9456 12112 9462 12124
rect 7377 12087 7435 12093
rect 7377 12084 7389 12087
rect 7248 12056 7389 12084
rect 7248 12044 7254 12056
rect 7377 12053 7389 12056
rect 7423 12053 7435 12087
rect 7377 12047 7435 12053
rect 7745 12087 7803 12093
rect 7745 12053 7757 12087
rect 7791 12053 7803 12087
rect 8110 12084 8116 12096
rect 8071 12056 8116 12084
rect 7745 12047 7803 12053
rect 8110 12044 8116 12056
rect 8168 12084 8174 12096
rect 8573 12087 8631 12093
rect 8573 12084 8585 12087
rect 8168 12056 8585 12084
rect 8168 12044 8174 12056
rect 8573 12053 8585 12056
rect 8619 12084 8631 12087
rect 10045 12087 10103 12093
rect 10045 12084 10057 12087
rect 8619 12056 10057 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 10045 12053 10057 12056
rect 10091 12084 10103 12087
rect 10502 12084 10508 12096
rect 10091 12056 10508 12084
rect 10091 12053 10103 12056
rect 10045 12047 10103 12053
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 10870 12084 10876 12096
rect 10831 12056 10876 12084
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 11333 12087 11391 12093
rect 11333 12053 11345 12087
rect 11379 12084 11391 12087
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11379 12056 11989 12084
rect 11379 12053 11391 12056
rect 11333 12047 11391 12053
rect 11977 12053 11989 12056
rect 12023 12053 12035 12087
rect 12084 12084 12112 12124
rect 12345 12121 12357 12155
rect 12391 12152 12403 12155
rect 12391 12124 12848 12152
rect 12391 12121 12403 12124
rect 12345 12115 12403 12121
rect 12710 12084 12716 12096
rect 12084 12056 12716 12084
rect 11977 12047 12035 12053
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 12820 12093 12848 12124
rect 12894 12112 12900 12164
rect 12952 12152 12958 12164
rect 17696 12152 17724 12183
rect 12952 12124 17724 12152
rect 12952 12112 12958 12124
rect 12805 12087 12863 12093
rect 12805 12053 12817 12087
rect 12851 12053 12863 12087
rect 12805 12047 12863 12053
rect 13262 12044 13268 12096
rect 13320 12084 13326 12096
rect 13320 12056 13365 12084
rect 13320 12044 13326 12056
rect 14090 12044 14096 12096
rect 14148 12084 14154 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 14148 12056 14473 12084
rect 14148 12044 14154 12056
rect 14461 12053 14473 12056
rect 14507 12084 14519 12087
rect 15381 12087 15439 12093
rect 15381 12084 15393 12087
rect 14507 12056 15393 12084
rect 14507 12053 14519 12056
rect 14461 12047 14519 12053
rect 15381 12053 15393 12056
rect 15427 12084 15439 12087
rect 15838 12084 15844 12096
rect 15427 12056 15844 12084
rect 15427 12053 15439 12056
rect 15381 12047 15439 12053
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 17957 12087 18015 12093
rect 17957 12053 17969 12087
rect 18003 12084 18015 12087
rect 18598 12084 18604 12096
rect 18003 12056 18604 12084
rect 18003 12053 18015 12056
rect 17957 12047 18015 12053
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 1104 11994 18860 12016
rect 1104 11942 5398 11994
rect 5450 11942 5462 11994
rect 5514 11942 5526 11994
rect 5578 11942 5590 11994
rect 5642 11942 5654 11994
rect 5706 11942 9846 11994
rect 9898 11942 9910 11994
rect 9962 11942 9974 11994
rect 10026 11942 10038 11994
rect 10090 11942 10102 11994
rect 10154 11942 14294 11994
rect 14346 11942 14358 11994
rect 14410 11942 14422 11994
rect 14474 11942 14486 11994
rect 14538 11942 14550 11994
rect 14602 11942 18860 11994
rect 1104 11920 18860 11942
rect 2682 11880 2688 11892
rect 2643 11852 2688 11880
rect 2682 11840 2688 11852
rect 2740 11840 2746 11892
rect 2958 11880 2964 11892
rect 2919 11852 2964 11880
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 3326 11880 3332 11892
rect 3287 11852 3332 11880
rect 3326 11840 3332 11852
rect 3384 11840 3390 11892
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 3510 11880 3516 11892
rect 3467 11852 3516 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 4338 11880 4344 11892
rect 4299 11852 4344 11880
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 4890 11840 4896 11892
rect 4948 11880 4954 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 4948 11852 5457 11880
rect 4948 11840 4954 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 5445 11843 5503 11849
rect 5813 11883 5871 11889
rect 5813 11849 5825 11883
rect 5859 11880 5871 11883
rect 6454 11880 6460 11892
rect 5859 11852 6460 11880
rect 5859 11849 5871 11852
rect 5813 11843 5871 11849
rect 6454 11840 6460 11852
rect 6512 11840 6518 11892
rect 6638 11880 6644 11892
rect 6599 11852 6644 11880
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 7098 11880 7104 11892
rect 7059 11852 7104 11880
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 8294 11880 8300 11892
rect 8255 11852 8300 11880
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 8404 11852 8616 11880
rect 2700 11812 2728 11840
rect 2056 11784 2728 11812
rect 4433 11815 4491 11821
rect 2056 11753 2084 11784
rect 4433 11781 4445 11815
rect 4479 11812 4491 11815
rect 6086 11812 6092 11824
rect 4479 11784 6092 11812
rect 4479 11781 4491 11784
rect 4433 11775 4491 11781
rect 6086 11772 6092 11784
rect 6144 11772 6150 11824
rect 8404 11812 8432 11852
rect 6840 11784 8432 11812
rect 8588 11812 8616 11852
rect 10410 11840 10416 11892
rect 10468 11880 10474 11892
rect 12434 11880 12440 11892
rect 10468 11852 12440 11880
rect 10468 11840 10474 11852
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12621 11883 12679 11889
rect 12621 11849 12633 11883
rect 12667 11880 12679 11883
rect 12894 11880 12900 11892
rect 12667 11852 12900 11880
rect 12667 11849 12679 11852
rect 12621 11843 12679 11849
rect 12161 11815 12219 11821
rect 12161 11812 12173 11815
rect 8588 11784 12173 11812
rect 2041 11747 2099 11753
rect 2041 11713 2053 11747
rect 2087 11713 2099 11747
rect 2041 11707 2099 11713
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2498 11744 2504 11756
rect 2455 11716 2504 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 2866 11704 2872 11756
rect 2924 11744 2930 11756
rect 3786 11744 3792 11756
rect 2924 11716 3792 11744
rect 2924 11704 2930 11716
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 4062 11704 4068 11756
rect 4120 11744 4126 11756
rect 5261 11747 5319 11753
rect 5261 11744 5273 11747
rect 4120 11716 5273 11744
rect 4120 11704 4126 11716
rect 5261 11713 5273 11716
rect 5307 11744 5319 11747
rect 6840 11744 6868 11784
rect 12161 11781 12173 11784
rect 12207 11812 12219 11815
rect 12636 11812 12664 11843
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 13081 11883 13139 11889
rect 13081 11849 13093 11883
rect 13127 11880 13139 11883
rect 13262 11880 13268 11892
rect 13127 11852 13268 11880
rect 13127 11849 13139 11852
rect 13081 11843 13139 11849
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15933 11883 15991 11889
rect 15933 11880 15945 11883
rect 15252 11852 15945 11880
rect 15252 11840 15258 11852
rect 15933 11849 15945 11852
rect 15979 11849 15991 11883
rect 16758 11880 16764 11892
rect 16719 11852 16764 11880
rect 15933 11843 15991 11849
rect 16758 11840 16764 11852
rect 16816 11880 16822 11892
rect 17402 11880 17408 11892
rect 16816 11852 17408 11880
rect 16816 11840 16822 11852
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 12207 11784 12664 11812
rect 12207 11781 12219 11784
rect 12161 11775 12219 11781
rect 13538 11772 13544 11824
rect 13596 11812 13602 11824
rect 17681 11815 17739 11821
rect 17681 11812 17693 11815
rect 13596 11784 17693 11812
rect 13596 11772 13602 11784
rect 17681 11781 17693 11784
rect 17727 11781 17739 11815
rect 17681 11775 17739 11781
rect 5307 11716 6868 11744
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11676 3663 11679
rect 4522 11676 4528 11688
rect 3651 11648 4528 11676
rect 3651 11645 3663 11648
rect 3605 11639 3663 11645
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 5920 11685 5948 11716
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7009 11747 7067 11753
rect 7009 11744 7021 11747
rect 6972 11716 7021 11744
rect 6972 11704 6978 11716
rect 7009 11713 7021 11716
rect 7055 11713 7067 11747
rect 7009 11707 7067 11713
rect 8570 11704 8576 11756
rect 8628 11744 8634 11756
rect 9125 11747 9183 11753
rect 9125 11744 9137 11747
rect 8628 11716 9137 11744
rect 8628 11704 8634 11716
rect 9125 11713 9137 11716
rect 9171 11713 9183 11747
rect 9125 11707 9183 11713
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 10410 11744 10416 11756
rect 9999 11716 10416 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 12713 11747 12771 11753
rect 12713 11713 12725 11747
rect 12759 11744 12771 11747
rect 12802 11744 12808 11756
rect 12759 11716 12808 11744
rect 12759 11713 12771 11716
rect 12713 11707 12771 11713
rect 12802 11704 12808 11716
rect 12860 11744 12866 11756
rect 13173 11747 13231 11753
rect 13173 11744 13185 11747
rect 12860 11716 13185 11744
rect 12860 11704 12866 11716
rect 13173 11713 13185 11716
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 15013 11747 15071 11753
rect 15013 11744 15025 11747
rect 14240 11716 15025 11744
rect 14240 11704 14246 11716
rect 15013 11713 15025 11716
rect 15059 11713 15071 11747
rect 15013 11707 15071 11713
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 6089 11679 6147 11685
rect 6089 11645 6101 11679
rect 6135 11645 6147 11679
rect 6089 11639 6147 11645
rect 1857 11611 1915 11617
rect 1857 11577 1869 11611
rect 1903 11608 1915 11611
rect 2774 11608 2780 11620
rect 1903 11580 2780 11608
rect 1903 11577 1915 11580
rect 1857 11571 1915 11577
rect 2774 11568 2780 11580
rect 2832 11568 2838 11620
rect 2866 11568 2872 11620
rect 2924 11568 2930 11620
rect 6104 11608 6132 11639
rect 6270 11636 6276 11688
rect 6328 11676 6334 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 6328 11648 7205 11676
rect 6328 11636 6334 11648
rect 7193 11645 7205 11648
rect 7239 11645 7251 11679
rect 7193 11639 7251 11645
rect 7282 11636 7288 11688
rect 7340 11676 7346 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 7340 11648 7757 11676
rect 7340 11636 7346 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11645 8171 11679
rect 8113 11639 8171 11645
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11676 8263 11679
rect 8251 11648 8524 11676
rect 8251 11645 8263 11648
rect 8205 11639 8263 11645
rect 7374 11608 7380 11620
rect 6104 11580 7380 11608
rect 7374 11568 7380 11580
rect 7432 11568 7438 11620
rect 8128 11608 8156 11639
rect 8386 11608 8392 11620
rect 8128 11580 8392 11608
rect 8386 11568 8392 11580
rect 8444 11568 8450 11620
rect 8496 11608 8524 11648
rect 8662 11636 8668 11688
rect 8720 11676 8726 11688
rect 9217 11679 9275 11685
rect 9217 11676 9229 11679
rect 8720 11648 9229 11676
rect 8720 11636 8726 11648
rect 9217 11645 9229 11648
rect 9263 11645 9275 11679
rect 9398 11676 9404 11688
rect 9359 11648 9404 11676
rect 9217 11639 9275 11645
rect 8757 11611 8815 11617
rect 8757 11608 8769 11611
rect 8496 11580 8769 11608
rect 8757 11577 8769 11580
rect 8803 11577 8815 11611
rect 9232 11608 9260 11639
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 10042 11676 10048 11688
rect 10003 11648 10048 11676
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 10226 11676 10232 11688
rect 10187 11648 10232 11676
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 12529 11679 12587 11685
rect 12529 11645 12541 11679
rect 12575 11676 12587 11679
rect 12618 11676 12624 11688
rect 12575 11648 12624 11676
rect 12575 11645 12587 11648
rect 12529 11639 12587 11645
rect 12618 11636 12624 11648
rect 12676 11676 12682 11688
rect 14642 11676 14648 11688
rect 12676 11648 14648 11676
rect 12676 11636 12682 11648
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11645 14979 11679
rect 15028 11676 15056 11707
rect 15102 11704 15108 11756
rect 15160 11744 15166 11756
rect 15746 11744 15752 11756
rect 15160 11716 15205 11744
rect 15304 11716 15752 11744
rect 15160 11704 15166 11716
rect 15304 11676 15332 11716
rect 15746 11704 15752 11716
rect 15804 11744 15810 11756
rect 16393 11747 16451 11753
rect 16393 11744 16405 11747
rect 15804 11716 16405 11744
rect 15804 11704 15810 11716
rect 16393 11713 16405 11716
rect 16439 11713 16451 11747
rect 17696 11744 17724 11775
rect 17865 11747 17923 11753
rect 17865 11744 17877 11747
rect 17696 11716 17877 11744
rect 16393 11707 16451 11713
rect 17865 11713 17877 11716
rect 17911 11713 17923 11747
rect 17865 11707 17923 11713
rect 16022 11676 16028 11688
rect 15028 11648 15332 11676
rect 15983 11648 16028 11676
rect 14921 11639 14979 11645
rect 9766 11608 9772 11620
rect 9232 11580 9772 11608
rect 8757 11571 8815 11577
rect 9766 11568 9772 11580
rect 9824 11568 9830 11620
rect 10502 11568 10508 11620
rect 10560 11608 10566 11620
rect 14090 11608 14096 11620
rect 10560 11580 14096 11608
rect 10560 11568 10566 11580
rect 14090 11568 14096 11580
rect 14148 11568 14154 11620
rect 14826 11568 14832 11620
rect 14884 11608 14890 11620
rect 14936 11608 14964 11639
rect 16022 11636 16028 11648
rect 16080 11636 16086 11688
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11645 16175 11679
rect 16117 11639 16175 11645
rect 16132 11608 16160 11639
rect 14884 11580 16160 11608
rect 14884 11568 14890 11580
rect 2225 11543 2283 11549
rect 2225 11509 2237 11543
rect 2271 11540 2283 11543
rect 2884 11540 2912 11568
rect 2271 11512 2912 11540
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 3050 11500 3056 11552
rect 3108 11540 3114 11552
rect 3973 11543 4031 11549
rect 3973 11540 3985 11543
rect 3108 11512 3985 11540
rect 3108 11500 3114 11512
rect 3973 11509 3985 11512
rect 4019 11509 4031 11543
rect 3973 11503 4031 11509
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 6270 11540 6276 11552
rect 5960 11512 6276 11540
rect 5960 11500 5966 11512
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 6454 11540 6460 11552
rect 6415 11512 6460 11540
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 7558 11540 7564 11552
rect 6972 11512 7564 11540
rect 6972 11500 6978 11512
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 8665 11543 8723 11549
rect 8665 11509 8677 11543
rect 8711 11540 8723 11543
rect 9306 11540 9312 11552
rect 8711 11512 9312 11540
rect 8711 11509 8723 11512
rect 8665 11503 8723 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 9548 11512 9597 11540
rect 9548 11500 9554 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 11790 11540 11796 11552
rect 9732 11512 11796 11540
rect 9732 11500 9738 11512
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 14553 11543 14611 11549
rect 14553 11540 14565 11543
rect 13872 11512 14565 11540
rect 13872 11500 13878 11512
rect 14553 11509 14565 11512
rect 14599 11540 14611 11543
rect 15102 11540 15108 11552
rect 14599 11512 15108 11540
rect 14599 11509 14611 11512
rect 14553 11503 14611 11509
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15473 11543 15531 11549
rect 15473 11540 15485 11543
rect 15436 11512 15485 11540
rect 15436 11500 15442 11512
rect 15473 11509 15485 11512
rect 15519 11509 15531 11543
rect 15473 11503 15531 11509
rect 15562 11500 15568 11552
rect 15620 11540 15626 11552
rect 15620 11512 15665 11540
rect 15620 11500 15626 11512
rect 16022 11500 16028 11552
rect 16080 11540 16086 11552
rect 16206 11540 16212 11552
rect 16080 11512 16212 11540
rect 16080 11500 16086 11512
rect 16206 11500 16212 11512
rect 16264 11540 16270 11552
rect 16945 11543 17003 11549
rect 16945 11540 16957 11543
rect 16264 11512 16957 11540
rect 16264 11500 16270 11512
rect 16945 11509 16957 11512
rect 16991 11509 17003 11543
rect 16945 11503 17003 11509
rect 18049 11543 18107 11549
rect 18049 11509 18061 11543
rect 18095 11540 18107 11543
rect 18230 11540 18236 11552
rect 18095 11512 18236 11540
rect 18095 11509 18107 11512
rect 18049 11503 18107 11509
rect 18230 11500 18236 11512
rect 18288 11500 18294 11552
rect 1104 11450 18860 11472
rect 1104 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 3302 11450
rect 3354 11398 3366 11450
rect 3418 11398 3430 11450
rect 3482 11398 7622 11450
rect 7674 11398 7686 11450
rect 7738 11398 7750 11450
rect 7802 11398 7814 11450
rect 7866 11398 7878 11450
rect 7930 11398 12070 11450
rect 12122 11398 12134 11450
rect 12186 11398 12198 11450
rect 12250 11398 12262 11450
rect 12314 11398 12326 11450
rect 12378 11398 16518 11450
rect 16570 11398 16582 11450
rect 16634 11398 16646 11450
rect 16698 11398 16710 11450
rect 16762 11398 16774 11450
rect 16826 11398 18860 11450
rect 1104 11376 18860 11398
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 6362 11336 6368 11348
rect 2556 11308 6368 11336
rect 2556 11296 2562 11308
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 6880 11308 7757 11336
rect 6880 11296 6886 11308
rect 7745 11305 7757 11308
rect 7791 11305 7803 11339
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 7745 11299 7803 11305
rect 7852 11308 8953 11336
rect 4525 11271 4583 11277
rect 4525 11237 4537 11271
rect 4571 11237 4583 11271
rect 4525 11231 4583 11237
rect 3050 11200 3056 11212
rect 3011 11172 3056 11200
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 3237 11203 3295 11209
rect 3237 11169 3249 11203
rect 3283 11200 3295 11203
rect 4540 11200 4568 11231
rect 7006 11228 7012 11280
rect 7064 11268 7070 11280
rect 7852 11268 7880 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 9398 11296 9404 11348
rect 9456 11336 9462 11348
rect 9582 11336 9588 11348
rect 9456 11308 9588 11336
rect 9456 11296 9462 11308
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 9766 11336 9772 11348
rect 9727 11308 9772 11336
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 15746 11336 15752 11348
rect 14200 11308 15752 11336
rect 9490 11268 9496 11280
rect 7064 11240 7880 11268
rect 8220 11240 9496 11268
rect 7064 11228 7070 11240
rect 4706 11200 4712 11212
rect 3283 11172 4712 11200
rect 3283 11169 3295 11172
rect 3237 11163 3295 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 6362 11160 6368 11212
rect 6420 11200 6426 11212
rect 7282 11200 7288 11212
rect 6420 11172 7288 11200
rect 6420 11160 6426 11172
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 8220 11209 8248 11240
rect 9490 11228 9496 11240
rect 9548 11228 9554 11280
rect 12710 11228 12716 11280
rect 12768 11268 12774 11280
rect 13078 11268 13084 11280
rect 12768 11240 13084 11268
rect 12768 11228 12774 11240
rect 13078 11228 13084 11240
rect 13136 11268 13142 11280
rect 14200 11268 14228 11308
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 15838 11296 15844 11348
rect 15896 11336 15902 11348
rect 15896 11308 17632 11336
rect 15896 11296 15902 11308
rect 16117 11271 16175 11277
rect 16117 11268 16129 11271
rect 13136 11240 14228 11268
rect 14568 11240 16129 11268
rect 13136 11228 13142 11240
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 8294 11160 8300 11212
rect 8352 11200 8358 11212
rect 8570 11200 8576 11212
rect 8352 11172 8397 11200
rect 8531 11172 8576 11200
rect 8352 11160 8358 11172
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 9582 11160 9588 11212
rect 9640 11200 9646 11212
rect 14568 11209 14596 11240
rect 16117 11237 16129 11240
rect 16163 11237 16175 11271
rect 16117 11231 16175 11237
rect 16945 11271 17003 11277
rect 16945 11237 16957 11271
rect 16991 11237 17003 11271
rect 16945 11231 17003 11237
rect 14553 11203 14611 11209
rect 9640 11172 9685 11200
rect 9640 11160 9646 11172
rect 14553 11169 14565 11203
rect 14599 11169 14611 11203
rect 14734 11200 14740 11212
rect 14695 11172 14740 11200
rect 14553 11163 14611 11169
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 15378 11200 15384 11212
rect 15339 11172 15384 11200
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 15473 11203 15531 11209
rect 15473 11169 15485 11203
rect 15519 11200 15531 11203
rect 15519 11172 15700 11200
rect 15519 11169 15531 11172
rect 15473 11163 15531 11169
rect 2958 11132 2964 11144
rect 2919 11104 2964 11132
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 4522 11092 4528 11144
rect 4580 11132 4586 11144
rect 5638 11135 5696 11141
rect 5638 11132 5650 11135
rect 4580 11104 5650 11132
rect 4580 11092 4586 11104
rect 5638 11101 5650 11104
rect 5684 11101 5696 11135
rect 5638 11095 5696 11101
rect 5810 11092 5816 11144
rect 5868 11132 5874 11144
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 5868 11104 5917 11132
rect 5868 11092 5874 11104
rect 5905 11101 5917 11104
rect 5951 11101 5963 11135
rect 5905 11095 5963 11101
rect 6178 11092 6184 11144
rect 6236 11132 6242 11144
rect 7653 11135 7711 11141
rect 7653 11132 7665 11135
rect 6236 11104 7665 11132
rect 6236 11092 6242 11104
rect 7653 11101 7665 11104
rect 7699 11132 7711 11135
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 7699 11104 8125 11132
rect 7699 11101 7711 11104
rect 7653 11095 7711 11101
rect 8113 11101 8125 11104
rect 8159 11132 8171 11135
rect 9306 11132 9312 11144
rect 8159 11104 8800 11132
rect 9267 11104 9312 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 6270 11024 6276 11076
rect 6328 11064 6334 11076
rect 8662 11064 8668 11076
rect 6328 11036 8668 11064
rect 6328 11024 6334 11036
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 8772 11064 8800 11104
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11132 9459 11135
rect 9447 11104 11284 11132
rect 9447 11101 9459 11104
rect 9401 11095 9459 11101
rect 9582 11064 9588 11076
rect 8772 11036 9588 11064
rect 9582 11024 9588 11036
rect 9640 11024 9646 11076
rect 9953 11067 10011 11073
rect 9953 11033 9965 11067
rect 9999 11064 10011 11067
rect 10042 11064 10048 11076
rect 9999 11036 10048 11064
rect 9999 11033 10011 11036
rect 9953 11027 10011 11033
rect 2590 10996 2596 11008
rect 2551 10968 2596 10996
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 4062 10956 4068 11008
rect 4120 10996 4126 11008
rect 9968 10996 9996 11027
rect 10042 11024 10048 11036
rect 10100 11064 10106 11076
rect 10962 11064 10968 11076
rect 10100 11036 10968 11064
rect 10100 11024 10106 11036
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 4120 10968 9996 10996
rect 11256 10996 11284 11104
rect 11514 11092 11520 11144
rect 11572 11132 11578 11144
rect 11701 11135 11759 11141
rect 11701 11132 11713 11135
rect 11572 11104 11713 11132
rect 11572 11092 11578 11104
rect 11701 11101 11713 11104
rect 11747 11101 11759 11135
rect 15289 11135 15347 11141
rect 11701 11095 11759 11101
rect 14384 11104 15240 11132
rect 11330 11024 11336 11076
rect 11388 11064 11394 11076
rect 11946 11067 12004 11073
rect 11946 11064 11958 11067
rect 11388 11036 11958 11064
rect 11388 11024 11394 11036
rect 11946 11033 11958 11036
rect 11992 11064 12004 11067
rect 14384 11064 14412 11104
rect 11992 11036 14412 11064
rect 14461 11067 14519 11073
rect 11992 11033 12004 11036
rect 11946 11027 12004 11033
rect 14461 11033 14473 11067
rect 14507 11064 14519 11067
rect 14642 11064 14648 11076
rect 14507 11036 14648 11064
rect 14507 11033 14519 11036
rect 14461 11027 14519 11033
rect 14642 11024 14648 11036
rect 14700 11024 14706 11076
rect 15212 11064 15240 11104
rect 15289 11101 15301 11135
rect 15335 11132 15347 11135
rect 15562 11132 15568 11144
rect 15335 11104 15568 11132
rect 15335 11101 15347 11104
rect 15289 11095 15347 11101
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 15672 11132 15700 11172
rect 15746 11160 15752 11212
rect 15804 11200 15810 11212
rect 16669 11203 16727 11209
rect 16669 11200 16681 11203
rect 15804 11172 16681 11200
rect 15804 11160 15810 11172
rect 16669 11169 16681 11172
rect 16715 11169 16727 11203
rect 16669 11163 16727 11169
rect 15838 11132 15844 11144
rect 15672 11104 15844 11132
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11132 16543 11135
rect 16960 11132 16988 11231
rect 17402 11200 17408 11212
rect 17363 11172 17408 11200
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 17497 11203 17555 11209
rect 17497 11169 17509 11203
rect 17543 11169 17555 11203
rect 17497 11163 17555 11169
rect 16531 11104 16988 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 17218 11064 17224 11076
rect 15212 11036 17224 11064
rect 17218 11024 17224 11036
rect 17276 11064 17282 11076
rect 17512 11064 17540 11163
rect 17276 11036 17540 11064
rect 17604 11064 17632 11308
rect 18049 11271 18107 11277
rect 18049 11237 18061 11271
rect 18095 11268 18107 11271
rect 18138 11268 18144 11280
rect 18095 11240 18144 11268
rect 18095 11237 18107 11240
rect 18049 11231 18107 11237
rect 18138 11228 18144 11240
rect 18196 11228 18202 11280
rect 17862 11132 17868 11144
rect 17823 11104 17868 11132
rect 17862 11092 17868 11104
rect 17920 11132 17926 11144
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 17920 11104 18245 11132
rect 17920 11092 17926 11104
rect 18233 11101 18245 11104
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 18506 11064 18512 11076
rect 17604 11036 18512 11064
rect 17276 11024 17282 11036
rect 14093 10999 14151 11005
rect 14093 10996 14105 10999
rect 11256 10968 14105 10996
rect 4120 10956 4126 10968
rect 14093 10965 14105 10968
rect 14139 10965 14151 10999
rect 14918 10996 14924 11008
rect 14879 10968 14924 10996
rect 14093 10959 14151 10965
rect 14918 10956 14924 10968
rect 14976 10956 14982 11008
rect 16577 10999 16635 11005
rect 16577 10965 16589 10999
rect 16623 10996 16635 10999
rect 16850 10996 16856 11008
rect 16623 10968 16856 10996
rect 16623 10965 16635 10968
rect 16577 10959 16635 10965
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 17313 10999 17371 11005
rect 17313 10965 17325 10999
rect 17359 10996 17371 10999
rect 17604 10996 17632 11036
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 17359 10968 17632 10996
rect 17359 10965 17371 10968
rect 17313 10959 17371 10965
rect 1104 10906 18860 10928
rect 1104 10854 5398 10906
rect 5450 10854 5462 10906
rect 5514 10854 5526 10906
rect 5578 10854 5590 10906
rect 5642 10854 5654 10906
rect 5706 10854 9846 10906
rect 9898 10854 9910 10906
rect 9962 10854 9974 10906
rect 10026 10854 10038 10906
rect 10090 10854 10102 10906
rect 10154 10854 14294 10906
rect 14346 10854 14358 10906
rect 14410 10854 14422 10906
rect 14474 10854 14486 10906
rect 14538 10854 14550 10906
rect 14602 10854 18860 10906
rect 1104 10832 18860 10854
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 2682 10792 2688 10804
rect 2363 10764 2688 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 2682 10752 2688 10764
rect 2740 10792 2746 10804
rect 2777 10795 2835 10801
rect 2777 10792 2789 10795
rect 2740 10764 2789 10792
rect 2740 10752 2746 10764
rect 2777 10761 2789 10764
rect 2823 10761 2835 10795
rect 2777 10755 2835 10761
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 6914 10792 6920 10804
rect 4120 10764 6920 10792
rect 4120 10752 4126 10764
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 8205 10795 8263 10801
rect 7116 10764 7328 10792
rect 1946 10684 1952 10736
rect 2004 10724 2010 10736
rect 2133 10727 2191 10733
rect 2133 10724 2145 10727
rect 2004 10696 2145 10724
rect 2004 10684 2010 10696
rect 2133 10693 2145 10696
rect 2179 10724 2191 10727
rect 3697 10727 3755 10733
rect 3697 10724 3709 10727
rect 2179 10696 3709 10724
rect 2179 10693 2191 10696
rect 2133 10687 2191 10693
rect 3697 10693 3709 10696
rect 3743 10724 3755 10727
rect 4154 10724 4160 10736
rect 3743 10696 4160 10724
rect 3743 10693 3755 10696
rect 3697 10687 3755 10693
rect 4154 10684 4160 10696
rect 4212 10684 4218 10736
rect 5902 10684 5908 10736
rect 5960 10733 5966 10736
rect 5960 10724 5972 10733
rect 6822 10724 6828 10736
rect 5960 10696 6828 10724
rect 5960 10687 5972 10696
rect 5960 10684 5966 10687
rect 6822 10684 6828 10696
rect 6880 10684 6886 10736
rect 3050 10616 3056 10668
rect 3108 10656 3114 10668
rect 7116 10665 7144 10764
rect 7300 10724 7328 10764
rect 8205 10761 8217 10795
rect 8251 10792 8263 10795
rect 9398 10792 9404 10804
rect 8251 10764 9404 10792
rect 8251 10761 8263 10764
rect 8205 10755 8263 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 11517 10795 11575 10801
rect 11517 10761 11529 10795
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 8386 10724 8392 10736
rect 7300 10696 8392 10724
rect 8386 10684 8392 10696
rect 8444 10684 8450 10736
rect 11532 10724 11560 10755
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 14369 10795 14427 10801
rect 14369 10792 14381 10795
rect 11756 10764 14381 10792
rect 11756 10752 11762 10764
rect 14369 10761 14381 10764
rect 14415 10761 14427 10795
rect 14642 10792 14648 10804
rect 14603 10764 14648 10792
rect 14369 10755 14427 10761
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 15105 10795 15163 10801
rect 15105 10761 15117 10795
rect 15151 10792 15163 10795
rect 16669 10795 16727 10801
rect 16669 10792 16681 10795
rect 15151 10764 16681 10792
rect 15151 10761 15163 10764
rect 15105 10755 15163 10761
rect 16669 10761 16681 10764
rect 16715 10761 16727 10795
rect 16669 10755 16727 10761
rect 13256 10727 13314 10733
rect 13256 10724 13268 10727
rect 11532 10696 13268 10724
rect 13256 10693 13268 10696
rect 13302 10724 13314 10727
rect 13354 10724 13360 10736
rect 13302 10696 13360 10724
rect 13302 10693 13314 10696
rect 13256 10687 13314 10693
rect 13354 10684 13360 10696
rect 13412 10684 13418 10736
rect 16482 10684 16488 10736
rect 16540 10724 16546 10736
rect 17037 10727 17095 10733
rect 17037 10724 17049 10727
rect 16540 10696 17049 10724
rect 16540 10684 16546 10696
rect 17037 10693 17049 10696
rect 17083 10724 17095 10727
rect 17494 10724 17500 10736
rect 17083 10696 17500 10724
rect 17083 10693 17095 10696
rect 17037 10687 17095 10693
rect 17494 10684 17500 10696
rect 17552 10684 17558 10736
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 3108 10628 3617 10656
rect 3108 10616 3114 10628
rect 3605 10625 3617 10628
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 7092 10659 7150 10665
rect 7092 10625 7104 10659
rect 7138 10625 7150 10659
rect 7092 10619 7150 10625
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 9410 10659 9468 10665
rect 9410 10656 9422 10659
rect 8260 10628 9422 10656
rect 8260 10616 8266 10628
rect 9410 10625 9422 10628
rect 9456 10625 9468 10659
rect 9410 10619 9468 10625
rect 10128 10659 10186 10665
rect 10128 10625 10140 10659
rect 10174 10656 10186 10659
rect 11698 10656 11704 10668
rect 10174 10628 11704 10656
rect 10174 10625 10186 10628
rect 10128 10619 10186 10625
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 12618 10616 12624 10668
rect 12676 10665 12682 10668
rect 12676 10656 12688 10665
rect 15013 10659 15071 10665
rect 12676 10628 12721 10656
rect 12676 10619 12688 10628
rect 15013 10625 15025 10659
rect 15059 10656 15071 10659
rect 16942 10656 16948 10668
rect 15059 10628 16948 10656
rect 15059 10625 15071 10628
rect 15013 10619 15071 10625
rect 12676 10616 12682 10619
rect 2222 10548 2228 10600
rect 2280 10588 2286 10600
rect 2866 10588 2872 10600
rect 2280 10560 2872 10588
rect 2280 10548 2286 10560
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10588 3019 10591
rect 3881 10591 3939 10597
rect 3881 10588 3893 10591
rect 3007 10560 3893 10588
rect 3007 10557 3019 10560
rect 2961 10551 3019 10557
rect 3881 10557 3893 10560
rect 3927 10588 3939 10591
rect 4982 10588 4988 10600
rect 3927 10560 4988 10588
rect 3927 10557 3939 10560
rect 3881 10551 3939 10557
rect 4982 10548 4988 10560
rect 5040 10548 5046 10600
rect 6181 10591 6239 10597
rect 6181 10557 6193 10591
rect 6227 10588 6239 10591
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6227 10560 6837 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 9674 10588 9680 10600
rect 9635 10560 9680 10588
rect 6825 10551 6883 10557
rect 2409 10455 2467 10461
rect 2409 10421 2421 10455
rect 2455 10452 2467 10455
rect 2498 10452 2504 10464
rect 2455 10424 2504 10452
rect 2455 10421 2467 10424
rect 2409 10415 2467 10421
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 2682 10412 2688 10464
rect 2740 10452 2746 10464
rect 3237 10455 3295 10461
rect 3237 10452 3249 10455
rect 2740 10424 3249 10452
rect 2740 10412 2746 10424
rect 3237 10421 3249 10424
rect 3283 10421 3295 10455
rect 4154 10452 4160 10464
rect 4115 10424 4160 10452
rect 3237 10415 3295 10421
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 4890 10452 4896 10464
rect 4847 10424 4896 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 4890 10412 4896 10424
rect 4948 10452 4954 10464
rect 5258 10452 5264 10464
rect 4948 10424 5264 10452
rect 4948 10412 4954 10424
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5810 10412 5816 10464
rect 5868 10452 5874 10464
rect 6196 10452 6224 10551
rect 9674 10548 9680 10560
rect 9732 10588 9738 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9732 10560 9873 10588
rect 9732 10548 9738 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 12894 10588 12900 10600
rect 12855 10560 12900 10588
rect 9861 10551 9919 10557
rect 12894 10548 12900 10560
rect 12952 10588 12958 10600
rect 12989 10591 13047 10597
rect 12989 10588 13001 10591
rect 12952 10560 13001 10588
rect 12952 10548 12958 10560
rect 12989 10557 13001 10560
rect 13035 10557 13047 10591
rect 14458 10588 14464 10600
rect 14419 10560 14464 10588
rect 12989 10551 13047 10557
rect 14458 10548 14464 10560
rect 14516 10588 14522 10600
rect 15028 10588 15056 10619
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17696 10628 17877 10656
rect 14516 10560 15056 10588
rect 15289 10591 15347 10597
rect 14516 10548 14522 10560
rect 15289 10557 15301 10591
rect 15335 10588 15347 10591
rect 15746 10588 15752 10600
rect 15335 10560 15752 10588
rect 15335 10557 15347 10560
rect 15289 10551 15347 10557
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 17129 10591 17187 10597
rect 17129 10557 17141 10591
rect 17175 10557 17187 10591
rect 17129 10551 17187 10557
rect 8297 10523 8355 10529
rect 8297 10489 8309 10523
rect 8343 10489 8355 10523
rect 8297 10483 8355 10489
rect 5868 10424 6224 10452
rect 5868 10412 5874 10424
rect 6822 10412 6828 10464
rect 6880 10452 6886 10464
rect 8312 10452 8340 10483
rect 10962 10480 10968 10532
rect 11020 10520 11026 10532
rect 16393 10523 16451 10529
rect 16393 10520 16405 10523
rect 11020 10492 11744 10520
rect 11020 10480 11026 10492
rect 6880 10424 8340 10452
rect 11241 10455 11299 10461
rect 6880 10412 6886 10424
rect 11241 10421 11253 10455
rect 11287 10452 11299 10455
rect 11606 10452 11612 10464
rect 11287 10424 11612 10452
rect 11287 10421 11299 10424
rect 11241 10415 11299 10421
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 11716 10452 11744 10492
rect 14384 10492 16405 10520
rect 14384 10452 14412 10492
rect 16393 10489 16405 10492
rect 16439 10520 16451 10523
rect 17144 10520 17172 10551
rect 17218 10548 17224 10600
rect 17276 10588 17282 10600
rect 17276 10560 17321 10588
rect 17276 10548 17282 10560
rect 17696 10529 17724 10628
rect 17865 10625 17877 10628
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 17681 10523 17739 10529
rect 17681 10520 17693 10523
rect 16439 10492 17693 10520
rect 16439 10489 16451 10492
rect 16393 10483 16451 10489
rect 17681 10489 17693 10492
rect 17727 10489 17739 10523
rect 17681 10483 17739 10489
rect 11716 10424 14412 10452
rect 15746 10412 15752 10464
rect 15804 10452 15810 10464
rect 15930 10452 15936 10464
rect 15804 10424 15936 10452
rect 15804 10412 15810 10424
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 18049 10455 18107 10461
rect 18049 10421 18061 10455
rect 18095 10452 18107 10455
rect 18322 10452 18328 10464
rect 18095 10424 18328 10452
rect 18095 10421 18107 10424
rect 18049 10415 18107 10421
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 1104 10362 18860 10384
rect 1104 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 3430 10362
rect 3482 10310 7622 10362
rect 7674 10310 7686 10362
rect 7738 10310 7750 10362
rect 7802 10310 7814 10362
rect 7866 10310 7878 10362
rect 7930 10310 12070 10362
rect 12122 10310 12134 10362
rect 12186 10310 12198 10362
rect 12250 10310 12262 10362
rect 12314 10310 12326 10362
rect 12378 10310 16518 10362
rect 16570 10310 16582 10362
rect 16634 10310 16646 10362
rect 16698 10310 16710 10362
rect 16762 10310 16774 10362
rect 16826 10310 18860 10362
rect 1104 10288 18860 10310
rect 6546 10248 6552 10260
rect 6507 10220 6552 10248
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 9033 10251 9091 10257
rect 9033 10248 9045 10251
rect 8260 10220 9045 10248
rect 8260 10208 8266 10220
rect 9033 10217 9045 10220
rect 9079 10217 9091 10251
rect 11425 10251 11483 10257
rect 11425 10248 11437 10251
rect 9033 10211 9091 10217
rect 9140 10220 11437 10248
rect 2406 10140 2412 10192
rect 2464 10180 2470 10192
rect 2464 10152 2636 10180
rect 2464 10140 2470 10152
rect 2498 10112 2504 10124
rect 2459 10084 2504 10112
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 2608 10121 2636 10152
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 9140 10180 9168 10220
rect 11425 10217 11437 10220
rect 11471 10248 11483 10251
rect 14734 10248 14740 10260
rect 11471 10220 14740 10248
rect 11471 10217 11483 10220
rect 11425 10211 11483 10217
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 15654 10208 15660 10260
rect 15712 10248 15718 10260
rect 16393 10251 16451 10257
rect 16393 10248 16405 10251
rect 15712 10220 16405 10248
rect 15712 10208 15718 10220
rect 16393 10217 16405 10220
rect 16439 10217 16451 10251
rect 16393 10211 16451 10217
rect 16577 10251 16635 10257
rect 16577 10217 16589 10251
rect 16623 10248 16635 10251
rect 16850 10248 16856 10260
rect 16623 10220 16856 10248
rect 16623 10217 16635 10220
rect 16577 10211 16635 10217
rect 8444 10152 9168 10180
rect 8444 10140 8450 10152
rect 2593 10115 2651 10121
rect 2593 10081 2605 10115
rect 2639 10081 2651 10115
rect 3050 10112 3056 10124
rect 3011 10084 3056 10112
rect 2593 10075 2651 10081
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 16408 10112 16436 10211
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 17402 10208 17408 10260
rect 17460 10248 17466 10260
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 17460 10220 17693 10248
rect 17460 10208 17466 10220
rect 17681 10217 17693 10220
rect 17727 10217 17739 10251
rect 17681 10211 17739 10217
rect 17034 10112 17040 10124
rect 16408 10084 17040 10112
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 17218 10112 17224 10124
rect 17179 10084 17224 10112
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 1946 10044 1952 10056
rect 1907 10016 1952 10044
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 2682 10044 2688 10056
rect 2455 10016 2688 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 2682 10004 2688 10016
rect 2740 10004 2746 10056
rect 4430 10004 4436 10056
rect 4488 10044 4494 10056
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4488 10016 4537 10044
rect 4488 10004 4494 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 4792 10047 4850 10053
rect 4792 10013 4804 10047
rect 4838 10013 4850 10047
rect 4792 10007 4850 10013
rect 4706 9936 4712 9988
rect 4764 9976 4770 9988
rect 4816 9976 4844 10007
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 7929 10047 7987 10053
rect 7929 10044 7941 10047
rect 6880 10016 7941 10044
rect 6880 10004 6886 10016
rect 7929 10013 7941 10016
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 10134 10004 10140 10056
rect 10192 10053 10198 10056
rect 10192 10044 10204 10053
rect 10410 10044 10416 10056
rect 10192 10016 10237 10044
rect 10371 10016 10416 10044
rect 10192 10007 10204 10016
rect 10192 10004 10198 10007
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 11514 10004 11520 10056
rect 11572 10044 11578 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 11572 10016 12817 10044
rect 11572 10004 11578 10016
rect 12805 10013 12817 10016
rect 12851 10044 12863 10047
rect 12894 10044 12900 10056
rect 12851 10016 12900 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 17696 10044 17724 10211
rect 17865 10047 17923 10053
rect 17865 10044 17877 10047
rect 17696 10016 17877 10044
rect 17865 10013 17877 10016
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 4764 9948 4844 9976
rect 5276 9948 6684 9976
rect 4764 9936 4770 9948
rect 1394 9868 1400 9920
rect 1452 9908 1458 9920
rect 1765 9911 1823 9917
rect 1765 9908 1777 9911
rect 1452 9880 1777 9908
rect 1452 9868 1458 9880
rect 1765 9877 1777 9880
rect 1811 9877 1823 9911
rect 1765 9871 1823 9877
rect 1854 9868 1860 9920
rect 1912 9908 1918 9920
rect 2041 9911 2099 9917
rect 2041 9908 2053 9911
rect 1912 9880 2053 9908
rect 1912 9868 1918 9880
rect 2041 9877 2053 9880
rect 2087 9877 2099 9911
rect 2041 9871 2099 9877
rect 2866 9868 2872 9920
rect 2924 9908 2930 9920
rect 3329 9911 3387 9917
rect 3329 9908 3341 9911
rect 2924 9880 3341 9908
rect 2924 9868 2930 9880
rect 3329 9877 3341 9880
rect 3375 9908 3387 9911
rect 5276 9908 5304 9948
rect 5902 9908 5908 9920
rect 3375 9880 5304 9908
rect 5863 9880 5908 9908
rect 3375 9877 3387 9880
rect 3329 9871 3387 9877
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 6656 9908 6684 9948
rect 7374 9936 7380 9988
rect 7432 9976 7438 9988
rect 7662 9979 7720 9985
rect 7662 9976 7674 9979
rect 7432 9948 7674 9976
rect 7432 9936 7438 9948
rect 7662 9945 7674 9948
rect 7708 9945 7720 9979
rect 12560 9979 12618 9985
rect 7662 9939 7720 9945
rect 10336 9948 12434 9976
rect 10336 9908 10364 9948
rect 6656 9880 10364 9908
rect 12406 9908 12434 9948
rect 12560 9945 12572 9979
rect 12606 9976 12618 9979
rect 13078 9976 13084 9988
rect 12606 9948 13084 9976
rect 12606 9945 12618 9948
rect 12560 9939 12618 9945
rect 13078 9936 13084 9948
rect 13136 9936 13142 9988
rect 14182 9908 14188 9920
rect 12406 9880 14188 9908
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 16390 9868 16396 9920
rect 16448 9908 16454 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 16448 9880 16957 9908
rect 16448 9868 16454 9880
rect 16945 9877 16957 9880
rect 16991 9908 17003 9911
rect 17494 9908 17500 9920
rect 16991 9880 17500 9908
rect 16991 9877 17003 9880
rect 16945 9871 17003 9877
rect 17494 9868 17500 9880
rect 17552 9868 17558 9920
rect 18049 9911 18107 9917
rect 18049 9877 18061 9911
rect 18095 9908 18107 9911
rect 18506 9908 18512 9920
rect 18095 9880 18512 9908
rect 18095 9877 18107 9880
rect 18049 9871 18107 9877
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 1104 9818 18860 9840
rect 1104 9766 5398 9818
rect 5450 9766 5462 9818
rect 5514 9766 5526 9818
rect 5578 9766 5590 9818
rect 5642 9766 5654 9818
rect 5706 9766 9846 9818
rect 9898 9766 9910 9818
rect 9962 9766 9974 9818
rect 10026 9766 10038 9818
rect 10090 9766 10102 9818
rect 10154 9766 14294 9818
rect 14346 9766 14358 9818
rect 14410 9766 14422 9818
rect 14474 9766 14486 9818
rect 14538 9766 14550 9818
rect 14602 9766 18860 9818
rect 1104 9744 18860 9766
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 16022 9704 16028 9716
rect 4212 9676 16028 9704
rect 4212 9664 4218 9676
rect 16022 9664 16028 9676
rect 16080 9664 16086 9716
rect 2682 9596 2688 9648
rect 2740 9636 2746 9648
rect 5568 9639 5626 9645
rect 2740 9608 2820 9636
rect 2740 9596 2746 9608
rect 1946 9528 1952 9580
rect 2004 9568 2010 9580
rect 2041 9571 2099 9577
rect 2041 9568 2053 9571
rect 2004 9540 2053 9568
rect 2004 9528 2010 9540
rect 2041 9537 2053 9540
rect 2087 9568 2099 9571
rect 2222 9568 2228 9580
rect 2087 9540 2228 9568
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2498 9528 2504 9580
rect 2556 9568 2562 9580
rect 2593 9571 2651 9577
rect 2593 9568 2605 9571
rect 2556 9540 2605 9568
rect 2556 9528 2562 9540
rect 2593 9537 2605 9540
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 2314 9460 2320 9512
rect 2372 9500 2378 9512
rect 2792 9509 2820 9608
rect 5568 9605 5580 9639
rect 5614 9636 5626 9639
rect 6546 9636 6552 9648
rect 5614 9608 6552 9636
rect 5614 9605 5626 9608
rect 5568 9599 5626 9605
rect 6546 9596 6552 9608
rect 6604 9596 6610 9648
rect 9582 9636 9588 9648
rect 8588 9608 9588 9636
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 7098 9568 7104 9580
rect 4120 9540 7104 9568
rect 4120 9528 4126 9540
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7282 9568 7288 9580
rect 7243 9540 7288 9568
rect 7282 9528 7288 9540
rect 7340 9568 7346 9580
rect 8018 9568 8024 9580
rect 7340 9540 8024 9568
rect 7340 9528 7346 9540
rect 8018 9528 8024 9540
rect 8076 9568 8082 9580
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 8076 9540 8401 9568
rect 8076 9528 8082 9540
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2372 9472 2697 9500
rect 2372 9460 2378 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 5810 9500 5816 9512
rect 2823 9472 4844 9500
rect 5771 9472 5816 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 1857 9435 1915 9441
rect 1857 9401 1869 9435
rect 1903 9432 1915 9435
rect 2866 9432 2872 9444
rect 1903 9404 2872 9432
rect 1903 9401 1915 9404
rect 1857 9395 1915 9401
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 4433 9435 4491 9441
rect 4433 9401 4445 9435
rect 4479 9432 4491 9435
rect 4522 9432 4528 9444
rect 4479 9404 4528 9432
rect 4479 9401 4491 9404
rect 4433 9395 4491 9401
rect 4522 9392 4528 9404
rect 4580 9392 4586 9444
rect 2222 9364 2228 9376
rect 2183 9336 2228 9364
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 4816 9364 4844 9472
rect 5810 9460 5816 9472
rect 5868 9500 5874 9512
rect 6822 9500 6828 9512
rect 5868 9472 6828 9500
rect 5868 9460 5874 9472
rect 6822 9460 6828 9472
rect 6880 9500 6886 9512
rect 8588 9509 8616 9608
rect 9582 9596 9588 9608
rect 9640 9636 9646 9648
rect 10410 9636 10416 9648
rect 9640 9608 10416 9636
rect 9640 9596 9646 9608
rect 10410 9596 10416 9608
rect 10468 9636 10474 9648
rect 11514 9636 11520 9648
rect 10468 9608 11520 9636
rect 10468 9596 10474 9608
rect 11514 9596 11520 9608
rect 11572 9596 11578 9648
rect 13020 9639 13078 9645
rect 13020 9605 13032 9639
rect 13066 9636 13078 9639
rect 14826 9636 14832 9648
rect 13066 9608 14832 9636
rect 13066 9605 13078 9608
rect 13020 9599 13078 9605
rect 14826 9596 14832 9608
rect 14884 9596 14890 9648
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 8829 9571 8887 9577
rect 8829 9568 8841 9571
rect 8720 9540 8841 9568
rect 8720 9528 8726 9540
rect 8829 9537 8841 9540
rect 8875 9537 8887 9571
rect 16114 9568 16120 9580
rect 8829 9531 8887 9537
rect 9600 9540 16120 9568
rect 7653 9503 7711 9509
rect 7653 9500 7665 9503
rect 6880 9472 7665 9500
rect 6880 9460 6886 9472
rect 7653 9469 7665 9472
rect 7699 9500 7711 9503
rect 8573 9503 8631 9509
rect 8573 9500 8585 9503
rect 7699 9472 8585 9500
rect 7699 9469 7711 9472
rect 7653 9463 7711 9469
rect 8573 9469 8585 9472
rect 8619 9469 8631 9503
rect 8573 9463 8631 9469
rect 6086 9364 6092 9376
rect 4816 9336 6092 9364
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 9600 9364 9628 9540
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 17678 9568 17684 9580
rect 17639 9540 17684 9568
rect 17678 9528 17684 9540
rect 17736 9568 17742 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17736 9540 17877 9568
rect 17736 9528 17742 9540
rect 17865 9537 17877 9540
rect 17911 9537 17923 9571
rect 17865 9531 17923 9537
rect 18233 9571 18291 9577
rect 18233 9537 18245 9571
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 13262 9500 13268 9512
rect 13223 9472 13268 9500
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 17954 9500 17960 9512
rect 13872 9472 17960 9500
rect 13872 9460 13878 9472
rect 17954 9460 17960 9472
rect 18012 9500 18018 9512
rect 18248 9500 18276 9531
rect 18012 9472 18276 9500
rect 18012 9460 18018 9472
rect 9674 9392 9680 9444
rect 9732 9432 9738 9444
rect 9732 9404 12020 9432
rect 9732 9392 9738 9404
rect 6236 9336 9628 9364
rect 6236 9324 6242 9336
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 9824 9336 9965 9364
rect 9824 9324 9830 9336
rect 9953 9333 9965 9336
rect 9999 9333 10011 9367
rect 11882 9364 11888 9376
rect 11843 9336 11888 9364
rect 9953 9327 10011 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 11992 9364 12020 9404
rect 14642 9364 14648 9376
rect 11992 9336 14648 9364
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 15381 9367 15439 9373
rect 15381 9333 15393 9367
rect 15427 9364 15439 9367
rect 16850 9364 16856 9376
rect 15427 9336 16856 9364
rect 15427 9333 15439 9336
rect 15381 9327 15439 9333
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 18046 9364 18052 9376
rect 18007 9336 18052 9364
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 18414 9364 18420 9376
rect 18375 9336 18420 9364
rect 18414 9324 18420 9336
rect 18472 9324 18478 9376
rect 1104 9274 18860 9296
rect 1104 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 3430 9274
rect 3482 9222 7622 9274
rect 7674 9222 7686 9274
rect 7738 9222 7750 9274
rect 7802 9222 7814 9274
rect 7866 9222 7878 9274
rect 7930 9222 12070 9274
rect 12122 9222 12134 9274
rect 12186 9222 12198 9274
rect 12250 9222 12262 9274
rect 12314 9222 12326 9274
rect 12378 9222 16518 9274
rect 16570 9222 16582 9274
rect 16634 9222 16646 9274
rect 16698 9222 16710 9274
rect 16762 9222 16774 9274
rect 16826 9222 18860 9274
rect 1104 9200 18860 9222
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 2133 9163 2191 9169
rect 2133 9160 2145 9163
rect 2004 9132 2145 9160
rect 2004 9120 2010 9132
rect 2133 9129 2145 9132
rect 2179 9129 2191 9163
rect 2498 9160 2504 9172
rect 2459 9132 2504 9160
rect 2133 9123 2191 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 6178 9160 6184 9172
rect 4304 9132 6184 9160
rect 4304 9120 4310 9132
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 7374 9160 7380 9172
rect 6871 9132 7380 9160
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 9674 9160 9680 9172
rect 7616 9132 9680 9160
rect 7616 9120 7622 9132
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10137 9163 10195 9169
rect 10137 9129 10149 9163
rect 10183 9160 10195 9163
rect 10226 9160 10232 9172
rect 10183 9132 10232 9160
rect 10183 9129 10195 9132
rect 10137 9123 10195 9129
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 11330 9160 11336 9172
rect 10612 9132 11336 9160
rect 2409 9095 2467 9101
rect 2409 9061 2421 9095
rect 2455 9092 2467 9095
rect 3142 9092 3148 9104
rect 2455 9064 3148 9092
rect 2455 9061 2467 9064
rect 2409 9055 2467 9061
rect 3142 9052 3148 9064
rect 3200 9092 3206 9104
rect 3970 9092 3976 9104
rect 3200 9064 3976 9092
rect 3200 9052 3206 9064
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 8757 9095 8815 9101
rect 8757 9061 8769 9095
rect 8803 9092 8815 9095
rect 10612 9092 10640 9132
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 11977 9163 12035 9169
rect 11977 9129 11989 9163
rect 12023 9160 12035 9163
rect 12618 9160 12624 9172
rect 12023 9132 12624 9160
rect 12023 9129 12035 9132
rect 11977 9123 12035 9129
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 14734 9120 14740 9172
rect 14792 9160 14798 9172
rect 15289 9163 15347 9169
rect 15289 9160 15301 9163
rect 14792 9132 15301 9160
rect 14792 9120 14798 9132
rect 15289 9129 15301 9132
rect 15335 9160 15347 9163
rect 16206 9160 16212 9172
rect 15335 9132 16212 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 16390 9160 16396 9172
rect 16351 9132 16396 9160
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 18012 9132 18061 9160
rect 18012 9120 18018 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 18049 9123 18107 9129
rect 8803 9064 10640 9092
rect 8803 9061 8815 9064
rect 8757 9055 8815 9061
rect 16114 9052 16120 9104
rect 16172 9092 16178 9104
rect 17126 9092 17132 9104
rect 16172 9064 17132 9092
rect 16172 9052 16178 9064
rect 17126 9052 17132 9064
rect 17184 9052 17190 9104
rect 2498 8984 2504 9036
rect 2556 9024 2562 9036
rect 3053 9027 3111 9033
rect 3053 9024 3065 9027
rect 2556 8996 3065 9024
rect 2556 8984 2562 8996
rect 3053 8993 3065 8996
rect 3099 8993 3111 9027
rect 11514 9024 11520 9036
rect 3053 8987 3111 8993
rect 6472 8996 7512 9024
rect 11475 8996 11520 9024
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 3970 8956 3976 8968
rect 3660 8928 3976 8956
rect 3660 8916 3666 8928
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 4448 8928 5365 8956
rect 4448 8900 4476 8928
rect 5353 8925 5365 8928
rect 5399 8956 5411 8959
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 5399 8928 5457 8956
rect 5399 8925 5411 8928
rect 5353 8919 5411 8925
rect 5445 8925 5457 8928
rect 5491 8956 5503 8959
rect 5491 8928 5856 8956
rect 5491 8925 5503 8928
rect 5445 8919 5503 8925
rect 5828 8900 5856 8928
rect 2869 8891 2927 8897
rect 2869 8857 2881 8891
rect 2915 8888 2927 8891
rect 3329 8891 3387 8897
rect 3329 8888 3341 8891
rect 2915 8860 3341 8888
rect 2915 8857 2927 8860
rect 2869 8851 2927 8857
rect 3329 8857 3341 8860
rect 3375 8857 3387 8891
rect 3329 8851 3387 8857
rect 4430 8848 4436 8900
rect 4488 8848 4494 8900
rect 4982 8848 4988 8900
rect 5040 8888 5046 8900
rect 5718 8897 5724 8900
rect 5086 8891 5144 8897
rect 5086 8888 5098 8891
rect 5040 8860 5098 8888
rect 5040 8848 5046 8860
rect 5086 8857 5098 8860
rect 5132 8857 5144 8891
rect 5712 8888 5724 8897
rect 5679 8860 5724 8888
rect 5086 8851 5144 8857
rect 5712 8851 5724 8860
rect 5718 8848 5724 8851
rect 5776 8848 5782 8900
rect 5810 8848 5816 8900
rect 5868 8848 5874 8900
rect 6472 8888 6500 8996
rect 6822 8916 6828 8968
rect 6880 8956 6886 8968
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 6880 8928 7389 8956
rect 6880 8916 6886 8928
rect 7377 8925 7389 8928
rect 7423 8925 7435 8959
rect 7484 8956 7512 8996
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 14553 9027 14611 9033
rect 14553 8993 14565 9027
rect 14599 9024 14611 9027
rect 16022 9024 16028 9036
rect 14599 8996 16028 9024
rect 14599 8993 14611 8996
rect 14553 8987 14611 8993
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 7484 8928 7788 8956
rect 7377 8919 7435 8925
rect 5920 8860 6500 8888
rect 2958 8820 2964 8832
rect 2871 8792 2964 8820
rect 2958 8780 2964 8792
rect 3016 8820 3022 8832
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3016 8792 3801 8820
rect 3016 8780 3022 8792
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 3973 8823 4031 8829
rect 3973 8789 3985 8823
rect 4019 8820 4031 8823
rect 4154 8820 4160 8832
rect 4019 8792 4160 8820
rect 4019 8789 4031 8792
rect 3973 8783 4031 8789
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 5920 8820 5948 8860
rect 7098 8848 7104 8900
rect 7156 8888 7162 8900
rect 7622 8891 7680 8897
rect 7622 8888 7634 8891
rect 7156 8860 7634 8888
rect 7156 8848 7162 8860
rect 7622 8857 7634 8860
rect 7668 8857 7680 8891
rect 7760 8888 7788 8928
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 11250 8959 11308 8965
rect 11250 8956 11262 8959
rect 9824 8928 11262 8956
rect 9824 8916 9830 8928
rect 11250 8925 11262 8928
rect 11296 8925 11308 8959
rect 11532 8956 11560 8984
rect 13262 8956 13268 8968
rect 11532 8928 13268 8956
rect 11250 8919 11308 8925
rect 13262 8916 13268 8928
rect 13320 8956 13326 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 13320 8928 13369 8956
rect 13320 8916 13326 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 14734 8956 14740 8968
rect 14695 8928 14740 8956
rect 13357 8919 13415 8925
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8956 15991 8959
rect 16850 8956 16856 8968
rect 15979 8928 16856 8956
rect 15979 8925 15991 8928
rect 15933 8919 15991 8925
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 17328 8928 17509 8956
rect 13112 8891 13170 8897
rect 7760 8860 12434 8888
rect 7622 8851 7680 8857
rect 5224 8792 5948 8820
rect 5224 8780 5230 8792
rect 6086 8780 6092 8832
rect 6144 8820 6150 8832
rect 8662 8820 8668 8832
rect 6144 8792 8668 8820
rect 6144 8780 6150 8792
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 12406 8820 12434 8860
rect 13112 8857 13124 8891
rect 13158 8888 13170 8891
rect 13446 8888 13452 8900
rect 13158 8860 13452 8888
rect 13158 8857 13170 8860
rect 13112 8851 13170 8857
rect 13446 8848 13452 8860
rect 13504 8848 13510 8900
rect 17328 8897 17356 8928
rect 17497 8925 17509 8928
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 17313 8891 17371 8897
rect 17313 8888 17325 8891
rect 14108 8860 17325 8888
rect 14108 8820 14136 8860
rect 17313 8857 17325 8860
rect 17359 8857 17371 8891
rect 17313 8851 17371 8857
rect 12406 8792 14136 8820
rect 14277 8823 14335 8829
rect 14277 8789 14289 8823
rect 14323 8820 14335 8823
rect 14642 8820 14648 8832
rect 14323 8792 14648 8820
rect 14323 8789 14335 8792
rect 14277 8783 14335 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 15102 8820 15108 8832
rect 15063 8792 15108 8820
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 15470 8820 15476 8832
rect 15431 8792 15476 8820
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 15841 8823 15899 8829
rect 15841 8789 15853 8823
rect 15887 8820 15899 8823
rect 16114 8820 16120 8832
rect 15887 8792 16120 8820
rect 15887 8789 15899 8792
rect 15841 8783 15899 8789
rect 16114 8780 16120 8792
rect 16172 8820 16178 8832
rect 16390 8820 16396 8832
rect 16172 8792 16396 8820
rect 16172 8780 16178 8792
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 17681 8823 17739 8829
rect 17681 8789 17693 8823
rect 17727 8820 17739 8823
rect 17770 8820 17776 8832
rect 17727 8792 17776 8820
rect 17727 8789 17739 8792
rect 17681 8783 17739 8789
rect 17770 8780 17776 8792
rect 17828 8780 17834 8832
rect 1104 8730 18860 8752
rect 1104 8678 5398 8730
rect 5450 8678 5462 8730
rect 5514 8678 5526 8730
rect 5578 8678 5590 8730
rect 5642 8678 5654 8730
rect 5706 8678 9846 8730
rect 9898 8678 9910 8730
rect 9962 8678 9974 8730
rect 10026 8678 10038 8730
rect 10090 8678 10102 8730
rect 10154 8678 14294 8730
rect 14346 8678 14358 8730
rect 14410 8678 14422 8730
rect 14474 8678 14486 8730
rect 14538 8678 14550 8730
rect 14602 8678 18860 8730
rect 1104 8656 18860 8678
rect 1857 8619 1915 8625
rect 1857 8585 1869 8619
rect 1903 8616 1915 8619
rect 2222 8616 2228 8628
rect 1903 8588 2228 8616
rect 1903 8585 1915 8588
rect 1857 8579 1915 8585
rect 2222 8576 2228 8588
rect 2280 8576 2286 8628
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 9766 8616 9772 8628
rect 2372 8588 2417 8616
rect 2608 8588 9772 8616
rect 2372 8576 2378 8588
rect 1946 8412 1952 8424
rect 1907 8384 1952 8412
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2133 8415 2191 8421
rect 2133 8381 2145 8415
rect 2179 8412 2191 8415
rect 2608 8412 2636 8588
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 12897 8619 12955 8625
rect 12897 8585 12909 8619
rect 12943 8585 12955 8619
rect 12897 8579 12955 8585
rect 14369 8619 14427 8625
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 14826 8616 14832 8628
rect 14415 8588 14832 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 2777 8551 2835 8557
rect 2777 8517 2789 8551
rect 2823 8548 2835 8551
rect 4065 8551 4123 8557
rect 4065 8548 4077 8551
rect 2823 8520 4077 8548
rect 2823 8517 2835 8520
rect 2777 8511 2835 8517
rect 4065 8517 4077 8520
rect 4111 8548 4123 8551
rect 4246 8548 4252 8560
rect 4111 8520 4252 8548
rect 4111 8517 4123 8520
rect 4065 8511 4123 8517
rect 4246 8508 4252 8520
rect 4304 8508 4310 8560
rect 4890 8508 4896 8560
rect 4948 8548 4954 8560
rect 4948 8520 5948 8548
rect 4948 8508 4954 8520
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8480 2743 8483
rect 3142 8480 3148 8492
rect 2731 8452 3148 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 2792 8424 2820 8452
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3510 8480 3516 8492
rect 3471 8452 3516 8480
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 4976 8483 5034 8489
rect 4976 8480 4988 8483
rect 3804 8452 4988 8480
rect 2179 8384 2636 8412
rect 2179 8381 2191 8384
rect 2133 8375 2191 8381
rect 2774 8372 2780 8424
rect 2832 8372 2838 8424
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8381 3019 8415
rect 3602 8412 3608 8424
rect 3563 8384 3608 8412
rect 2961 8375 3019 8381
rect 1489 8347 1547 8353
rect 1489 8313 1501 8347
rect 1535 8344 1547 8347
rect 1762 8344 1768 8356
rect 1535 8316 1768 8344
rect 1535 8313 1547 8316
rect 1489 8307 1547 8313
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 2222 8304 2228 8356
rect 2280 8344 2286 8356
rect 2498 8344 2504 8356
rect 2280 8316 2504 8344
rect 2280 8304 2286 8316
rect 2498 8304 2504 8316
rect 2556 8344 2562 8356
rect 2976 8344 3004 8375
rect 3602 8372 3608 8384
rect 3660 8372 3666 8424
rect 3804 8421 3832 8452
rect 4976 8449 4988 8452
rect 5022 8480 5034 8483
rect 5810 8480 5816 8492
rect 5022 8452 5816 8480
rect 5022 8449 5034 8452
rect 4976 8443 5034 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 5920 8480 5948 8520
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 9300 8551 9358 8557
rect 6880 8520 7788 8548
rect 6880 8508 6886 8520
rect 7760 8489 7788 8520
rect 9300 8517 9312 8551
rect 9346 8548 9358 8551
rect 9398 8548 9404 8560
rect 9346 8520 9404 8548
rect 9346 8517 9358 8520
rect 9300 8511 9358 8517
rect 9398 8508 9404 8520
rect 9456 8508 9462 8560
rect 12912 8548 12940 8579
rect 14826 8576 14832 8588
rect 14884 8576 14890 8628
rect 15749 8619 15807 8625
rect 15749 8585 15761 8619
rect 15795 8616 15807 8619
rect 16298 8616 16304 8628
rect 15795 8588 16304 8616
rect 15795 8585 15807 8588
rect 15749 8579 15807 8585
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 17034 8576 17040 8628
rect 17092 8616 17098 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17092 8588 17509 8616
rect 17092 8576 17098 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 13256 8551 13314 8557
rect 13256 8548 13268 8551
rect 11532 8520 12434 8548
rect 12912 8520 13268 8548
rect 11532 8492 11560 8520
rect 7478 8483 7536 8489
rect 7478 8480 7490 8483
rect 5920 8452 7490 8480
rect 7478 8449 7490 8452
rect 7524 8449 7536 8483
rect 7478 8443 7536 8449
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8480 7803 8483
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 7791 8452 9045 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 9033 8449 9045 8452
rect 9079 8449 9091 8483
rect 11514 8480 11520 8492
rect 11475 8452 11520 8480
rect 9033 8443 9091 8449
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 11773 8483 11831 8489
rect 11773 8480 11785 8483
rect 11664 8452 11785 8480
rect 11664 8440 11670 8452
rect 11773 8449 11785 8452
rect 11819 8449 11831 8483
rect 12406 8480 12434 8520
rect 13256 8517 13268 8520
rect 13302 8548 13314 8551
rect 16022 8548 16028 8560
rect 13302 8520 16028 8548
rect 13302 8517 13314 8520
rect 13256 8511 13314 8517
rect 16022 8508 16028 8520
rect 16080 8508 16086 8560
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12406 8452 13001 8480
rect 11773 8443 11831 8449
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 17512 8480 17540 8579
rect 17681 8483 17739 8489
rect 17681 8480 17693 8483
rect 17512 8452 17693 8480
rect 12989 8443 13047 8449
rect 17681 8449 17693 8452
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 3804 8344 3832 8375
rect 4430 8372 4436 8424
rect 4488 8412 4494 8424
rect 4709 8415 4767 8421
rect 4709 8412 4721 8415
rect 4488 8384 4721 8412
rect 4488 8372 4494 8384
rect 4709 8381 4721 8384
rect 4755 8381 4767 8415
rect 4709 8375 4767 8381
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 14734 8412 14740 8424
rect 14608 8384 14740 8412
rect 14608 8372 14614 8384
rect 14734 8372 14740 8384
rect 14792 8372 14798 8424
rect 15841 8415 15899 8421
rect 15841 8381 15853 8415
rect 15887 8381 15899 8415
rect 16022 8412 16028 8424
rect 15983 8384 16028 8412
rect 15841 8375 15899 8381
rect 6086 8344 6092 8356
rect 2556 8316 3832 8344
rect 6047 8316 6092 8344
rect 2556 8304 2562 8316
rect 6086 8304 6092 8316
rect 6144 8304 6150 8356
rect 15194 8344 15200 8356
rect 10244 8316 10548 8344
rect 15155 8316 15200 8344
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3145 8279 3203 8285
rect 3145 8276 3157 8279
rect 3016 8248 3157 8276
rect 3016 8236 3022 8248
rect 3145 8245 3157 8248
rect 3191 8245 3203 8279
rect 3145 8239 3203 8245
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 6365 8279 6423 8285
rect 6365 8276 6377 8279
rect 5776 8248 6377 8276
rect 5776 8236 5782 8248
rect 6365 8245 6377 8248
rect 6411 8245 6423 8279
rect 6365 8239 6423 8245
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 10244 8276 10272 8316
rect 10410 8276 10416 8288
rect 8628 8248 10272 8276
rect 10371 8248 10416 8276
rect 8628 8236 8634 8248
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 10520 8276 10548 8316
rect 15194 8304 15200 8316
rect 15252 8344 15258 8356
rect 15856 8344 15884 8375
rect 16022 8372 16028 8384
rect 16080 8372 16086 8424
rect 15252 8316 15884 8344
rect 15252 8304 15258 8316
rect 17678 8304 17684 8356
rect 17736 8344 17742 8356
rect 17865 8347 17923 8353
rect 17865 8344 17877 8347
rect 17736 8316 17877 8344
rect 17736 8304 17742 8316
rect 17865 8313 17877 8316
rect 17911 8313 17923 8347
rect 17865 8307 17923 8313
rect 14734 8276 14740 8288
rect 10520 8248 14740 8276
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 15378 8276 15384 8288
rect 15339 8248 15384 8276
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 1104 8186 18860 8208
rect 1104 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 3430 8186
rect 3482 8134 7622 8186
rect 7674 8134 7686 8186
rect 7738 8134 7750 8186
rect 7802 8134 7814 8186
rect 7866 8134 7878 8186
rect 7930 8134 12070 8186
rect 12122 8134 12134 8186
rect 12186 8134 12198 8186
rect 12250 8134 12262 8186
rect 12314 8134 12326 8186
rect 12378 8134 16518 8186
rect 16570 8134 16582 8186
rect 16634 8134 16646 8186
rect 16698 8134 16710 8186
rect 16762 8134 16774 8186
rect 16826 8134 18860 8186
rect 1104 8112 18860 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 1765 8075 1823 8081
rect 1765 8072 1777 8075
rect 1636 8044 1777 8072
rect 1636 8032 1642 8044
rect 1765 8041 1777 8044
rect 1811 8041 1823 8075
rect 1765 8035 1823 8041
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 2004 8044 2145 8072
rect 2004 8032 2010 8044
rect 2133 8041 2145 8044
rect 2179 8041 2191 8075
rect 2133 8035 2191 8041
rect 14734 8032 14740 8084
rect 14792 8072 14798 8084
rect 18046 8072 18052 8084
rect 14792 8044 18052 8072
rect 14792 8032 14798 8044
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 1670 7964 1676 8016
rect 1728 8004 1734 8016
rect 2041 8007 2099 8013
rect 2041 8004 2053 8007
rect 1728 7976 2053 8004
rect 1728 7964 1734 7976
rect 2041 7973 2053 7976
rect 2087 7973 2099 8007
rect 4522 8004 4528 8016
rect 2041 7967 2099 7973
rect 2516 7976 4528 8004
rect 1486 7896 1492 7948
rect 1544 7936 1550 7948
rect 2516 7936 2544 7976
rect 4522 7964 4528 7976
rect 4580 7964 4586 8016
rect 16942 8004 16948 8016
rect 16903 7976 16948 8004
rect 16942 7964 16948 7976
rect 17000 7964 17006 8016
rect 2682 7936 2688 7948
rect 1544 7908 2544 7936
rect 2643 7908 2688 7936
rect 1544 7896 1550 7908
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 14826 7896 14832 7948
rect 14884 7936 14890 7948
rect 14921 7939 14979 7945
rect 14921 7936 14933 7939
rect 14884 7908 14933 7936
rect 14884 7896 14890 7908
rect 14921 7905 14933 7908
rect 14967 7905 14979 7939
rect 14921 7899 14979 7905
rect 15105 7939 15163 7945
rect 15105 7905 15117 7939
rect 15151 7936 15163 7939
rect 15378 7936 15384 7948
rect 15151 7908 15384 7936
rect 15151 7905 15163 7908
rect 15105 7899 15163 7905
rect 15378 7896 15384 7908
rect 15436 7896 15442 7948
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2958 7868 2964 7880
rect 2639 7840 2964 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 4488 7840 4537 7868
rect 4488 7828 4494 7840
rect 4525 7837 4537 7840
rect 4571 7868 4583 7871
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 4571 7840 6929 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 6917 7837 6929 7840
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8352 7840 8953 7868
rect 8352 7828 8358 7840
rect 8941 7837 8953 7840
rect 8987 7868 8999 7871
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 8987 7840 10517 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 10505 7837 10517 7840
rect 10551 7868 10563 7871
rect 10594 7868 10600 7880
rect 10551 7840 10600 7868
rect 10551 7837 10563 7840
rect 10505 7831 10563 7837
rect 10594 7828 10600 7840
rect 10652 7868 10658 7880
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 10652 7840 12081 7868
rect 10652 7828 10658 7840
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 15197 7871 15255 7877
rect 12069 7831 12127 7837
rect 12176 7840 15148 7868
rect 2406 7760 2412 7812
rect 2464 7800 2470 7812
rect 2682 7800 2688 7812
rect 2464 7772 2688 7800
rect 2464 7760 2470 7772
rect 2682 7760 2688 7772
rect 2740 7800 2746 7812
rect 4154 7800 4160 7812
rect 2740 7772 4160 7800
rect 2740 7760 2746 7772
rect 4154 7760 4160 7772
rect 4212 7800 4218 7812
rect 4770 7803 4828 7809
rect 4770 7800 4782 7803
rect 4212 7772 4782 7800
rect 4212 7760 4218 7772
rect 4770 7769 4782 7772
rect 4816 7769 4828 7803
rect 4770 7763 4828 7769
rect 7184 7803 7242 7809
rect 7184 7769 7196 7803
rect 7230 7800 7242 7803
rect 7466 7800 7472 7812
rect 7230 7772 7472 7800
rect 7230 7769 7242 7772
rect 7184 7763 7242 7769
rect 7466 7760 7472 7772
rect 7524 7760 7530 7812
rect 9186 7803 9244 7809
rect 9186 7800 9198 7803
rect 8496 7772 9198 7800
rect 8496 7744 8524 7772
rect 9186 7769 9198 7772
rect 9232 7769 9244 7803
rect 9186 7763 9244 7769
rect 10410 7760 10416 7812
rect 10468 7800 10474 7812
rect 10750 7803 10808 7809
rect 10750 7800 10762 7803
rect 10468 7772 10762 7800
rect 10468 7760 10474 7772
rect 10750 7769 10762 7772
rect 10796 7800 10808 7803
rect 12176 7800 12204 7840
rect 10796 7772 12204 7800
rect 12336 7803 12394 7809
rect 10796 7769 10808 7772
rect 10750 7763 10808 7769
rect 12336 7769 12348 7803
rect 12382 7800 12394 7803
rect 13262 7800 13268 7812
rect 12382 7772 13268 7800
rect 12382 7769 12394 7772
rect 12336 7763 12394 7769
rect 13262 7760 13268 7772
rect 13320 7760 13326 7812
rect 15120 7800 15148 7840
rect 15197 7837 15209 7871
rect 15243 7868 15255 7871
rect 15470 7868 15476 7880
rect 15243 7840 15476 7868
rect 15243 7837 15255 7840
rect 15197 7831 15255 7837
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 16960 7868 16988 7964
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 16960 7840 17049 7868
rect 17037 7837 17049 7840
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 16114 7800 16120 7812
rect 15120 7772 16120 7800
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 2130 7692 2136 7744
rect 2188 7732 2194 7744
rect 2501 7735 2559 7741
rect 2501 7732 2513 7735
rect 2188 7704 2513 7732
rect 2188 7692 2194 7704
rect 2501 7701 2513 7704
rect 2547 7701 2559 7735
rect 2501 7695 2559 7701
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 3145 7735 3203 7741
rect 3145 7732 3157 7735
rect 2832 7704 3157 7732
rect 2832 7692 2838 7704
rect 3145 7701 3157 7704
rect 3191 7732 3203 7735
rect 3878 7732 3884 7744
rect 3191 7704 3884 7732
rect 3191 7701 3203 7704
rect 3145 7695 3203 7701
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 5626 7692 5632 7744
rect 5684 7732 5690 7744
rect 5905 7735 5963 7741
rect 5905 7732 5917 7735
rect 5684 7704 5917 7732
rect 5684 7692 5690 7704
rect 5905 7701 5917 7704
rect 5951 7732 5963 7735
rect 6086 7732 6092 7744
rect 5951 7704 6092 7732
rect 5951 7701 5963 7704
rect 5905 7695 5963 7701
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 8297 7735 8355 7741
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 8478 7732 8484 7744
rect 8343 7704 8484 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 9306 7692 9312 7744
rect 9364 7732 9370 7744
rect 10321 7735 10379 7741
rect 10321 7732 10333 7735
rect 9364 7704 10333 7732
rect 9364 7692 9370 7704
rect 10321 7701 10333 7704
rect 10367 7701 10379 7735
rect 10321 7695 10379 7701
rect 11885 7735 11943 7741
rect 11885 7701 11897 7735
rect 11931 7732 11943 7735
rect 12250 7732 12256 7744
rect 11931 7704 12256 7732
rect 11931 7701 11943 7704
rect 11885 7695 11943 7701
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 13446 7732 13452 7744
rect 13407 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 14734 7732 14740 7744
rect 14608 7704 14740 7732
rect 14608 7692 14614 7704
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 15378 7692 15384 7744
rect 15436 7732 15442 7744
rect 15565 7735 15623 7741
rect 15565 7732 15577 7735
rect 15436 7704 15577 7732
rect 15436 7692 15442 7704
rect 15565 7701 15577 7704
rect 15611 7701 15623 7735
rect 17218 7732 17224 7744
rect 17179 7704 17224 7732
rect 15565 7695 15623 7701
rect 17218 7692 17224 7704
rect 17276 7692 17282 7744
rect 1104 7642 18860 7664
rect 1104 7590 5398 7642
rect 5450 7590 5462 7642
rect 5514 7590 5526 7642
rect 5578 7590 5590 7642
rect 5642 7590 5654 7642
rect 5706 7590 9846 7642
rect 9898 7590 9910 7642
rect 9962 7590 9974 7642
rect 10026 7590 10038 7642
rect 10090 7590 10102 7642
rect 10154 7590 14294 7642
rect 14346 7590 14358 7642
rect 14410 7590 14422 7642
rect 14474 7590 14486 7642
rect 14538 7590 14550 7642
rect 14602 7590 18860 7642
rect 1104 7568 18860 7590
rect 1486 7488 1492 7540
rect 1544 7528 1550 7540
rect 1765 7531 1823 7537
rect 1765 7528 1777 7531
rect 1544 7500 1777 7528
rect 1544 7488 1550 7500
rect 1765 7497 1777 7500
rect 1811 7497 1823 7531
rect 2130 7528 2136 7540
rect 2091 7500 2136 7528
rect 1765 7491 1823 7497
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 2593 7531 2651 7537
rect 2593 7497 2605 7531
rect 2639 7528 2651 7531
rect 2774 7528 2780 7540
rect 2639 7500 2780 7528
rect 2639 7497 2651 7500
rect 2593 7491 2651 7497
rect 2774 7488 2780 7500
rect 2832 7488 2838 7540
rect 2961 7531 3019 7537
rect 2961 7497 2973 7531
rect 3007 7528 3019 7531
rect 3602 7528 3608 7540
rect 3007 7500 3608 7528
rect 3007 7497 3019 7500
rect 2961 7491 3019 7497
rect 3602 7488 3608 7500
rect 3660 7488 3666 7540
rect 3786 7488 3792 7540
rect 3844 7528 3850 7540
rect 3970 7528 3976 7540
rect 3844 7500 3976 7528
rect 3844 7488 3850 7500
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 14182 7528 14188 7540
rect 4580 7500 14188 7528
rect 4580 7488 4586 7500
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 14553 7531 14611 7537
rect 14553 7497 14565 7531
rect 14599 7528 14611 7531
rect 14921 7531 14979 7537
rect 14921 7528 14933 7531
rect 14599 7500 14933 7528
rect 14599 7497 14611 7500
rect 14553 7491 14611 7497
rect 14921 7497 14933 7500
rect 14967 7497 14979 7531
rect 15378 7528 15384 7540
rect 15339 7500 15384 7528
rect 14921 7491 14979 7497
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 17126 7528 17132 7540
rect 17039 7500 17132 7528
rect 17126 7488 17132 7500
rect 17184 7528 17190 7540
rect 17497 7531 17555 7537
rect 17497 7528 17509 7531
rect 17184 7500 17509 7528
rect 17184 7488 17190 7500
rect 17497 7497 17509 7500
rect 17543 7497 17555 7531
rect 17497 7491 17555 7497
rect 1670 7420 1676 7472
rect 1728 7460 1734 7472
rect 2501 7463 2559 7469
rect 2501 7460 2513 7463
rect 1728 7432 2513 7460
rect 1728 7420 1734 7432
rect 2222 7392 2228 7404
rect 1504 7364 2228 7392
rect 1504 7333 1532 7364
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 1489 7327 1547 7333
rect 1489 7293 1501 7327
rect 1535 7293 1547 7327
rect 1670 7324 1676 7336
rect 1631 7296 1676 7324
rect 1489 7287 1547 7293
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 2332 7188 2360 7432
rect 2501 7429 2513 7432
rect 2547 7429 2559 7463
rect 2501 7423 2559 7429
rect 4430 7420 4436 7472
rect 4488 7460 4494 7472
rect 4488 7432 5948 7460
rect 4488 7420 4494 7432
rect 3602 7392 3608 7404
rect 3344 7364 3608 7392
rect 2409 7327 2467 7333
rect 2409 7293 2421 7327
rect 2455 7293 2467 7327
rect 2409 7287 2467 7293
rect 2424 7256 2452 7287
rect 2424 7228 3096 7256
rect 2774 7188 2780 7200
rect 2332 7160 2780 7188
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 3068 7197 3096 7228
rect 3053 7191 3111 7197
rect 3053 7157 3065 7191
rect 3099 7188 3111 7191
rect 3344 7188 3372 7364
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 4177 7395 4235 7401
rect 4177 7361 4189 7395
rect 4223 7392 4235 7395
rect 5166 7392 5172 7404
rect 4223 7364 5172 7392
rect 4223 7361 4235 7364
rect 4177 7355 4235 7361
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 5626 7352 5632 7404
rect 5684 7401 5690 7404
rect 5920 7401 5948 7432
rect 6454 7420 6460 7472
rect 6512 7460 6518 7472
rect 6730 7460 6736 7472
rect 6512 7432 6736 7460
rect 6512 7420 6518 7432
rect 6730 7420 6736 7432
rect 6788 7420 6794 7472
rect 11882 7420 11888 7472
rect 11940 7460 11946 7472
rect 12314 7463 12372 7469
rect 12314 7460 12326 7463
rect 11940 7432 12326 7460
rect 11940 7420 11946 7432
rect 12314 7429 12326 7432
rect 12360 7460 12372 7463
rect 12360 7432 15608 7460
rect 12360 7429 12372 7432
rect 12314 7423 12372 7429
rect 5684 7392 5696 7401
rect 5905 7395 5963 7401
rect 5684 7364 5729 7392
rect 5684 7355 5696 7364
rect 5905 7361 5917 7395
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 7857 7395 7915 7401
rect 7857 7361 7869 7395
rect 7903 7392 7915 7395
rect 8018 7392 8024 7404
rect 7903 7364 8024 7392
rect 7903 7361 7915 7364
rect 7857 7355 7915 7361
rect 5684 7352 5690 7355
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 10330 7395 10388 7401
rect 10330 7392 10342 7395
rect 9364 7364 10342 7392
rect 9364 7352 9370 7364
rect 10330 7361 10342 7364
rect 10376 7361 10388 7395
rect 10594 7392 10600 7404
rect 10555 7364 10600 7392
rect 10330 7355 10388 7361
rect 10594 7352 10600 7364
rect 10652 7392 10658 7404
rect 11974 7392 11980 7404
rect 10652 7364 11980 7392
rect 10652 7352 10658 7364
rect 11974 7352 11980 7364
rect 12032 7392 12038 7404
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 12032 7364 12081 7392
rect 12032 7352 12038 7364
rect 12069 7361 12081 7364
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14918 7392 14924 7404
rect 14507 7364 14924 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7392 15347 7395
rect 15470 7392 15476 7404
rect 15335 7364 15476 7392
rect 15335 7361 15347 7364
rect 15289 7355 15347 7361
rect 15470 7352 15476 7364
rect 15528 7352 15534 7404
rect 4430 7324 4436 7336
rect 4391 7296 4436 7324
rect 4430 7284 4436 7296
rect 4488 7284 4494 7336
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8294 7324 8300 7336
rect 8159 7296 8300 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 15580 7333 15608 7432
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17681 7395 17739 7401
rect 17681 7392 17693 7395
rect 17083 7364 17693 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17681 7361 17693 7364
rect 17727 7392 17739 7395
rect 17865 7395 17923 7401
rect 17865 7392 17877 7395
rect 17727 7364 17877 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 17865 7361 17877 7364
rect 17911 7361 17923 7395
rect 17865 7355 17923 7361
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 13464 7296 14657 7324
rect 13464 7265 13492 7296
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7324 15623 7327
rect 15838 7324 15844 7336
rect 15611 7296 15844 7324
rect 15611 7293 15623 7296
rect 15565 7287 15623 7293
rect 15838 7284 15844 7296
rect 15896 7284 15902 7336
rect 16390 7324 16396 7336
rect 16351 7296 16396 7324
rect 16390 7284 16396 7296
rect 16448 7324 16454 7336
rect 17052 7324 17080 7355
rect 18046 7352 18052 7404
rect 18104 7392 18110 7404
rect 18233 7395 18291 7401
rect 18233 7392 18245 7395
rect 18104 7364 18245 7392
rect 18104 7352 18110 7364
rect 18233 7361 18245 7364
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 16448 7296 17080 7324
rect 17221 7327 17279 7333
rect 16448 7284 16454 7296
rect 17221 7293 17233 7327
rect 17267 7293 17279 7327
rect 17221 7287 17279 7293
rect 13449 7259 13507 7265
rect 13449 7225 13461 7259
rect 13495 7225 13507 7259
rect 13449 7219 13507 7225
rect 3099 7160 3372 7188
rect 3099 7157 3111 7160
rect 3053 7151 3111 7157
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 4212 7160 4537 7188
rect 4212 7148 4218 7160
rect 4525 7157 4537 7160
rect 4571 7188 4583 7191
rect 4982 7188 4988 7200
rect 4571 7160 4988 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 5997 7191 6055 7197
rect 5997 7188 6009 7191
rect 5224 7160 6009 7188
rect 5224 7148 5230 7160
rect 5997 7157 6009 7160
rect 6043 7157 6055 7191
rect 5997 7151 6055 7157
rect 6733 7191 6791 7197
rect 6733 7157 6745 7191
rect 6779 7188 6791 7191
rect 7466 7188 7472 7200
rect 6779 7160 7472 7188
rect 6779 7157 6791 7160
rect 6733 7151 6791 7157
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 9217 7191 9275 7197
rect 9217 7157 9229 7191
rect 9263 7188 9275 7191
rect 9398 7188 9404 7200
rect 9263 7160 9404 7188
rect 9263 7157 9275 7160
rect 9217 7151 9275 7157
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 13464 7188 13492 7219
rect 16206 7216 16212 7268
rect 16264 7256 16270 7268
rect 16669 7259 16727 7265
rect 16669 7256 16681 7259
rect 16264 7228 16681 7256
rect 16264 7216 16270 7228
rect 16669 7225 16681 7228
rect 16715 7225 16727 7259
rect 17236 7256 17264 7287
rect 16669 7219 16727 7225
rect 17144 7228 17264 7256
rect 17144 7200 17172 7228
rect 10284 7160 13492 7188
rect 10284 7148 10290 7160
rect 13814 7148 13820 7200
rect 13872 7188 13878 7200
rect 14093 7191 14151 7197
rect 14093 7188 14105 7191
rect 13872 7160 14105 7188
rect 13872 7148 13878 7160
rect 14093 7157 14105 7160
rect 14139 7157 14151 7191
rect 14093 7151 14151 7157
rect 17126 7148 17132 7200
rect 17184 7148 17190 7200
rect 18046 7188 18052 7200
rect 18007 7160 18052 7188
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 18414 7188 18420 7200
rect 18375 7160 18420 7188
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 1104 7098 18860 7120
rect 1104 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 3430 7098
rect 3482 7046 7622 7098
rect 7674 7046 7686 7098
rect 7738 7046 7750 7098
rect 7802 7046 7814 7098
rect 7866 7046 7878 7098
rect 7930 7046 12070 7098
rect 12122 7046 12134 7098
rect 12186 7046 12198 7098
rect 12250 7046 12262 7098
rect 12314 7046 12326 7098
rect 12378 7046 16518 7098
rect 16570 7046 16582 7098
rect 16634 7046 16646 7098
rect 16698 7046 16710 7098
rect 16762 7046 16774 7098
rect 16826 7046 18860 7098
rect 1104 7024 18860 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 1949 6987 2007 6993
rect 1949 6984 1961 6987
rect 1728 6956 1961 6984
rect 1728 6944 1734 6956
rect 1949 6953 1961 6956
rect 1995 6953 2007 6987
rect 1949 6947 2007 6953
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 5810 6984 5816 6996
rect 2280 6956 5672 6984
rect 5771 6956 5816 6984
rect 2280 6944 2286 6956
rect 1486 6876 1492 6928
rect 1544 6916 1550 6928
rect 5644 6916 5672 6956
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 11974 6944 11980 6996
rect 12032 6984 12038 6996
rect 15381 6987 15439 6993
rect 12032 6956 12664 6984
rect 12032 6944 12038 6956
rect 6270 6916 6276 6928
rect 1544 6888 4108 6916
rect 5644 6888 6276 6916
rect 1544 6876 1550 6888
rect 2424 6857 2452 6888
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2593 6851 2651 6857
rect 2455 6820 2489 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2593 6817 2605 6851
rect 2639 6848 2651 6851
rect 2869 6851 2927 6857
rect 2869 6848 2881 6851
rect 2639 6820 2881 6848
rect 2639 6817 2651 6820
rect 2593 6811 2651 6817
rect 2869 6817 2881 6820
rect 2915 6817 2927 6851
rect 2869 6811 2927 6817
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6780 1547 6783
rect 1857 6783 1915 6789
rect 1857 6780 1869 6783
rect 1535 6752 1869 6780
rect 1535 6749 1547 6752
rect 1489 6743 1547 6749
rect 1857 6749 1869 6752
rect 1903 6780 1915 6783
rect 1946 6780 1952 6792
rect 1903 6752 1952 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2608 6712 2636 6811
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 3970 6848 3976 6860
rect 3016 6820 3976 6848
rect 3016 6808 3022 6820
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 4080 6848 4108 6888
rect 6270 6876 6276 6888
rect 6328 6876 6334 6928
rect 12360 6857 12388 6956
rect 12437 6919 12495 6925
rect 12437 6885 12449 6919
rect 12483 6885 12495 6919
rect 12437 6879 12495 6885
rect 12345 6851 12403 6857
rect 4080 6820 4568 6848
rect 3145 6783 3203 6789
rect 2746 6752 3096 6780
rect 2746 6712 2774 6752
rect 2608 6684 2774 6712
rect 3068 6712 3096 6752
rect 3145 6749 3157 6783
rect 3191 6780 3203 6783
rect 3881 6783 3939 6789
rect 3881 6780 3893 6783
rect 3191 6752 3893 6780
rect 3191 6749 3203 6752
rect 3145 6743 3203 6749
rect 3881 6749 3893 6752
rect 3927 6780 3939 6783
rect 4246 6780 4252 6792
rect 3927 6752 4252 6780
rect 3927 6749 3939 6752
rect 3881 6743 3939 6749
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4430 6780 4436 6792
rect 4391 6752 4436 6780
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 4540 6780 4568 6820
rect 12345 6817 12357 6851
rect 12391 6817 12403 6851
rect 12345 6811 12403 6817
rect 6822 6780 6828 6792
rect 4540 6752 6828 6780
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 8444 6752 8493 6780
rect 8444 6740 8450 6752
rect 8481 6749 8493 6752
rect 8527 6780 8539 6783
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 8527 6752 9321 6780
rect 8527 6749 8539 6752
rect 8481 6743 8539 6749
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9565 6783 9623 6789
rect 9565 6780 9577 6783
rect 9456 6752 9577 6780
rect 9456 6740 9462 6752
rect 9565 6749 9577 6752
rect 9611 6749 9623 6783
rect 11330 6780 11336 6792
rect 9565 6743 9623 6749
rect 9692 6752 11336 6780
rect 3602 6712 3608 6724
rect 3068 6684 3608 6712
rect 3602 6672 3608 6684
rect 3660 6712 3666 6724
rect 4678 6715 4736 6721
rect 4678 6712 4690 6715
rect 3660 6684 4690 6712
rect 3660 6672 3666 6684
rect 4678 6681 4690 6684
rect 4724 6681 4736 6715
rect 4678 6675 4736 6681
rect 6178 6672 6184 6724
rect 6236 6712 6242 6724
rect 8236 6715 8294 6721
rect 8236 6712 8248 6715
rect 6236 6684 8248 6712
rect 6236 6672 6242 6684
rect 8236 6681 8248 6684
rect 8282 6712 8294 6715
rect 9692 6712 9720 6752
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 8282 6684 9720 6712
rect 10704 6684 11192 6712
rect 8282 6681 8294 6684
rect 8236 6675 8294 6681
rect 1578 6604 1584 6656
rect 1636 6644 1642 6656
rect 1673 6647 1731 6653
rect 1673 6644 1685 6647
rect 1636 6616 1685 6644
rect 1636 6604 1642 6616
rect 1673 6613 1685 6616
rect 1719 6613 1731 6647
rect 1673 6607 1731 6613
rect 2317 6647 2375 6653
rect 2317 6613 2329 6647
rect 2363 6644 2375 6647
rect 2958 6644 2964 6656
rect 2363 6616 2964 6644
rect 2363 6613 2375 6616
rect 2317 6607 2375 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 3142 6644 3148 6656
rect 3099 6616 3148 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 3510 6644 3516 6656
rect 3471 6616 3516 6644
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3970 6644 3976 6656
rect 3931 6616 3976 6644
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4249 6647 4307 6653
rect 4249 6613 4261 6647
rect 4295 6644 4307 6647
rect 4338 6644 4344 6656
rect 4295 6616 4344 6644
rect 4295 6613 4307 6616
rect 4249 6607 4307 6613
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 7098 6644 7104 6656
rect 7059 6616 7104 6644
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 10704 6653 10732 6684
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 10468 6616 10701 6644
rect 10468 6604 10474 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10689 6607 10747 6613
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 10965 6647 11023 6653
rect 10965 6644 10977 6647
rect 10836 6616 10977 6644
rect 10836 6604 10842 6616
rect 10965 6613 10977 6616
rect 11011 6613 11023 6647
rect 11164 6644 11192 6684
rect 11974 6672 11980 6724
rect 12032 6712 12038 6724
rect 12078 6715 12136 6721
rect 12078 6712 12090 6715
rect 12032 6684 12090 6712
rect 12032 6672 12038 6684
rect 12078 6681 12090 6684
rect 12124 6712 12136 6715
rect 12452 6712 12480 6879
rect 12636 6780 12664 6956
rect 15381 6953 15393 6987
rect 15427 6984 15439 6987
rect 15470 6984 15476 6996
rect 15427 6956 15476 6984
rect 15427 6953 15439 6956
rect 15381 6947 15439 6953
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 18138 6984 18144 6996
rect 18099 6956 18144 6984
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 14826 6916 14832 6928
rect 14752 6888 14832 6916
rect 14752 6857 14780 6888
rect 14826 6876 14832 6888
rect 14884 6876 14890 6928
rect 14737 6851 14795 6857
rect 14737 6817 14749 6851
rect 14783 6817 14795 6851
rect 14737 6811 14795 6817
rect 14921 6851 14979 6857
rect 14921 6817 14933 6851
rect 14967 6848 14979 6851
rect 15102 6848 15108 6860
rect 14967 6820 15108 6848
rect 14967 6817 14979 6820
rect 14921 6811 14979 6817
rect 15102 6808 15108 6820
rect 15160 6808 15166 6860
rect 16206 6848 16212 6860
rect 16167 6820 16212 6848
rect 16206 6808 16212 6820
rect 16264 6808 16270 6860
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6817 16359 6851
rect 17126 6848 17132 6860
rect 17087 6820 17132 6848
rect 16301 6811 16359 6817
rect 13817 6783 13875 6789
rect 13817 6780 13829 6783
rect 12636 6752 13829 6780
rect 13817 6749 13829 6752
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 16316 6780 16344 6811
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 17034 6780 17040 6792
rect 15528 6752 16344 6780
rect 16995 6752 17040 6780
rect 15528 6740 15534 6752
rect 17034 6740 17040 6752
rect 17092 6780 17098 6792
rect 17310 6780 17316 6792
rect 17092 6752 17316 6780
rect 17092 6740 17098 6752
rect 17310 6740 17316 6752
rect 17368 6780 17374 6792
rect 17405 6783 17463 6789
rect 17405 6780 17417 6783
rect 17368 6752 17417 6780
rect 17368 6740 17374 6752
rect 17405 6749 17417 6752
rect 17451 6749 17463 6783
rect 17405 6743 17463 6749
rect 13550 6715 13608 6721
rect 13550 6712 13562 6715
rect 12124 6684 12480 6712
rect 13004 6684 13562 6712
rect 12124 6681 12136 6684
rect 12078 6675 12136 6681
rect 13004 6644 13032 6684
rect 13550 6681 13562 6684
rect 13596 6681 13608 6715
rect 16022 6712 16028 6724
rect 13550 6675 13608 6681
rect 14016 6684 16028 6712
rect 11164 6616 13032 6644
rect 10965 6607 11023 6613
rect 13078 6604 13084 6656
rect 13136 6644 13142 6656
rect 14016 6644 14044 6684
rect 16022 6672 16028 6684
rect 16080 6672 16086 6724
rect 16117 6715 16175 6721
rect 16117 6681 16129 6715
rect 16163 6712 16175 6715
rect 16163 6684 16620 6712
rect 16163 6681 16175 6684
rect 16117 6675 16175 6681
rect 13136 6616 14044 6644
rect 13136 6604 13142 6616
rect 14090 6604 14096 6656
rect 14148 6644 14154 6656
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 14148 6616 14473 6644
rect 14148 6604 14154 6616
rect 14461 6613 14473 6616
rect 14507 6644 14519 6647
rect 14826 6644 14832 6656
rect 14507 6616 14832 6644
rect 14507 6613 14519 6616
rect 14461 6607 14519 6613
rect 14826 6604 14832 6616
rect 14884 6644 14890 6656
rect 15013 6647 15071 6653
rect 15013 6644 15025 6647
rect 14884 6616 15025 6644
rect 14884 6604 14890 6616
rect 15013 6613 15025 6616
rect 15059 6613 15071 6647
rect 15746 6644 15752 6656
rect 15707 6616 15752 6644
rect 15013 6607 15071 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 16592 6653 16620 6684
rect 16577 6647 16635 6653
rect 16577 6613 16589 6647
rect 16623 6613 16635 6647
rect 16942 6644 16948 6656
rect 16903 6616 16948 6644
rect 16577 6607 16635 6613
rect 16942 6604 16948 6616
rect 17000 6604 17006 6656
rect 1104 6554 18860 6576
rect 1104 6502 5398 6554
rect 5450 6502 5462 6554
rect 5514 6502 5526 6554
rect 5578 6502 5590 6554
rect 5642 6502 5654 6554
rect 5706 6502 9846 6554
rect 9898 6502 9910 6554
rect 9962 6502 9974 6554
rect 10026 6502 10038 6554
rect 10090 6502 10102 6554
rect 10154 6502 14294 6554
rect 14346 6502 14358 6554
rect 14410 6502 14422 6554
rect 14474 6502 14486 6554
rect 14538 6502 14550 6554
rect 14602 6502 18860 6554
rect 1104 6480 18860 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 3053 6443 3111 6449
rect 3053 6440 3065 6443
rect 2363 6412 3065 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 3053 6409 3065 6412
rect 3099 6409 3111 6443
rect 3053 6403 3111 6409
rect 3421 6443 3479 6449
rect 3421 6409 3433 6443
rect 3467 6440 3479 6443
rect 3881 6443 3939 6449
rect 3881 6440 3893 6443
rect 3467 6412 3893 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 3881 6409 3893 6412
rect 3927 6409 3939 6443
rect 4246 6440 4252 6452
rect 4159 6412 4252 6440
rect 3881 6403 3939 6409
rect 4246 6400 4252 6412
rect 4304 6440 4310 6452
rect 6546 6440 6552 6452
rect 4304 6412 6552 6440
rect 4304 6400 4310 6412
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 13078 6440 13084 6452
rect 6788 6412 13084 6440
rect 6788 6400 6794 6412
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 13262 6440 13268 6452
rect 13223 6412 13268 6440
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 14001 6443 14059 6449
rect 14001 6409 14013 6443
rect 14047 6440 14059 6443
rect 14369 6443 14427 6449
rect 14369 6440 14381 6443
rect 14047 6412 14381 6440
rect 14047 6409 14059 6412
rect 14001 6403 14059 6409
rect 14369 6409 14381 6412
rect 14415 6409 14427 6443
rect 14369 6403 14427 6409
rect 14829 6443 14887 6449
rect 14829 6409 14841 6443
rect 14875 6440 14887 6443
rect 15197 6443 15255 6449
rect 15197 6440 15209 6443
rect 14875 6412 15209 6440
rect 14875 6409 14887 6412
rect 14829 6403 14887 6409
rect 15197 6409 15209 6412
rect 15243 6409 15255 6443
rect 15197 6403 15255 6409
rect 16022 6400 16028 6452
rect 16080 6440 16086 6452
rect 16209 6443 16267 6449
rect 16209 6440 16221 6443
rect 16080 6412 16221 6440
rect 16080 6400 16086 6412
rect 16209 6409 16221 6412
rect 16255 6409 16267 6443
rect 16942 6440 16948 6452
rect 16903 6412 16948 6440
rect 16209 6403 16267 6409
rect 4430 6332 4436 6384
rect 4488 6372 4494 6384
rect 8294 6372 8300 6384
rect 4488 6344 6224 6372
rect 4488 6332 4494 6344
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 2222 6304 2228 6316
rect 2183 6276 2228 6304
rect 1765 6267 1823 6273
rect 1780 6236 1808 6267
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6304 3019 6307
rect 3786 6304 3792 6316
rect 3007 6276 3792 6304
rect 3007 6273 3019 6276
rect 2961 6267 3019 6273
rect 3786 6264 3792 6276
rect 3844 6304 3850 6316
rect 4062 6304 4068 6316
rect 3844 6276 4068 6304
rect 3844 6264 3850 6276
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 5626 6304 5632 6316
rect 4540 6276 5632 6304
rect 2406 6236 2412 6248
rect 1780 6208 2412 6236
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 2682 6236 2688 6248
rect 2547 6208 2688 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 2682 6196 2688 6208
rect 2740 6196 2746 6248
rect 2774 6196 2780 6248
rect 2832 6196 2838 6248
rect 3510 6236 3516 6248
rect 3471 6208 3516 6236
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 4154 6236 4160 6248
rect 3660 6208 4160 6236
rect 3660 6196 3666 6208
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 4338 6236 4344 6248
rect 4299 6208 4344 6236
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 4540 6245 4568 6276
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 5902 6264 5908 6316
rect 5960 6313 5966 6316
rect 6196 6313 6224 6344
rect 7576 6344 8300 6372
rect 5960 6304 5972 6313
rect 6181 6307 6239 6313
rect 5960 6276 6005 6304
rect 5960 6267 5972 6276
rect 6181 6273 6193 6307
rect 6227 6304 6239 6307
rect 7576 6304 7604 6344
rect 7944 6313 7972 6344
rect 8294 6332 8300 6344
rect 8352 6372 8358 6384
rect 12152 6375 12210 6381
rect 8352 6344 10272 6372
rect 8352 6332 8358 6344
rect 6227 6276 7604 6304
rect 7673 6307 7731 6313
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 7673 6273 7685 6307
rect 7719 6304 7731 6307
rect 7929 6307 7987 6313
rect 7719 6276 7880 6304
rect 7719 6273 7731 6276
rect 7673 6267 7731 6273
rect 5960 6264 5966 6267
rect 4525 6239 4583 6245
rect 4525 6205 4537 6239
rect 4571 6205 4583 6239
rect 4525 6199 4583 6205
rect 6457 6239 6515 6245
rect 6457 6205 6469 6239
rect 6503 6236 6515 6239
rect 6546 6236 6552 6248
rect 6503 6208 6552 6236
rect 6503 6205 6515 6208
rect 6457 6199 6515 6205
rect 2792 6168 2820 6196
rect 2958 6168 2964 6180
rect 2792 6140 2964 6168
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 4540 6168 4568 6199
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 7852 6236 7880 6276
rect 7929 6273 7941 6307
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 9973 6307 10031 6313
rect 9973 6273 9985 6307
rect 10019 6304 10031 6307
rect 10134 6304 10140 6316
rect 10019 6276 10140 6304
rect 10019 6273 10031 6276
rect 9973 6267 10031 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10244 6313 10272 6344
rect 12152 6341 12164 6375
rect 12198 6372 12210 6375
rect 12342 6372 12348 6384
rect 12198 6344 12348 6372
rect 12198 6341 12210 6344
rect 12152 6335 12210 6341
rect 12342 6332 12348 6344
rect 12400 6372 12406 6384
rect 12400 6332 12434 6372
rect 10229 6307 10287 6313
rect 10229 6273 10241 6307
rect 10275 6304 10287 6307
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 10275 6276 11897 6304
rect 10275 6273 10287 6276
rect 10229 6267 10287 6273
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 12406 6304 12434 6332
rect 13170 6304 13176 6316
rect 12406 6276 13176 6304
rect 11885 6267 11943 6273
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 13280 6304 13308 6400
rect 13909 6375 13967 6381
rect 13909 6341 13921 6375
rect 13955 6372 13967 6375
rect 15746 6372 15752 6384
rect 13955 6344 15752 6372
rect 13955 6341 13967 6344
rect 13909 6335 13967 6341
rect 15746 6332 15752 6344
rect 15804 6332 15810 6384
rect 16224 6372 16252 6403
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 16850 6372 16856 6384
rect 16224 6344 16856 6372
rect 16850 6332 16856 6344
rect 16908 6332 16914 6384
rect 14737 6307 14795 6313
rect 13280 6276 14263 6304
rect 7852 6208 8892 6236
rect 6730 6168 6736 6180
rect 4120 6140 4568 6168
rect 4632 6140 4936 6168
rect 4120 6128 4126 6140
rect 1857 6103 1915 6109
rect 1857 6069 1869 6103
rect 1903 6100 1915 6103
rect 1946 6100 1952 6112
rect 1903 6072 1952 6100
rect 1903 6069 1915 6072
rect 1857 6063 1915 6069
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 2832 6072 2877 6100
rect 2832 6060 2838 6072
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 4338 6100 4344 6112
rect 3200 6072 4344 6100
rect 3200 6060 3206 6072
rect 4338 6060 4344 6072
rect 4396 6100 4402 6112
rect 4632 6100 4660 6140
rect 4396 6072 4660 6100
rect 4396 6060 4402 6072
rect 4706 6060 4712 6112
rect 4764 6100 4770 6112
rect 4801 6103 4859 6109
rect 4801 6100 4813 6103
rect 4764 6072 4813 6100
rect 4764 6060 4770 6072
rect 4801 6069 4813 6072
rect 4847 6069 4859 6103
rect 4908 6100 4936 6140
rect 6196 6140 6736 6168
rect 5810 6100 5816 6112
rect 4908 6072 5816 6100
rect 4801 6063 4859 6069
rect 5810 6060 5816 6072
rect 5868 6100 5874 6112
rect 6196 6100 6224 6140
rect 6730 6128 6736 6140
rect 6788 6128 6794 6180
rect 8864 6112 8892 6208
rect 13446 6196 13452 6248
rect 13504 6236 13510 6248
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13504 6208 14105 6236
rect 13504 6196 13510 6208
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14235 6236 14263 6276
rect 14737 6273 14749 6307
rect 14783 6304 14795 6307
rect 15102 6304 15108 6316
rect 14783 6276 15108 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6304 15623 6307
rect 16390 6304 16396 6316
rect 15611 6276 16396 6304
rect 15611 6273 15623 6276
rect 15565 6267 15623 6273
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 14921 6239 14979 6245
rect 14921 6236 14933 6239
rect 14235 6208 14933 6236
rect 14093 6199 14151 6205
rect 14921 6205 14933 6208
rect 14967 6236 14979 6239
rect 15470 6236 15476 6248
rect 14967 6208 15476 6236
rect 14967 6205 14979 6208
rect 14921 6199 14979 6205
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 15654 6236 15660 6248
rect 15615 6208 15660 6236
rect 15654 6196 15660 6208
rect 15712 6196 15718 6248
rect 15746 6196 15752 6248
rect 15804 6236 15810 6248
rect 17126 6236 17132 6248
rect 15804 6208 17132 6236
rect 15804 6196 15810 6208
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 13078 6128 13084 6180
rect 13136 6168 13142 6180
rect 13541 6171 13599 6177
rect 13541 6168 13553 6171
rect 13136 6140 13553 6168
rect 13136 6128 13142 6140
rect 13541 6137 13553 6140
rect 13587 6137 13599 6171
rect 13541 6131 13599 6137
rect 14826 6128 14832 6180
rect 14884 6168 14890 6180
rect 18049 6171 18107 6177
rect 18049 6168 18061 6171
rect 14884 6140 18061 6168
rect 14884 6128 14890 6140
rect 18049 6137 18061 6140
rect 18095 6168 18107 6171
rect 18138 6168 18144 6180
rect 18095 6140 18144 6168
rect 18095 6137 18107 6140
rect 18049 6131 18107 6137
rect 18138 6128 18144 6140
rect 18196 6128 18202 6180
rect 5868 6072 6224 6100
rect 6549 6103 6607 6109
rect 5868 6060 5874 6072
rect 6549 6069 6561 6103
rect 6595 6100 6607 6103
rect 8018 6100 8024 6112
rect 6595 6072 8024 6100
rect 6595 6069 6607 6072
rect 6549 6063 6607 6069
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 8846 6100 8852 6112
rect 8807 6072 8852 6100
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 15194 6100 15200 6112
rect 13044 6072 15200 6100
rect 13044 6060 13050 6072
rect 15194 6060 15200 6072
rect 15252 6100 15258 6112
rect 16022 6100 16028 6112
rect 15252 6072 16028 6100
rect 15252 6060 15258 6072
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 1104 6010 18860 6032
rect 1104 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 3430 6010
rect 3482 5958 7622 6010
rect 7674 5958 7686 6010
rect 7738 5958 7750 6010
rect 7802 5958 7814 6010
rect 7866 5958 7878 6010
rect 7930 5958 12070 6010
rect 12122 5958 12134 6010
rect 12186 5958 12198 6010
rect 12250 5958 12262 6010
rect 12314 5958 12326 6010
rect 12378 5958 16518 6010
rect 16570 5958 16582 6010
rect 16634 5958 16646 6010
rect 16698 5958 16710 6010
rect 16762 5958 16774 6010
rect 16826 5958 18860 6010
rect 1104 5936 18860 5958
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 2823 5868 3464 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 2593 5831 2651 5837
rect 2593 5797 2605 5831
rect 2639 5828 2651 5831
rect 2958 5828 2964 5840
rect 2639 5800 2964 5828
rect 2639 5797 2651 5800
rect 2593 5791 2651 5797
rect 2958 5788 2964 5800
rect 3016 5828 3022 5840
rect 3142 5828 3148 5840
rect 3016 5800 3148 5828
rect 3016 5788 3022 5800
rect 3142 5788 3148 5800
rect 3200 5788 3206 5840
rect 3436 5828 3464 5868
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 3605 5899 3663 5905
rect 3605 5896 3617 5899
rect 3568 5868 3617 5896
rect 3568 5856 3574 5868
rect 3605 5865 3617 5868
rect 3651 5865 3663 5899
rect 3605 5859 3663 5865
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 3878 5896 3884 5908
rect 3752 5868 3884 5896
rect 3752 5856 3758 5868
rect 3878 5856 3884 5868
rect 3936 5896 3942 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3936 5868 4077 5896
rect 3936 5856 3942 5868
rect 4065 5865 4077 5868
rect 4111 5896 4123 5899
rect 4111 5868 5488 5896
rect 4111 5865 4123 5868
rect 4065 5859 4123 5865
rect 3786 5828 3792 5840
rect 3436 5800 3792 5828
rect 3786 5788 3792 5800
rect 3844 5788 3850 5840
rect 5460 5828 5488 5868
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 5905 5899 5963 5905
rect 5905 5896 5917 5899
rect 5776 5868 5917 5896
rect 5776 5856 5782 5868
rect 5905 5865 5917 5868
rect 5951 5896 5963 5899
rect 6178 5896 6184 5908
rect 5951 5868 6184 5896
rect 5951 5865 5963 5868
rect 5905 5859 5963 5865
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 14182 5896 14188 5908
rect 14143 5868 14188 5896
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 15102 5896 15108 5908
rect 15063 5868 15108 5896
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15565 5899 15623 5905
rect 15565 5865 15577 5899
rect 15611 5896 15623 5899
rect 15654 5896 15660 5908
rect 15611 5868 15660 5896
rect 15611 5865 15623 5868
rect 15565 5859 15623 5865
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 16390 5896 16396 5908
rect 16351 5868 16396 5896
rect 16390 5856 16396 5868
rect 16448 5856 16454 5908
rect 17494 5896 17500 5908
rect 17455 5868 17500 5896
rect 17494 5856 17500 5868
rect 17552 5856 17558 5908
rect 18046 5896 18052 5908
rect 18007 5868 18052 5896
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 6270 5828 6276 5840
rect 5460 5800 6276 5828
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 7374 5788 7380 5840
rect 7432 5828 7438 5840
rect 7837 5831 7895 5837
rect 7837 5828 7849 5831
rect 7432 5800 7849 5828
rect 7432 5788 7438 5800
rect 7837 5797 7849 5800
rect 7883 5828 7895 5831
rect 7929 5831 7987 5837
rect 7929 5828 7941 5831
rect 7883 5800 7941 5828
rect 7883 5797 7895 5800
rect 7837 5791 7895 5797
rect 7929 5797 7941 5800
rect 7975 5828 7987 5831
rect 8110 5828 8116 5840
rect 7975 5800 8116 5828
rect 7975 5797 7987 5800
rect 7929 5791 7987 5797
rect 8110 5788 8116 5800
rect 8168 5828 8174 5840
rect 8665 5831 8723 5837
rect 8665 5828 8677 5831
rect 8168 5800 8677 5828
rect 8168 5788 8174 5800
rect 8665 5797 8677 5800
rect 8711 5828 8723 5831
rect 9677 5831 9735 5837
rect 9677 5828 9689 5831
rect 8711 5800 9689 5828
rect 8711 5797 8723 5800
rect 8665 5791 8723 5797
rect 9677 5797 9689 5800
rect 9723 5828 9735 5831
rect 10137 5831 10195 5837
rect 10137 5828 10149 5831
rect 9723 5800 10149 5828
rect 9723 5797 9735 5800
rect 9677 5791 9735 5797
rect 10137 5797 10149 5800
rect 10183 5828 10195 5831
rect 10321 5831 10379 5837
rect 10321 5828 10333 5831
rect 10183 5800 10333 5828
rect 10183 5797 10195 5800
rect 10137 5791 10195 5797
rect 10321 5797 10333 5800
rect 10367 5797 10379 5831
rect 12986 5828 12992 5840
rect 10321 5791 10379 5797
rect 12406 5800 12992 5828
rect 1946 5760 1952 5772
rect 1907 5732 1952 5760
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 2133 5763 2191 5769
rect 2133 5729 2145 5763
rect 2179 5729 2191 5763
rect 2133 5723 2191 5729
rect 3053 5763 3111 5769
rect 3053 5729 3065 5763
rect 3099 5760 3111 5763
rect 4062 5760 4068 5772
rect 3099 5732 4068 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 1854 5692 1860 5704
rect 1815 5664 1860 5692
rect 1854 5652 1860 5664
rect 1912 5652 1918 5704
rect 2148 5692 2176 5723
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 4430 5720 4436 5772
rect 4488 5760 4494 5772
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 4488 5732 4537 5760
rect 4488 5720 4494 5732
rect 4525 5729 4537 5732
rect 4571 5729 4583 5763
rect 4525 5723 4583 5729
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 5960 5732 6745 5760
rect 5960 5720 5966 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 12406 5760 12434 5800
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 13170 5788 13176 5840
rect 13228 5828 13234 5840
rect 15746 5828 15752 5840
rect 13228 5800 15752 5828
rect 13228 5788 13234 5800
rect 6733 5723 6791 5729
rect 6840 5732 12434 5760
rect 12529 5763 12587 5769
rect 6086 5692 6092 5704
rect 2148 5664 6092 5692
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5692 6699 5695
rect 6840 5692 6868 5732
rect 12529 5729 12541 5763
rect 12575 5760 12587 5763
rect 12802 5760 12808 5772
rect 12575 5732 12808 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 12802 5720 12808 5732
rect 12860 5760 12866 5772
rect 14476 5769 14504 5800
rect 15746 5788 15752 5800
rect 15804 5788 15810 5840
rect 16298 5788 16304 5840
rect 16356 5828 16362 5840
rect 17221 5831 17279 5837
rect 17221 5828 17233 5831
rect 16356 5800 17233 5828
rect 16356 5788 16362 5800
rect 17221 5797 17233 5800
rect 17267 5797 17279 5831
rect 17221 5791 17279 5797
rect 13633 5763 13691 5769
rect 13633 5760 13645 5763
rect 12860 5732 13645 5760
rect 12860 5720 12866 5732
rect 13633 5729 13645 5732
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 14461 5763 14519 5769
rect 14461 5729 14473 5763
rect 14507 5729 14519 5763
rect 14461 5723 14519 5729
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5760 14703 5763
rect 15286 5760 15292 5772
rect 14691 5732 15292 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 16114 5760 16120 5772
rect 16075 5732 16120 5760
rect 16114 5720 16120 5732
rect 16172 5760 16178 5772
rect 16945 5763 17003 5769
rect 16945 5760 16957 5763
rect 16172 5732 16957 5760
rect 16172 5720 16178 5732
rect 16945 5729 16957 5732
rect 16991 5729 17003 5763
rect 16945 5723 17003 5729
rect 7466 5692 7472 5704
rect 6687 5664 6868 5692
rect 7427 5664 7472 5692
rect 6687 5661 6699 5664
rect 6641 5655 6699 5661
rect 3142 5624 3148 5636
rect 3055 5596 3148 5624
rect 3142 5584 3148 5596
rect 3200 5624 3206 5636
rect 3200 5596 4660 5624
rect 3200 5584 3206 5596
rect 1489 5559 1547 5565
rect 1489 5525 1501 5559
rect 1535 5556 1547 5559
rect 1670 5556 1676 5568
rect 1535 5528 1676 5556
rect 1535 5525 1547 5528
rect 1489 5519 1547 5525
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 2406 5556 2412 5568
rect 2367 5528 2412 5556
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 3694 5556 3700 5568
rect 3283 5528 3700 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 3881 5559 3939 5565
rect 3881 5525 3893 5559
rect 3927 5556 3939 5559
rect 4338 5556 4344 5568
rect 3927 5528 4344 5556
rect 3927 5525 3939 5528
rect 3881 5519 3939 5525
rect 4338 5516 4344 5528
rect 4396 5516 4402 5568
rect 4632 5556 4660 5596
rect 4706 5584 4712 5636
rect 4764 5633 4770 5636
rect 4764 5627 4828 5633
rect 4764 5593 4782 5627
rect 4816 5593 4828 5627
rect 4764 5587 4828 5593
rect 5997 5627 6055 5633
rect 5997 5593 6009 5627
rect 6043 5624 6055 5627
rect 6656 5624 6684 5655
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 9306 5692 9312 5704
rect 9267 5664 9312 5692
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5692 10747 5695
rect 11974 5692 11980 5704
rect 10735 5664 11980 5692
rect 10735 5661 10747 5664
rect 10689 5655 10747 5661
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 14182 5652 14188 5704
rect 14240 5692 14246 5704
rect 14734 5692 14740 5704
rect 14240 5664 14740 5692
rect 14240 5652 14246 5664
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 16022 5692 16028 5704
rect 15983 5664 16028 5692
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 16850 5692 16856 5704
rect 16811 5664 16856 5692
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 17494 5652 17500 5704
rect 17552 5652 17558 5704
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 17696 5664 17877 5692
rect 8205 5627 8263 5633
rect 8205 5624 8217 5627
rect 6043 5596 6684 5624
rect 6748 5596 8217 5624
rect 6043 5593 6055 5596
rect 5997 5587 6055 5593
rect 4764 5584 4770 5587
rect 6012 5556 6040 5587
rect 6178 5556 6184 5568
rect 4632 5528 6040 5556
rect 6139 5528 6184 5556
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 6270 5516 6276 5568
rect 6328 5556 6334 5568
rect 6549 5559 6607 5565
rect 6549 5556 6561 5559
rect 6328 5528 6561 5556
rect 6328 5516 6334 5528
rect 6549 5525 6561 5528
rect 6595 5556 6607 5559
rect 6748 5556 6776 5596
rect 8205 5593 8217 5596
rect 8251 5624 8263 5627
rect 11057 5627 11115 5633
rect 8251 5596 9352 5624
rect 8251 5593 8263 5596
rect 8205 5587 8263 5593
rect 7374 5556 7380 5568
rect 6595 5528 6776 5556
rect 7335 5528 7380 5556
rect 6595 5525 6607 5528
rect 6549 5519 6607 5525
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 9214 5556 9220 5568
rect 9175 5528 9220 5556
rect 9214 5516 9220 5528
rect 9272 5516 9278 5568
rect 9324 5556 9352 5596
rect 11057 5593 11069 5627
rect 11103 5624 11115 5627
rect 11238 5624 11244 5636
rect 11103 5596 11244 5624
rect 11103 5593 11115 5596
rect 11057 5587 11115 5593
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 12618 5584 12624 5636
rect 12676 5624 12682 5636
rect 12676 5596 12721 5624
rect 12676 5584 12682 5596
rect 13354 5584 13360 5636
rect 13412 5624 13418 5636
rect 13541 5627 13599 5633
rect 13541 5624 13553 5627
rect 13412 5596 13553 5624
rect 13412 5584 13418 5596
rect 13541 5593 13553 5596
rect 13587 5593 13599 5627
rect 15933 5627 15991 5633
rect 15933 5624 15945 5627
rect 13541 5587 13599 5593
rect 14936 5596 15945 5624
rect 14936 5556 14964 5596
rect 15933 5593 15945 5596
rect 15979 5624 15991 5627
rect 16298 5624 16304 5636
rect 15979 5596 16304 5624
rect 15979 5593 15991 5596
rect 15933 5587 15991 5593
rect 16298 5584 16304 5596
rect 16356 5584 16362 5636
rect 16761 5627 16819 5633
rect 16761 5593 16773 5627
rect 16807 5624 16819 5627
rect 17512 5624 17540 5652
rect 16807 5596 17540 5624
rect 16807 5593 16819 5596
rect 16761 5587 16819 5593
rect 9324 5528 14964 5556
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 15252 5528 15297 5556
rect 15252 5516 15258 5528
rect 17494 5516 17500 5568
rect 17552 5556 17558 5568
rect 17696 5565 17724 5664
rect 17865 5661 17877 5664
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 18138 5652 18144 5704
rect 18196 5692 18202 5704
rect 18233 5695 18291 5701
rect 18233 5692 18245 5695
rect 18196 5664 18245 5692
rect 18196 5652 18202 5664
rect 18233 5661 18245 5664
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 17681 5559 17739 5565
rect 17681 5556 17693 5559
rect 17552 5528 17693 5556
rect 17552 5516 17558 5528
rect 17681 5525 17693 5528
rect 17727 5525 17739 5559
rect 18414 5556 18420 5568
rect 18375 5528 18420 5556
rect 17681 5519 17739 5525
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 1104 5466 18860 5488
rect 1104 5414 5398 5466
rect 5450 5414 5462 5466
rect 5514 5414 5526 5466
rect 5578 5414 5590 5466
rect 5642 5414 5654 5466
rect 5706 5414 9846 5466
rect 9898 5414 9910 5466
rect 9962 5414 9974 5466
rect 10026 5414 10038 5466
rect 10090 5414 10102 5466
rect 10154 5414 14294 5466
rect 14346 5414 14358 5466
rect 14410 5414 14422 5466
rect 14474 5414 14486 5466
rect 14538 5414 14550 5466
rect 14602 5414 18860 5466
rect 1104 5392 18860 5414
rect 1765 5355 1823 5361
rect 1765 5321 1777 5355
rect 1811 5352 1823 5355
rect 1854 5352 1860 5364
rect 1811 5324 1860 5352
rect 1811 5321 1823 5324
rect 1765 5315 1823 5321
rect 1854 5312 1860 5324
rect 1912 5352 1918 5364
rect 2130 5352 2136 5364
rect 1912 5324 2136 5352
rect 1912 5312 1918 5324
rect 2130 5312 2136 5324
rect 2188 5312 2194 5364
rect 2222 5312 2228 5364
rect 2280 5352 2286 5364
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 2280 5324 2605 5352
rect 2280 5312 2286 5324
rect 2593 5321 2605 5324
rect 2639 5321 2651 5355
rect 2593 5315 2651 5321
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3513 5355 3571 5361
rect 3513 5352 3525 5355
rect 3099 5324 3525 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3513 5321 3525 5324
rect 3559 5321 3571 5355
rect 3513 5315 3571 5321
rect 3878 5312 3884 5364
rect 3936 5352 3942 5364
rect 3973 5355 4031 5361
rect 3973 5352 3985 5355
rect 3936 5324 3985 5352
rect 3936 5312 3942 5324
rect 3973 5321 3985 5324
rect 4019 5321 4031 5355
rect 3973 5315 4031 5321
rect 4893 5355 4951 5361
rect 4893 5321 4905 5355
rect 4939 5352 4951 5355
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 4939 5324 5365 5352
rect 4939 5321 4951 5324
rect 4893 5315 4951 5321
rect 5353 5321 5365 5324
rect 5399 5321 5411 5355
rect 5353 5315 5411 5321
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 6546 5352 6552 5364
rect 5767 5324 6552 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 4801 5287 4859 5293
rect 2240 5256 4752 5284
rect 2240 5225 2268 5256
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2225 5219 2283 5225
rect 2225 5216 2237 5219
rect 2179 5188 2237 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 2225 5185 2237 5188
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 2314 5176 2320 5228
rect 2372 5216 2378 5228
rect 2501 5219 2559 5225
rect 2501 5216 2513 5219
rect 2372 5188 2513 5216
rect 2372 5176 2378 5188
rect 2501 5185 2513 5188
rect 2547 5216 2559 5219
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 2547 5188 2973 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 2961 5185 2973 5188
rect 3007 5216 3019 5219
rect 3786 5216 3792 5228
rect 3007 5188 3792 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5185 3939 5219
rect 4724 5216 4752 5256
rect 4801 5253 4813 5287
rect 4847 5284 4859 5287
rect 6178 5284 6184 5296
rect 4847 5256 6184 5284
rect 4847 5253 4859 5256
rect 4801 5247 4859 5253
rect 6178 5244 6184 5256
rect 6236 5244 6242 5296
rect 6288 5216 6316 5324
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 6917 5355 6975 5361
rect 6917 5352 6929 5355
rect 6880 5324 6929 5352
rect 6880 5312 6886 5324
rect 6917 5321 6929 5324
rect 6963 5321 6975 5355
rect 6917 5315 6975 5321
rect 7653 5355 7711 5361
rect 7653 5321 7665 5355
rect 7699 5352 7711 5355
rect 11057 5355 11115 5361
rect 7699 5324 10180 5352
rect 7699 5321 7711 5324
rect 7653 5315 7711 5321
rect 7098 5244 7104 5296
rect 7156 5284 7162 5296
rect 7156 5256 7880 5284
rect 7156 5244 7162 5256
rect 4724 5188 6316 5216
rect 6825 5219 6883 5225
rect 3881 5179 3939 5185
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 7466 5216 7472 5228
rect 6871 5188 7472 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5148 3295 5151
rect 3602 5148 3608 5160
rect 3283 5120 3608 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 3602 5108 3608 5120
rect 3660 5108 3666 5160
rect 1946 5012 1952 5024
rect 1907 4984 1952 5012
rect 1946 4972 1952 4984
rect 2004 4972 2010 5024
rect 3896 5012 3924 5179
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4706 5148 4712 5160
rect 4120 5120 4165 5148
rect 4667 5120 4712 5148
rect 4120 5108 4126 5120
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 5810 5148 5816 5160
rect 5771 5120 5816 5148
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 5960 5120 6005 5148
rect 5960 5108 5966 5120
rect 6086 5108 6092 5160
rect 6144 5148 6150 5160
rect 6638 5148 6644 5160
rect 6144 5120 6644 5148
rect 6144 5108 6150 5120
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 7009 5151 7067 5157
rect 7009 5117 7021 5151
rect 7055 5117 7067 5151
rect 7009 5111 7067 5117
rect 5920 5080 5948 5108
rect 7024 5080 7052 5111
rect 7098 5108 7104 5160
rect 7156 5148 7162 5160
rect 7852 5157 7880 5256
rect 8110 5216 8116 5228
rect 8071 5188 8116 5216
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 8478 5216 8484 5228
rect 8439 5188 8484 5216
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 9398 5216 9404 5228
rect 9359 5188 9404 5216
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 7745 5151 7803 5157
rect 7745 5148 7757 5151
rect 7156 5120 7757 5148
rect 7156 5108 7162 5120
rect 7745 5117 7757 5120
rect 7791 5117 7803 5151
rect 7745 5111 7803 5117
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5117 7895 5151
rect 7837 5111 7895 5117
rect 5920 5052 7052 5080
rect 8128 5080 8156 5176
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 9582 5148 9588 5160
rect 8895 5120 9588 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 9732 5120 9777 5148
rect 9732 5108 9738 5120
rect 9033 5083 9091 5089
rect 9033 5080 9045 5083
rect 8128 5052 9045 5080
rect 9033 5049 9045 5052
rect 9079 5080 9091 5083
rect 9766 5080 9772 5092
rect 9079 5052 9772 5080
rect 9079 5049 9091 5052
rect 9033 5043 9091 5049
rect 9766 5040 9772 5052
rect 9824 5080 9830 5092
rect 9861 5083 9919 5089
rect 9861 5080 9873 5083
rect 9824 5052 9873 5080
rect 9824 5040 9830 5052
rect 9861 5049 9873 5052
rect 9907 5080 9919 5083
rect 10045 5083 10103 5089
rect 10045 5080 10057 5083
rect 9907 5052 10057 5080
rect 9907 5049 9919 5052
rect 9861 5043 9919 5049
rect 10045 5049 10057 5052
rect 10091 5049 10103 5083
rect 10152 5080 10180 5324
rect 11057 5321 11069 5355
rect 11103 5352 11115 5355
rect 11146 5352 11152 5364
rect 11103 5324 11152 5352
rect 11103 5321 11115 5324
rect 11057 5315 11115 5321
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 11287 5355 11345 5361
rect 11287 5321 11299 5355
rect 11333 5352 11345 5355
rect 12618 5352 12624 5364
rect 11333 5324 12624 5352
rect 11333 5321 11345 5324
rect 11287 5315 11345 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 13265 5355 13323 5361
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13633 5355 13691 5361
rect 13633 5352 13645 5355
rect 13311 5324 13645 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13633 5321 13645 5324
rect 13679 5321 13691 5355
rect 13633 5315 13691 5321
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 14001 5355 14059 5361
rect 14001 5352 14013 5355
rect 13780 5324 14013 5352
rect 13780 5312 13786 5324
rect 14001 5321 14013 5324
rect 14047 5321 14059 5355
rect 14001 5315 14059 5321
rect 14093 5355 14151 5361
rect 14093 5321 14105 5355
rect 14139 5352 14151 5355
rect 14366 5352 14372 5364
rect 14139 5324 14372 5352
rect 14139 5321 14151 5324
rect 14093 5315 14151 5321
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 14461 5355 14519 5361
rect 14461 5321 14473 5355
rect 14507 5321 14519 5355
rect 14461 5315 14519 5321
rect 14829 5355 14887 5361
rect 14829 5321 14841 5355
rect 14875 5352 14887 5355
rect 15194 5352 15200 5364
rect 14875 5324 15200 5352
rect 14875 5321 14887 5324
rect 14829 5315 14887 5321
rect 11164 5284 11192 5312
rect 11609 5287 11667 5293
rect 11609 5284 11621 5287
rect 11164 5256 11621 5284
rect 11609 5253 11621 5256
rect 11655 5253 11667 5287
rect 11609 5247 11667 5253
rect 11701 5287 11759 5293
rect 11701 5253 11713 5287
rect 11747 5284 11759 5287
rect 11790 5284 11796 5296
rect 11747 5256 11796 5284
rect 11747 5253 11759 5256
rect 11701 5247 11759 5253
rect 11790 5244 11796 5256
rect 11848 5244 11854 5296
rect 13173 5287 13231 5293
rect 13173 5253 13185 5287
rect 13219 5284 13231 5287
rect 14476 5284 14504 5315
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 15286 5312 15292 5364
rect 15344 5352 15350 5364
rect 17586 5352 17592 5364
rect 15344 5324 15389 5352
rect 17547 5324 17592 5352
rect 15344 5312 15350 5324
rect 17586 5312 17592 5324
rect 17644 5312 17650 5364
rect 13219 5256 14504 5284
rect 13219 5253 13231 5256
rect 13173 5247 13231 5253
rect 15378 5244 15384 5296
rect 15436 5284 15442 5296
rect 15657 5287 15715 5293
rect 15657 5284 15669 5287
rect 15436 5256 15669 5284
rect 15436 5244 15442 5256
rect 15657 5253 15669 5256
rect 15703 5253 15715 5287
rect 15657 5247 15715 5253
rect 16022 5244 16028 5296
rect 16080 5284 16086 5296
rect 16080 5256 16160 5284
rect 16080 5244 16086 5256
rect 10410 5216 10416 5228
rect 10371 5188 10416 5216
rect 10410 5176 10416 5188
rect 10468 5176 10474 5228
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11184 5219 11242 5225
rect 11184 5216 11196 5219
rect 11112 5188 11196 5216
rect 11112 5176 11118 5188
rect 11184 5185 11196 5188
rect 11230 5185 11242 5219
rect 15749 5219 15807 5225
rect 11184 5179 11242 5185
rect 12636 5188 13952 5216
rect 10781 5151 10839 5157
rect 10781 5117 10793 5151
rect 10827 5148 10839 5151
rect 11882 5148 11888 5160
rect 10827 5120 11888 5148
rect 10827 5117 10839 5120
rect 10781 5111 10839 5117
rect 11882 5108 11888 5120
rect 11940 5108 11946 5160
rect 12636 5157 12664 5188
rect 12621 5151 12679 5157
rect 12621 5117 12633 5151
rect 12667 5117 12679 5151
rect 12621 5111 12679 5117
rect 13357 5151 13415 5157
rect 13357 5117 13369 5151
rect 13403 5117 13415 5151
rect 13357 5111 13415 5117
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 10152 5052 12817 5080
rect 10045 5043 10103 5049
rect 12805 5049 12817 5052
rect 12851 5049 12863 5083
rect 12805 5043 12863 5049
rect 4430 5012 4436 5024
rect 3896 4984 4436 5012
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 5261 5015 5319 5021
rect 5261 4981 5273 5015
rect 5307 5012 5319 5015
rect 5718 5012 5724 5024
rect 5307 4984 5724 5012
rect 5307 4981 5319 4984
rect 5261 4975 5319 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6457 5015 6515 5021
rect 6457 4981 6469 5015
rect 6503 5012 6515 5015
rect 6730 5012 6736 5024
rect 6503 4984 6736 5012
rect 6503 4981 6515 4984
rect 6457 4975 6515 4981
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7285 5015 7343 5021
rect 7285 5012 7297 5015
rect 6972 4984 7297 5012
rect 6972 4972 6978 4984
rect 7285 4981 7297 4984
rect 7331 4981 7343 5015
rect 7285 4975 7343 4981
rect 11330 4972 11336 5024
rect 11388 5012 11394 5024
rect 13372 5012 13400 5111
rect 13924 5080 13952 5188
rect 14200 5188 15056 5216
rect 14200 5160 14228 5188
rect 14182 5148 14188 5160
rect 14143 5120 14188 5148
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 15028 5157 15056 5188
rect 15749 5185 15761 5219
rect 15795 5216 15807 5219
rect 15930 5216 15936 5228
rect 15795 5188 15936 5216
rect 15795 5185 15807 5188
rect 15749 5179 15807 5185
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16132 5225 16160 5256
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16206 5216 16212 5228
rect 16163 5188 16212 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16206 5176 16212 5188
rect 16264 5176 16270 5228
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 16850 5216 16856 5228
rect 16715 5188 16856 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 16850 5176 16856 5188
rect 16908 5216 16914 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16908 5188 17049 5216
rect 16908 5176 16914 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 17604 5216 17632 5312
rect 17773 5219 17831 5225
rect 17773 5216 17785 5219
rect 17604 5188 17785 5216
rect 17037 5179 17095 5185
rect 17773 5185 17785 5188
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 14921 5151 14979 5157
rect 14921 5117 14933 5151
rect 14967 5117 14979 5151
rect 14921 5111 14979 5117
rect 15013 5151 15071 5157
rect 15013 5117 15025 5151
rect 15059 5117 15071 5151
rect 15013 5111 15071 5117
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 16022 5148 16028 5160
rect 15887 5120 16028 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 14826 5080 14832 5092
rect 13924 5052 14832 5080
rect 14826 5040 14832 5052
rect 14884 5040 14890 5092
rect 14936 5080 14964 5111
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 15746 5080 15752 5092
rect 14936 5052 15752 5080
rect 11388 4984 13400 5012
rect 11388 4972 11394 4984
rect 13538 4972 13544 5024
rect 13596 5012 13602 5024
rect 14936 5012 14964 5052
rect 15746 5040 15752 5052
rect 15804 5040 15810 5092
rect 16298 5012 16304 5024
rect 13596 4984 14964 5012
rect 16259 4984 16304 5012
rect 13596 4972 13602 4984
rect 16298 4972 16304 4984
rect 16356 4972 16362 5024
rect 16850 5012 16856 5024
rect 16811 4984 16856 5012
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 17954 5012 17960 5024
rect 17915 4984 17960 5012
rect 17954 4972 17960 4984
rect 18012 4972 18018 5024
rect 1104 4922 18860 4944
rect 1104 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 3430 4922
rect 3482 4870 7622 4922
rect 7674 4870 7686 4922
rect 7738 4870 7750 4922
rect 7802 4870 7814 4922
rect 7866 4870 7878 4922
rect 7930 4870 12070 4922
rect 12122 4870 12134 4922
rect 12186 4870 12198 4922
rect 12250 4870 12262 4922
rect 12314 4870 12326 4922
rect 12378 4870 16518 4922
rect 16570 4870 16582 4922
rect 16634 4870 16646 4922
rect 16698 4870 16710 4922
rect 16762 4870 16774 4922
rect 16826 4870 18860 4922
rect 1104 4848 18860 4870
rect 2593 4811 2651 4817
rect 2593 4777 2605 4811
rect 2639 4808 2651 4811
rect 5261 4811 5319 4817
rect 2639 4780 4476 4808
rect 2639 4777 2651 4780
rect 2593 4771 2651 4777
rect 2222 4740 2228 4752
rect 2183 4712 2228 4740
rect 2222 4700 2228 4712
rect 2280 4700 2286 4752
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4604 1731 4607
rect 1854 4604 1860 4616
rect 1719 4576 1860 4604
rect 1719 4573 1731 4576
rect 1673 4567 1731 4573
rect 1854 4564 1860 4576
rect 1912 4564 1918 4616
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2608 4604 2636 4771
rect 4448 4752 4476 4780
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5810 4808 5816 4820
rect 5307 4780 5816 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 6181 4811 6239 4817
rect 6181 4777 6193 4811
rect 6227 4808 6239 4811
rect 7098 4808 7104 4820
rect 6227 4780 7104 4808
rect 6227 4777 6239 4780
rect 6181 4771 6239 4777
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 13538 4808 13544 4820
rect 7208 4780 13544 4808
rect 2777 4743 2835 4749
rect 2777 4709 2789 4743
rect 2823 4740 2835 4743
rect 3786 4740 3792 4752
rect 2823 4712 3792 4740
rect 2823 4709 2835 4712
rect 2777 4703 2835 4709
rect 3786 4700 3792 4712
rect 3844 4700 3850 4752
rect 4430 4700 4436 4752
rect 4488 4740 4494 4752
rect 7208 4740 7236 4780
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 13630 4768 13636 4820
rect 13688 4808 13694 4820
rect 14274 4808 14280 4820
rect 13688 4780 14280 4808
rect 13688 4768 13694 4780
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 14458 4768 14464 4820
rect 14516 4808 14522 4820
rect 14553 4811 14611 4817
rect 14553 4808 14565 4811
rect 14516 4780 14565 4808
rect 14516 4768 14522 4780
rect 14553 4777 14565 4780
rect 14599 4808 14611 4811
rect 14734 4808 14740 4820
rect 14599 4780 14740 4808
rect 14599 4777 14611 4780
rect 14553 4771 14611 4777
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 15746 4768 15752 4820
rect 15804 4808 15810 4820
rect 16117 4811 16175 4817
rect 16117 4808 16129 4811
rect 15804 4780 16129 4808
rect 15804 4768 15810 4780
rect 16117 4777 16129 4780
rect 16163 4777 16175 4811
rect 16117 4771 16175 4777
rect 16206 4768 16212 4820
rect 16264 4808 16270 4820
rect 16301 4811 16359 4817
rect 16301 4808 16313 4811
rect 16264 4780 16313 4808
rect 16264 4768 16270 4780
rect 16301 4777 16313 4780
rect 16347 4777 16359 4811
rect 16301 4771 16359 4777
rect 14090 4740 14096 4752
rect 4488 4712 7236 4740
rect 7300 4712 14096 4740
rect 4488 4700 4494 4712
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4672 3203 4675
rect 3694 4672 3700 4684
rect 3191 4644 3700 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 2455 4576 2636 4604
rect 2961 4607 3019 4613
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2961 4573 2973 4607
rect 3007 4604 3019 4607
rect 3160 4604 3188 4635
rect 3694 4632 3700 4644
rect 3752 4632 3758 4684
rect 5534 4672 5540 4684
rect 5495 4644 5540 4672
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 5718 4672 5724 4684
rect 5679 4644 5724 4672
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 6730 4672 6736 4684
rect 6691 4644 6736 4672
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4672 6883 4675
rect 7300 4672 7328 4712
rect 14090 4700 14096 4712
rect 14148 4700 14154 4752
rect 15378 4700 15384 4752
rect 15436 4740 15442 4752
rect 16485 4743 16543 4749
rect 16485 4740 16497 4743
rect 15436 4712 16497 4740
rect 15436 4700 15442 4712
rect 16485 4709 16497 4712
rect 16531 4709 16543 4743
rect 16485 4703 16543 4709
rect 6871 4644 7328 4672
rect 7377 4675 7435 4681
rect 6871 4641 6883 4644
rect 6825 4635 6883 4641
rect 7377 4641 7389 4675
rect 7423 4672 7435 4675
rect 7466 4672 7472 4684
rect 7423 4644 7472 4672
rect 7423 4641 7435 4644
rect 7377 4635 7435 4641
rect 3007 4576 3188 4604
rect 3421 4607 3479 4613
rect 3007 4573 3019 4576
rect 2961 4567 3019 4573
rect 3421 4573 3433 4607
rect 3467 4604 3479 4607
rect 3878 4604 3884 4616
rect 3467 4576 3884 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 1578 4428 1584 4480
rect 1636 4468 1642 4480
rect 1857 4471 1915 4477
rect 1857 4468 1869 4471
rect 1636 4440 1869 4468
rect 1636 4428 1642 4440
rect 1857 4437 1869 4440
rect 1903 4437 1915 4471
rect 2056 4468 2084 4567
rect 3878 4564 3884 4576
rect 3936 4564 3942 4616
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 6840 4604 6868 4635
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 9677 4675 9735 4681
rect 8076 4644 9352 4672
rect 8076 4632 8082 4644
rect 4764 4576 6868 4604
rect 4764 4564 4770 4576
rect 9214 4564 9220 4616
rect 9272 4564 9278 4616
rect 9324 4613 9352 4644
rect 9677 4641 9689 4675
rect 9723 4672 9735 4675
rect 9766 4672 9772 4684
rect 9723 4644 9772 4672
rect 9723 4641 9735 4644
rect 9677 4635 9735 4641
rect 9766 4632 9772 4644
rect 9824 4672 9830 4684
rect 9861 4675 9919 4681
rect 9861 4672 9873 4675
rect 9824 4644 9873 4672
rect 9824 4632 9830 4644
rect 9861 4641 9873 4644
rect 9907 4672 9919 4675
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 9907 4644 10057 4672
rect 9907 4641 9919 4644
rect 9861 4635 9919 4641
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 10778 4672 10784 4684
rect 10045 4635 10103 4641
rect 10428 4644 10784 4672
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 10428 4613 10456 4644
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 10962 4672 10968 4684
rect 10923 4644 10968 4672
rect 10962 4632 10968 4644
rect 11020 4672 11026 4684
rect 12066 4672 12072 4684
rect 11020 4644 12072 4672
rect 11020 4632 11026 4644
rect 12066 4632 12072 4644
rect 12124 4632 12130 4684
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4672 12311 4675
rect 12526 4672 12532 4684
rect 12299 4644 12532 4672
rect 12299 4641 12311 4644
rect 12253 4635 12311 4641
rect 12526 4632 12532 4644
rect 12584 4672 12590 4684
rect 13265 4675 13323 4681
rect 12584 4644 13124 4672
rect 12584 4632 12590 4644
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 10284 4576 10425 4604
rect 10284 4564 10290 4576
rect 10413 4573 10425 4576
rect 10459 4573 10471 4607
rect 10413 4567 10471 4573
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 13096 4604 13124 4644
rect 13265 4641 13277 4675
rect 13311 4672 13323 4675
rect 14235 4672 14366 4684
rect 17402 4672 17408 4684
rect 13311 4656 17408 4672
rect 13311 4644 14263 4656
rect 14338 4644 17408 4656
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 17402 4632 17408 4644
rect 17460 4632 17466 4684
rect 13633 4607 13691 4613
rect 13633 4604 13645 4607
rect 11940 4576 12112 4604
rect 13096 4576 13645 4604
rect 11940 4564 11946 4576
rect 5813 4539 5871 4545
rect 5813 4505 5825 4539
rect 5859 4536 5871 4539
rect 8021 4539 8079 4545
rect 5859 4508 6316 4536
rect 5859 4505 5871 4508
rect 5813 4499 5871 4505
rect 3605 4471 3663 4477
rect 3605 4468 3617 4471
rect 2056 4440 3617 4468
rect 1857 4431 1915 4437
rect 3605 4437 3617 4440
rect 3651 4468 3663 4471
rect 6086 4468 6092 4480
rect 3651 4440 6092 4468
rect 3651 4437 3663 4440
rect 3605 4431 3663 4437
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 6288 4477 6316 4508
rect 8021 4505 8033 4539
rect 8067 4536 8079 4539
rect 8110 4536 8116 4548
rect 8067 4508 8116 4536
rect 8067 4505 8079 4508
rect 8021 4499 8079 4505
rect 8110 4496 8116 4508
rect 8168 4536 8174 4548
rect 8481 4539 8539 4545
rect 8481 4536 8493 4539
rect 8168 4508 8493 4536
rect 8168 4496 8174 4508
rect 8481 4505 8493 4508
rect 8527 4536 8539 4539
rect 8665 4539 8723 4545
rect 8665 4536 8677 4539
rect 8527 4508 8677 4536
rect 8527 4505 8539 4508
rect 8481 4499 8539 4505
rect 8665 4505 8677 4508
rect 8711 4505 8723 4539
rect 9232 4536 9260 4564
rect 10778 4536 10784 4548
rect 9232 4508 10640 4536
rect 10739 4508 10784 4536
rect 8665 4499 8723 4505
rect 6273 4471 6331 4477
rect 6273 4437 6285 4471
rect 6319 4437 6331 4471
rect 6638 4468 6644 4480
rect 6599 4440 6644 4468
rect 6273 4431 6331 4437
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 7193 4471 7251 4477
rect 7193 4468 7205 4471
rect 6880 4440 7205 4468
rect 6880 4428 6886 4440
rect 7193 4437 7205 4440
rect 7239 4468 7251 4471
rect 8202 4468 8208 4480
rect 7239 4440 8208 4468
rect 7239 4437 7251 4440
rect 7193 4431 7251 4437
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 9122 4428 9128 4480
rect 9180 4468 9186 4480
rect 9217 4471 9275 4477
rect 9217 4468 9229 4471
rect 9180 4440 9229 4468
rect 9180 4428 9186 4440
rect 9217 4437 9229 4440
rect 9263 4437 9275 4471
rect 10612 4468 10640 4508
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 11054 4496 11060 4548
rect 11112 4536 11118 4548
rect 11977 4539 12035 4545
rect 11112 4508 11205 4536
rect 11112 4496 11118 4508
rect 11977 4505 11989 4539
rect 12023 4505 12035 4539
rect 12084 4536 12112 4576
rect 13633 4573 13645 4576
rect 13679 4573 13691 4607
rect 13633 4567 13691 4573
rect 14274 4564 14280 4616
rect 14332 4604 14338 4616
rect 15930 4604 15936 4616
rect 14332 4576 14688 4604
rect 15891 4576 15936 4604
rect 14332 4564 14338 4576
rect 12345 4539 12403 4545
rect 12345 4536 12357 4539
rect 12084 4508 12357 4536
rect 11977 4499 12035 4505
rect 12345 4505 12357 4508
rect 12391 4505 12403 4539
rect 14660 4536 14688 4576
rect 15930 4564 15936 4576
rect 15988 4604 15994 4616
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 15988 4576 17509 4604
rect 15988 4564 15994 4576
rect 17497 4573 17509 4576
rect 17543 4604 17555 4607
rect 17681 4607 17739 4613
rect 17681 4604 17693 4607
rect 17543 4576 17693 4604
rect 17543 4573 17555 4576
rect 17497 4567 17555 4573
rect 17681 4573 17693 4576
rect 17727 4573 17739 4607
rect 17681 4567 17739 4573
rect 14829 4539 14887 4545
rect 14829 4536 14841 4539
rect 12345 4499 12403 4505
rect 13372 4508 14596 4536
rect 14660 4508 14841 4536
rect 11072 4468 11100 4496
rect 10612 4440 11100 4468
rect 9217 4431 9275 4437
rect 11146 4428 11152 4480
rect 11204 4468 11210 4480
rect 11790 4468 11796 4480
rect 11204 4440 11796 4468
rect 11204 4428 11210 4440
rect 11790 4428 11796 4440
rect 11848 4428 11854 4480
rect 11992 4468 12020 4499
rect 13372 4468 13400 4508
rect 11992 4440 13400 4468
rect 13541 4471 13599 4477
rect 13541 4437 13553 4471
rect 13587 4468 13599 4471
rect 13722 4468 13728 4480
rect 13587 4440 13728 4468
rect 13587 4437 13599 4440
rect 13541 4431 13599 4437
rect 13722 4428 13728 4440
rect 13780 4428 13786 4480
rect 14568 4468 14596 4508
rect 14829 4505 14841 4508
rect 14875 4505 14887 4539
rect 14829 4499 14887 4505
rect 14918 4496 14924 4548
rect 14976 4536 14982 4548
rect 15841 4539 15899 4545
rect 14976 4508 15021 4536
rect 14976 4496 14982 4508
rect 15841 4505 15853 4539
rect 15887 4536 15899 4539
rect 17126 4536 17132 4548
rect 15887 4508 17132 4536
rect 15887 4505 15899 4508
rect 15841 4499 15899 4505
rect 17126 4496 17132 4508
rect 17184 4496 17190 4548
rect 16022 4468 16028 4480
rect 14568 4440 16028 4468
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 17770 4428 17776 4480
rect 17828 4468 17834 4480
rect 17865 4471 17923 4477
rect 17865 4468 17877 4471
rect 17828 4440 17877 4468
rect 17828 4428 17834 4440
rect 17865 4437 17877 4440
rect 17911 4437 17923 4471
rect 17865 4431 17923 4437
rect 1104 4378 18860 4400
rect 1104 4326 5398 4378
rect 5450 4326 5462 4378
rect 5514 4326 5526 4378
rect 5578 4326 5590 4378
rect 5642 4326 5654 4378
rect 5706 4326 9846 4378
rect 9898 4326 9910 4378
rect 9962 4326 9974 4378
rect 10026 4326 10038 4378
rect 10090 4326 10102 4378
rect 10154 4326 14294 4378
rect 14346 4326 14358 4378
rect 14410 4326 14422 4378
rect 14474 4326 14486 4378
rect 14538 4326 14550 4378
rect 14602 4326 18860 4378
rect 1104 4304 18860 4326
rect 5902 4224 5908 4276
rect 5960 4264 5966 4276
rect 6089 4267 6147 4273
rect 6089 4264 6101 4267
rect 5960 4236 6101 4264
rect 5960 4224 5966 4236
rect 6089 4233 6101 4236
rect 6135 4233 6147 4267
rect 6089 4227 6147 4233
rect 6457 4267 6515 4273
rect 6457 4233 6469 4267
rect 6503 4264 6515 4267
rect 6546 4264 6552 4276
rect 6503 4236 6552 4264
rect 6503 4233 6515 4236
rect 6457 4227 6515 4233
rect 6104 4196 6132 4227
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 8021 4267 8079 4273
rect 8021 4233 8033 4267
rect 8067 4264 8079 4267
rect 8110 4264 8116 4276
rect 8067 4236 8116 4264
rect 8067 4233 8079 4236
rect 8021 4227 8079 4233
rect 8110 4224 8116 4236
rect 8168 4224 8174 4276
rect 8202 4224 8208 4276
rect 8260 4264 8266 4276
rect 11054 4264 11060 4276
rect 8260 4236 11060 4264
rect 8260 4224 8266 4236
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 14550 4264 14556 4276
rect 11256 4236 14556 4264
rect 6638 4196 6644 4208
rect 6104 4168 6644 4196
rect 6638 4156 6644 4168
rect 6696 4156 6702 4208
rect 1670 4128 1676 4140
rect 1631 4100 1676 4128
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4097 2559 4131
rect 2501 4091 2559 4097
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3050 4128 3056 4140
rect 2915 4100 3056 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 1854 4060 1860 4072
rect 1815 4032 1860 4060
rect 1854 4020 1860 4032
rect 1912 4020 1918 4072
rect 2516 4060 2544 4091
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 3234 4128 3240 4140
rect 3195 4100 3240 4128
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 8128 4128 8156 4224
rect 9122 4196 9128 4208
rect 9083 4168 9128 4196
rect 9122 4156 9128 4168
rect 9180 4156 9186 4208
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 11256 4205 11284 4236
rect 14550 4224 14556 4236
rect 14608 4224 14614 4276
rect 14642 4224 14648 4276
rect 14700 4264 14706 4276
rect 14700 4236 15884 4264
rect 14700 4224 14706 4236
rect 10321 4199 10379 4205
rect 10321 4196 10333 4199
rect 9640 4168 10333 4196
rect 9640 4156 9646 4168
rect 10321 4165 10333 4168
rect 10367 4165 10379 4199
rect 10321 4159 10379 4165
rect 11241 4199 11299 4205
rect 11241 4165 11253 4199
rect 11287 4165 11299 4199
rect 11241 4159 11299 4165
rect 11698 4156 11704 4208
rect 11756 4196 11762 4208
rect 12526 4196 12532 4208
rect 11756 4168 12296 4196
rect 12487 4168 12532 4196
rect 11756 4156 11762 4168
rect 8481 4131 8539 4137
rect 8128 4100 8432 4128
rect 3252 4060 3280 4088
rect 8110 4060 8116 4072
rect 2516 4032 3280 4060
rect 8071 4032 8116 4060
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 8404 4060 8432 4100
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 8846 4128 8852 4140
rect 8527 4100 8852 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 9030 4060 9036 4072
rect 8404 4032 8892 4060
rect 8991 4032 9036 4060
rect 2314 3992 2320 4004
rect 2275 3964 2320 3992
rect 2314 3952 2320 3964
rect 2372 3952 2378 4004
rect 5718 3952 5724 4004
rect 5776 3992 5782 4004
rect 8864 4001 8892 4032
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 10042 4060 10048 4072
rect 10003 4032 10048 4060
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 10318 4060 10324 4072
rect 10275 4032 10324 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10318 4020 10324 4032
rect 10376 4020 10382 4072
rect 11698 4020 11704 4072
rect 11756 4060 11762 4072
rect 11885 4063 11943 4069
rect 11885 4060 11897 4063
rect 11756 4032 11897 4060
rect 11756 4020 11762 4032
rect 11885 4029 11897 4032
rect 11931 4029 11943 4063
rect 12066 4060 12072 4072
rect 12027 4032 12072 4060
rect 11885 4023 11943 4029
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 12268 4060 12296 4168
rect 12526 4156 12532 4168
rect 12584 4156 12590 4208
rect 14783 4199 14841 4205
rect 14783 4165 14795 4199
rect 14829 4196 14841 4199
rect 15105 4199 15163 4205
rect 15105 4196 15117 4199
rect 14829 4168 15117 4196
rect 14829 4165 14841 4168
rect 14783 4159 14841 4165
rect 15105 4165 15117 4168
rect 15151 4165 15163 4199
rect 15105 4159 15163 4165
rect 14680 4130 14738 4136
rect 14680 4096 14692 4130
rect 14726 4096 14738 4130
rect 15856 4128 15884 4236
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 15856 4100 17693 4128
rect 14680 4090 14738 4096
rect 17681 4097 17693 4100
rect 17727 4128 17739 4131
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 17727 4100 17785 4128
rect 17727 4097 17739 4100
rect 17681 4091 17739 4097
rect 17773 4097 17785 4100
rect 17819 4097 17831 4131
rect 17773 4091 17831 4097
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12268 4032 12449 4060
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 13446 4060 13452 4072
rect 13407 4032 13452 4060
rect 12437 4023 12495 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 14695 4060 14723 4090
rect 15013 4063 15071 4069
rect 15013 4060 15025 4063
rect 14476 4032 14723 4060
rect 14752 4032 15025 4060
rect 8849 3995 8907 4001
rect 5776 3964 8800 3992
rect 5776 3952 5782 3964
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 2866 3924 2872 3936
rect 2731 3896 2872 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 8772 3924 8800 3964
rect 8849 3961 8861 3995
rect 8895 3961 8907 3995
rect 8849 3955 8907 3961
rect 10226 3924 10232 3936
rect 8772 3896 10232 3924
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10336 3924 10364 4020
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 10836 3964 12121 3992
rect 10836 3952 10842 3964
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 10336 3896 11529 3924
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 12093 3924 12121 3964
rect 14476 3936 14504 4032
rect 14752 3936 14780 4032
rect 15013 4029 15025 4032
rect 15059 4029 15071 4063
rect 15562 4060 15568 4072
rect 15523 4032 15568 4060
rect 15013 4023 15071 4029
rect 15562 4020 15568 4032
rect 15620 4020 15626 4072
rect 14458 3924 14464 3936
rect 12093 3896 14464 3924
rect 11517 3887 11575 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 14553 3927 14611 3933
rect 14553 3893 14565 3927
rect 14599 3924 14611 3927
rect 14734 3924 14740 3936
rect 14599 3896 14740 3924
rect 14599 3893 14611 3896
rect 14553 3887 14611 3893
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 17954 3924 17960 3936
rect 17915 3896 17960 3924
rect 17954 3884 17960 3896
rect 18012 3884 18018 3936
rect 1104 3834 18860 3856
rect 1104 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 3430 3834
rect 3482 3782 7622 3834
rect 7674 3782 7686 3834
rect 7738 3782 7750 3834
rect 7802 3782 7814 3834
rect 7866 3782 7878 3834
rect 7930 3782 12070 3834
rect 12122 3782 12134 3834
rect 12186 3782 12198 3834
rect 12250 3782 12262 3834
rect 12314 3782 12326 3834
rect 12378 3782 16518 3834
rect 16570 3782 16582 3834
rect 16634 3782 16646 3834
rect 16698 3782 16710 3834
rect 16762 3782 16774 3834
rect 16826 3782 18860 3834
rect 1104 3760 18860 3782
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 8202 3720 8208 3732
rect 3476 3692 8208 3720
rect 3476 3680 3482 3692
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 8938 3720 8944 3732
rect 8899 3692 8944 3720
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 10137 3723 10195 3729
rect 10137 3720 10149 3723
rect 9088 3692 10149 3720
rect 9088 3680 9094 3692
rect 10137 3689 10149 3692
rect 10183 3689 10195 3723
rect 10137 3683 10195 3689
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 14918 3720 14924 3732
rect 14148 3692 14924 3720
rect 14148 3680 14154 3692
rect 14918 3680 14924 3692
rect 14976 3680 14982 3732
rect 15746 3720 15752 3732
rect 15707 3692 15752 3720
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 8956 3652 8984 3680
rect 7760 3624 8984 3652
rect 2777 3587 2835 3593
rect 2777 3584 2789 3587
rect 2148 3556 2789 3584
rect 2148 3525 2176 3556
rect 2777 3553 2789 3556
rect 2823 3584 2835 3587
rect 7282 3584 7288 3596
rect 2823 3556 7288 3584
rect 2823 3553 2835 3556
rect 2777 3547 2835 3553
rect 7282 3544 7288 3556
rect 7340 3544 7346 3596
rect 7760 3593 7788 3624
rect 10042 3612 10048 3664
rect 10100 3652 10106 3664
rect 15470 3652 15476 3664
rect 10100 3624 15476 3652
rect 10100 3612 10106 3624
rect 15470 3612 15476 3624
rect 15528 3612 15534 3664
rect 7745 3587 7803 3593
rect 7745 3553 7757 3587
rect 7791 3553 7803 3587
rect 7745 3547 7803 3553
rect 8757 3587 8815 3593
rect 8757 3553 8769 3587
rect 8803 3584 8815 3587
rect 12986 3584 12992 3596
rect 8803 3556 12992 3584
rect 8803 3553 8815 3556
rect 8757 3547 8815 3553
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 13354 3544 13360 3596
rect 13412 3584 13418 3596
rect 14185 3587 14243 3593
rect 14185 3584 14197 3587
rect 13412 3556 14197 3584
rect 13412 3544 13418 3556
rect 14185 3553 14197 3556
rect 14231 3553 14243 3587
rect 15010 3584 15016 3596
rect 14971 3556 15016 3584
rect 14185 3547 14243 3553
rect 15010 3544 15016 3556
rect 15068 3544 15074 3596
rect 15764 3584 15792 3680
rect 16025 3587 16083 3593
rect 16025 3584 16037 3587
rect 15764 3556 16037 3584
rect 16025 3553 16037 3556
rect 16071 3553 16083 3587
rect 16025 3547 16083 3553
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3516 2559 3519
rect 2682 3516 2688 3528
rect 2547 3488 2688 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3516 5871 3519
rect 6914 3516 6920 3528
rect 5859 3488 6920 3516
rect 5859 3485 5871 3488
rect 5813 3479 5871 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7444 3519 7502 3525
rect 7444 3485 7456 3519
rect 7490 3516 7502 3519
rect 7490 3488 7604 3516
rect 7490 3485 7502 3488
rect 7444 3479 7502 3485
rect 1857 3451 1915 3457
rect 1857 3417 1869 3451
rect 1903 3448 1915 3451
rect 2866 3448 2872 3460
rect 1903 3420 2872 3448
rect 1903 3417 1915 3420
rect 1857 3411 1915 3417
rect 2866 3408 2872 3420
rect 2924 3408 2930 3460
rect 3050 3408 3056 3460
rect 3108 3448 3114 3460
rect 5537 3451 5595 3457
rect 5537 3448 5549 3451
rect 3108 3420 5549 3448
rect 3108 3408 3114 3420
rect 5537 3417 5549 3420
rect 5583 3417 5595 3451
rect 7576 3448 7604 3488
rect 9122 3476 9128 3528
rect 9180 3525 9186 3528
rect 9180 3519 9218 3525
rect 9206 3485 9218 3519
rect 9180 3479 9218 3485
rect 9180 3476 9186 3479
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 10908 3519 10966 3525
rect 10908 3516 10920 3519
rect 9640 3488 10920 3516
rect 9640 3476 9646 3488
rect 10908 3485 10920 3488
rect 10954 3485 10966 3519
rect 10908 3479 10966 3485
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 11882 3516 11888 3528
rect 11296 3488 11888 3516
rect 11296 3476 11302 3488
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 12526 3476 12532 3528
rect 12584 3516 12590 3528
rect 13116 3519 13174 3525
rect 13116 3516 13128 3519
rect 12584 3488 13128 3516
rect 12584 3476 12590 3488
rect 13116 3485 13128 3488
rect 13162 3485 13174 3519
rect 13116 3479 13174 3485
rect 7837 3451 7895 3457
rect 7576 3420 7696 3448
rect 5537 3411 5595 3417
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 7558 3389 7564 3392
rect 2317 3383 2375 3389
rect 2317 3380 2329 3383
rect 1452 3352 2329 3380
rect 1452 3340 1458 3352
rect 2317 3349 2329 3352
rect 2363 3349 2375 3383
rect 2317 3343 2375 3349
rect 7515 3383 7564 3389
rect 7515 3349 7527 3383
rect 7561 3349 7564 3383
rect 7515 3343 7564 3349
rect 7558 3340 7564 3343
rect 7616 3340 7622 3392
rect 7668 3380 7696 3420
rect 7837 3417 7849 3451
rect 7883 3448 7895 3451
rect 8110 3448 8116 3460
rect 7883 3420 8116 3448
rect 7883 3417 7895 3420
rect 7837 3411 7895 3417
rect 7852 3380 7880 3411
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 11606 3408 11612 3460
rect 11664 3448 11670 3460
rect 12713 3451 12771 3457
rect 12713 3448 12725 3451
rect 11664 3420 12725 3448
rect 11664 3408 11670 3420
rect 12713 3417 12725 3420
rect 12759 3417 12771 3451
rect 12713 3411 12771 3417
rect 13219 3451 13277 3457
rect 13219 3417 13231 3451
rect 13265 3448 13277 3451
rect 14277 3451 14335 3457
rect 13265 3420 14136 3448
rect 13265 3417 13277 3420
rect 13219 3411 13277 3417
rect 7668 3352 7880 3380
rect 9263 3383 9321 3389
rect 9263 3349 9275 3383
rect 9309 3380 9321 3383
rect 9766 3380 9772 3392
rect 9309 3352 9772 3380
rect 9309 3349 9321 3352
rect 9263 3343 9321 3349
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 11011 3383 11069 3389
rect 11011 3349 11023 3383
rect 11057 3380 11069 3383
rect 11974 3380 11980 3392
rect 11057 3352 11980 3380
rect 11057 3349 11069 3352
rect 11011 3343 11069 3349
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 13354 3340 13360 3392
rect 13412 3380 13418 3392
rect 13817 3383 13875 3389
rect 13817 3380 13829 3383
rect 13412 3352 13829 3380
rect 13412 3340 13418 3352
rect 13817 3349 13829 3352
rect 13863 3349 13875 3383
rect 14108 3380 14136 3420
rect 14277 3417 14289 3451
rect 14323 3417 14335 3451
rect 14277 3411 14335 3417
rect 14292 3380 14320 3411
rect 14458 3408 14464 3460
rect 14516 3448 14522 3460
rect 16117 3451 16175 3457
rect 16117 3448 16129 3451
rect 14516 3420 16129 3448
rect 14516 3408 14522 3420
rect 16117 3417 16129 3420
rect 16163 3417 16175 3451
rect 16117 3411 16175 3417
rect 17037 3451 17095 3457
rect 17037 3417 17049 3451
rect 17083 3448 17095 3451
rect 17862 3448 17868 3460
rect 17083 3420 17868 3448
rect 17083 3417 17095 3420
rect 17037 3411 17095 3417
rect 17862 3408 17868 3420
rect 17920 3408 17926 3460
rect 14108 3352 14320 3380
rect 13817 3343 13875 3349
rect 1104 3290 18860 3312
rect 1104 3238 5398 3290
rect 5450 3238 5462 3290
rect 5514 3238 5526 3290
rect 5578 3238 5590 3290
rect 5642 3238 5654 3290
rect 5706 3238 9846 3290
rect 9898 3238 9910 3290
rect 9962 3238 9974 3290
rect 10026 3238 10038 3290
rect 10090 3238 10102 3290
rect 10154 3238 14294 3290
rect 14346 3238 14358 3290
rect 14410 3238 14422 3290
rect 14474 3238 14486 3290
rect 14538 3238 14550 3290
rect 14602 3238 18860 3290
rect 1104 3216 18860 3238
rect 3602 3136 3608 3188
rect 3660 3176 3666 3188
rect 8110 3176 8116 3188
rect 3660 3148 5948 3176
rect 3660 3136 3666 3148
rect 3694 3068 3700 3120
rect 3752 3108 3758 3120
rect 5537 3111 5595 3117
rect 5537 3108 5549 3111
rect 3752 3080 5549 3108
rect 3752 3068 3758 3080
rect 5537 3077 5549 3080
rect 5583 3077 5595 3111
rect 5537 3071 5595 3077
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 1762 3040 1768 3052
rect 1719 3012 1768 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2590 3040 2596 3052
rect 2547 3012 2596 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3040 3387 3043
rect 3418 3040 3424 3052
rect 3375 3012 3424 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 3418 3000 3424 3012
rect 3476 3000 3482 3052
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3040 4859 3043
rect 5074 3040 5080 3052
rect 4847 3012 5080 3040
rect 4847 3009 4859 3012
rect 4801 3003 4859 3009
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3009 5227 3043
rect 5169 3003 5227 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 934 2932 940 2984
rect 992 2972 998 2984
rect 1857 2975 1915 2981
rect 1857 2972 1869 2975
rect 992 2944 1869 2972
rect 992 2932 998 2944
rect 1857 2941 1869 2944
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 2314 2932 2320 2984
rect 2372 2972 2378 2984
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 2372 2944 2697 2972
rect 2372 2932 2378 2944
rect 2685 2941 2697 2944
rect 2731 2941 2743 2975
rect 4614 2972 4620 2984
rect 4575 2944 4620 2972
rect 2685 2935 2743 2941
rect 4614 2932 4620 2944
rect 4672 2932 4678 2984
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3145 2839 3203 2845
rect 3145 2836 3157 2839
rect 2832 2808 3157 2836
rect 2832 2796 2838 2808
rect 3145 2805 3157 2808
rect 3191 2805 3203 2839
rect 3145 2799 3203 2805
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 4985 2839 5043 2845
rect 4985 2836 4997 2839
rect 3568 2808 4997 2836
rect 3568 2796 3574 2808
rect 4985 2805 4997 2808
rect 5031 2805 5043 2839
rect 5184 2836 5212 3003
rect 5828 2904 5856 3003
rect 5920 2972 5948 3148
rect 6656 3148 8116 3176
rect 6656 3049 6684 3148
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 11790 3176 11796 3188
rect 8720 3148 11796 3176
rect 8720 3136 8726 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 11940 3148 13400 3176
rect 11940 3136 11946 3148
rect 7558 3068 7564 3120
rect 7616 3108 7622 3120
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 7616 3080 7849 3108
rect 7616 3068 7622 3080
rect 7837 3077 7849 3080
rect 7883 3077 7895 3111
rect 8754 3108 8760 3120
rect 8715 3080 8760 3108
rect 7837 3071 7895 3077
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 9306 3108 9312 3120
rect 9267 3080 9312 3108
rect 9306 3068 9312 3080
rect 9364 3068 9370 3120
rect 9766 3068 9772 3120
rect 9824 3108 9830 3120
rect 10229 3111 10287 3117
rect 10229 3108 10241 3111
rect 9824 3080 10241 3108
rect 9824 3068 9830 3080
rect 10229 3077 10241 3080
rect 10275 3077 10287 3111
rect 10229 3071 10287 3077
rect 11238 3068 11244 3120
rect 11296 3068 11302 3120
rect 11698 3108 11704 3120
rect 11659 3080 11704 3108
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 12066 3068 12072 3120
rect 12124 3108 12130 3120
rect 12124 3080 12572 3108
rect 12124 3068 12130 3080
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 7006 3000 7012 3052
rect 7064 3040 7070 3052
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 7064 3012 7205 3040
rect 7064 3000 7070 3012
rect 7193 3009 7205 3012
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3040 7343 3043
rect 7374 3040 7380 3052
rect 7331 3012 7380 3040
rect 7331 3009 7343 3012
rect 7285 3003 7343 3009
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 9214 3040 9220 3052
rect 9175 3012 9220 3040
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 10778 3040 10784 3052
rect 10739 3012 10784 3040
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11256 3040 11284 3068
rect 11195 3012 11284 3040
rect 12544 3040 12572 3080
rect 12618 3068 12624 3120
rect 12676 3108 12682 3120
rect 12943 3111 13001 3117
rect 12676 3080 12721 3108
rect 12676 3068 12682 3080
rect 12943 3077 12955 3111
rect 12989 3108 13001 3111
rect 13265 3111 13323 3117
rect 13265 3108 13277 3111
rect 12989 3080 13277 3108
rect 12989 3077 13001 3080
rect 12943 3071 13001 3077
rect 13265 3077 13277 3080
rect 13311 3077 13323 3111
rect 13372 3108 13400 3148
rect 13446 3136 13452 3188
rect 13504 3176 13510 3188
rect 13504 3148 17080 3176
rect 13504 3136 13510 3148
rect 14090 3108 14096 3120
rect 13372 3080 14096 3108
rect 13265 3071 13323 3077
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 14182 3068 14188 3120
rect 14240 3108 14246 3120
rect 14369 3111 14427 3117
rect 14369 3108 14381 3111
rect 14240 3080 14381 3108
rect 14240 3068 14246 3080
rect 14369 3077 14381 3080
rect 14415 3077 14427 3111
rect 14369 3071 14427 3077
rect 14461 3111 14519 3117
rect 14461 3077 14473 3111
rect 14507 3108 14519 3111
rect 14550 3108 14556 3120
rect 14507 3080 14556 3108
rect 14507 3077 14519 3080
rect 14461 3071 14519 3077
rect 14550 3068 14556 3080
rect 14608 3068 14614 3120
rect 14642 3068 14648 3120
rect 14700 3108 14706 3120
rect 14700 3080 16068 3108
rect 14700 3068 14706 3080
rect 12840 3043 12898 3049
rect 12840 3040 12852 3043
rect 12544 3012 12852 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 12840 3009 12852 3012
rect 12886 3009 12898 3043
rect 15470 3040 15476 3052
rect 15431 3012 15476 3040
rect 12840 3003 12898 3009
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 16040 3049 16068 3080
rect 16025 3043 16083 3049
rect 16025 3009 16037 3043
rect 16071 3009 16083 3043
rect 16025 3003 16083 3009
rect 16114 3000 16120 3052
rect 16172 3040 16178 3052
rect 17052 3049 17080 3148
rect 17126 3068 17132 3120
rect 17184 3108 17190 3120
rect 17184 3080 18276 3108
rect 17184 3068 17190 3080
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16172 3012 16681 3040
rect 16172 3000 16178 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3009 17095 3043
rect 17402 3040 17408 3052
rect 17363 3012 17408 3040
rect 17037 3003 17095 3009
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 17862 3040 17868 3052
rect 17823 3012 17868 3040
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 18248 3049 18276 3080
rect 18233 3043 18291 3049
rect 18233 3009 18245 3043
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 5920 2944 6929 2972
rect 6917 2941 6929 2944
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 7745 2975 7803 2981
rect 7745 2941 7757 2975
rect 7791 2960 7803 2975
rect 9398 2972 9404 2984
rect 7852 2960 9404 2972
rect 7791 2944 9404 2960
rect 7791 2941 7880 2944
rect 7745 2935 7880 2941
rect 7760 2932 7880 2935
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2972 10379 2975
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 10367 2944 11253 2972
rect 10367 2941 10379 2944
rect 10321 2935 10379 2941
rect 11241 2941 11253 2944
rect 11287 2972 11299 2975
rect 11287 2944 11560 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11532 2916 11560 2944
rect 11606 2932 11612 2984
rect 11664 2972 11670 2984
rect 11882 2972 11888 2984
rect 11664 2944 11888 2972
rect 11664 2932 11670 2944
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 13173 2975 13231 2981
rect 13173 2941 13185 2975
rect 13219 2941 13231 2975
rect 13998 2972 14004 2984
rect 13959 2944 14004 2972
rect 13173 2935 13231 2941
rect 5828 2876 7696 2904
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5184 2808 5917 2836
rect 4985 2799 5043 2805
rect 5905 2805 5917 2808
rect 5951 2836 5963 2839
rect 6362 2836 6368 2848
rect 5951 2808 6368 2836
rect 5951 2805 5963 2808
rect 5905 2799 5963 2805
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 6457 2839 6515 2845
rect 6457 2805 6469 2839
rect 6503 2836 6515 2839
rect 6914 2836 6920 2848
rect 6503 2808 6920 2836
rect 6503 2805 6515 2808
rect 6457 2799 6515 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7466 2836 7472 2848
rect 7427 2808 7472 2836
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 7668 2836 7696 2876
rect 10226 2864 10232 2916
rect 10284 2904 10290 2916
rect 10965 2907 11023 2913
rect 10965 2904 10977 2907
rect 10284 2876 10977 2904
rect 10284 2864 10290 2876
rect 10965 2873 10977 2876
rect 11011 2873 11023 2907
rect 10965 2867 11023 2873
rect 11514 2864 11520 2916
rect 11572 2864 11578 2916
rect 11790 2864 11796 2916
rect 11848 2904 11854 2916
rect 13078 2904 13084 2916
rect 11848 2876 13084 2904
rect 11848 2864 11854 2876
rect 13078 2864 13084 2876
rect 13136 2864 13142 2916
rect 8662 2836 8668 2848
rect 7668 2808 8668 2836
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 8754 2796 8760 2848
rect 8812 2836 8818 2848
rect 9033 2839 9091 2845
rect 9033 2836 9045 2839
rect 8812 2808 9045 2836
rect 8812 2796 8818 2808
rect 9033 2805 9045 2808
rect 9079 2805 9091 2839
rect 10594 2836 10600 2848
rect 10555 2808 10600 2836
rect 9033 2799 9091 2805
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 13188 2836 13216 2935
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 14645 2975 14703 2981
rect 14645 2972 14657 2975
rect 14235 2944 14657 2972
rect 13906 2864 13912 2916
rect 13964 2904 13970 2916
rect 14235 2904 14263 2944
rect 14645 2941 14657 2944
rect 14691 2941 14703 2975
rect 14645 2935 14703 2941
rect 13964 2876 14263 2904
rect 13964 2864 13970 2876
rect 14366 2864 14372 2916
rect 14424 2904 14430 2916
rect 15470 2904 15476 2916
rect 14424 2876 15476 2904
rect 14424 2864 14430 2876
rect 15470 2864 15476 2876
rect 15528 2864 15534 2916
rect 15841 2907 15899 2913
rect 15841 2904 15853 2907
rect 15580 2876 15853 2904
rect 13814 2836 13820 2848
rect 13188 2808 13820 2836
rect 13814 2796 13820 2808
rect 13872 2836 13878 2848
rect 15580 2836 15608 2876
rect 15841 2873 15853 2876
rect 15887 2873 15899 2907
rect 15841 2867 15899 2873
rect 18049 2907 18107 2913
rect 18049 2873 18061 2907
rect 18095 2904 18107 2907
rect 18874 2904 18880 2916
rect 18095 2876 18880 2904
rect 18095 2873 18107 2876
rect 18049 2867 18107 2873
rect 18874 2864 18880 2876
rect 18932 2864 18938 2916
rect 13872 2808 15608 2836
rect 15657 2839 15715 2845
rect 13872 2796 13878 2808
rect 15657 2805 15669 2839
rect 15703 2836 15715 2839
rect 15746 2836 15752 2848
rect 15703 2808 15752 2836
rect 15703 2805 15715 2808
rect 15657 2799 15715 2805
rect 15746 2796 15752 2808
rect 15804 2796 15810 2848
rect 16209 2839 16267 2845
rect 16209 2805 16221 2839
rect 16255 2836 16267 2839
rect 16390 2836 16396 2848
rect 16255 2808 16396 2836
rect 16255 2805 16267 2808
rect 16209 2799 16267 2805
rect 16390 2796 16396 2808
rect 16448 2796 16454 2848
rect 16853 2839 16911 2845
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 17034 2836 17040 2848
rect 16899 2808 17040 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 17221 2839 17279 2845
rect 17221 2805 17233 2839
rect 17267 2836 17279 2839
rect 17494 2836 17500 2848
rect 17267 2808 17500 2836
rect 17267 2805 17279 2808
rect 17221 2799 17279 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 17589 2839 17647 2845
rect 17589 2805 17601 2839
rect 17635 2836 17647 2839
rect 17954 2836 17960 2848
rect 17635 2808 17960 2836
rect 17635 2805 17647 2808
rect 17589 2799 17647 2805
rect 17954 2796 17960 2808
rect 18012 2796 18018 2848
rect 18414 2836 18420 2848
rect 18375 2808 18420 2836
rect 18414 2796 18420 2808
rect 18472 2796 18478 2848
rect 1104 2746 18860 2768
rect 1104 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 3430 2746
rect 3482 2694 7622 2746
rect 7674 2694 7686 2746
rect 7738 2694 7750 2746
rect 7802 2694 7814 2746
rect 7866 2694 7878 2746
rect 7930 2694 12070 2746
rect 12122 2694 12134 2746
rect 12186 2694 12198 2746
rect 12250 2694 12262 2746
rect 12314 2694 12326 2746
rect 12378 2694 16518 2746
rect 16570 2694 16582 2746
rect 16634 2694 16646 2746
rect 16698 2694 16710 2746
rect 16762 2694 16774 2746
rect 16826 2694 18860 2746
rect 1104 2672 18860 2694
rect 11195 2635 11253 2641
rect 11195 2601 11207 2635
rect 11241 2632 11253 2635
rect 11698 2632 11704 2644
rect 11241 2604 11704 2632
rect 11241 2601 11253 2604
rect 11195 2595 11253 2601
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 14323 2635 14381 2641
rect 14323 2601 14335 2635
rect 14369 2632 14381 2635
rect 14458 2632 14464 2644
rect 14369 2604 14464 2632
rect 14369 2601 14381 2604
rect 14323 2595 14381 2601
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 15470 2632 15476 2644
rect 15431 2604 15476 2632
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 17681 2635 17739 2641
rect 17681 2632 17693 2635
rect 16546 2604 17693 2632
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 10505 2567 10563 2573
rect 10505 2564 10517 2567
rect 9732 2536 10517 2564
rect 9732 2524 9738 2536
rect 10505 2533 10517 2536
rect 10551 2533 10563 2567
rect 10870 2564 10876 2576
rect 10505 2527 10563 2533
rect 10612 2536 10876 2564
rect 10612 2496 10640 2536
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 11054 2524 11060 2576
rect 11112 2564 11118 2576
rect 14645 2567 14703 2573
rect 11112 2536 14596 2564
rect 11112 2524 11118 2536
rect 11698 2496 11704 2508
rect 7024 2468 10640 2496
rect 10704 2468 11704 2496
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 4890 2428 4896 2440
rect 2179 2400 4896 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 7024 2437 7052 2468
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 9122 2428 9128 2440
rect 7883 2400 9128 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 9490 2428 9496 2440
rect 9263 2400 9496 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 9766 2388 9772 2440
rect 9824 2428 9830 2440
rect 10704 2437 10732 2468
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 12894 2496 12900 2508
rect 12855 2468 12900 2496
rect 12894 2456 12900 2468
rect 12952 2456 12958 2508
rect 12986 2456 12992 2508
rect 13044 2496 13050 2508
rect 14568 2496 14596 2536
rect 14645 2533 14657 2567
rect 14691 2564 14703 2567
rect 15194 2564 15200 2576
rect 14691 2536 15200 2564
rect 14691 2533 14703 2536
rect 14645 2527 14703 2533
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 16546 2496 16574 2604
rect 17681 2601 17693 2604
rect 17727 2601 17739 2635
rect 17681 2595 17739 2601
rect 13044 2468 14504 2496
rect 14568 2468 16574 2496
rect 13044 2456 13050 2468
rect 11146 2437 11152 2440
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 9824 2400 10241 2428
rect 9824 2388 9830 2400
rect 10229 2397 10241 2400
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2397 10747 2431
rect 10689 2391 10747 2397
rect 11124 2431 11152 2437
rect 11124 2397 11136 2431
rect 11124 2391 11152 2397
rect 11146 2388 11152 2391
rect 11204 2388 11210 2440
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14476 2437 14504 2468
rect 14220 2431 14278 2437
rect 14220 2428 14232 2431
rect 14148 2400 14232 2428
rect 14148 2388 14154 2400
rect 14220 2397 14232 2400
rect 14266 2397 14278 2431
rect 14220 2391 14278 2397
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2397 14519 2431
rect 14826 2428 14832 2440
rect 14787 2400 14832 2428
rect 14461 2391 14519 2397
rect 14826 2388 14832 2400
rect 14884 2388 14890 2440
rect 17696 2428 17724 2595
rect 17865 2431 17923 2437
rect 17865 2428 17877 2431
rect 17696 2400 17877 2428
rect 17865 2397 17877 2400
rect 17911 2397 17923 2431
rect 17865 2391 17923 2397
rect 1394 2320 1400 2372
rect 1452 2360 1458 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 1452 2332 1869 2360
rect 1452 2320 1458 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 4212 2332 6745 2360
rect 4212 2320 4218 2332
rect 6733 2329 6745 2332
rect 6779 2329 6791 2363
rect 9398 2360 9404 2372
rect 9311 2332 9404 2360
rect 6733 2323 6791 2329
rect 9398 2320 9404 2332
rect 9456 2360 9462 2372
rect 11885 2363 11943 2369
rect 9456 2332 11100 2360
rect 9456 2320 9462 2332
rect 11072 2304 11100 2332
rect 11885 2329 11897 2363
rect 11931 2329 11943 2363
rect 11885 2323 11943 2329
rect 7374 2252 7380 2304
rect 7432 2292 7438 2304
rect 7653 2295 7711 2301
rect 7653 2292 7665 2295
rect 7432 2264 7665 2292
rect 7432 2252 7438 2264
rect 7653 2261 7665 2264
rect 7699 2261 7711 2295
rect 7653 2255 7711 2261
rect 8294 2252 8300 2304
rect 8352 2292 8358 2304
rect 9033 2295 9091 2301
rect 9033 2292 9045 2295
rect 8352 2264 9045 2292
rect 8352 2252 8358 2264
rect 9033 2261 9045 2264
rect 9079 2261 9091 2295
rect 9033 2255 9091 2261
rect 9490 2252 9496 2304
rect 9548 2292 9554 2304
rect 10045 2295 10103 2301
rect 10045 2292 10057 2295
rect 9548 2264 10057 2292
rect 9548 2252 9554 2264
rect 10045 2261 10057 2264
rect 10091 2261 10103 2295
rect 10045 2255 10103 2261
rect 11054 2252 11060 2304
rect 11112 2252 11118 2304
rect 11900 2292 11928 2323
rect 11974 2320 11980 2372
rect 12032 2360 12038 2372
rect 16114 2360 16120 2372
rect 12032 2332 12077 2360
rect 15028 2332 16120 2360
rect 12032 2320 12038 2332
rect 12434 2292 12440 2304
rect 11900 2264 12440 2292
rect 12434 2252 12440 2264
rect 12492 2292 12498 2304
rect 15028 2301 15056 2332
rect 16114 2320 16120 2332
rect 16172 2320 16178 2372
rect 12989 2295 13047 2301
rect 12989 2292 13001 2295
rect 12492 2264 13001 2292
rect 12492 2252 12498 2264
rect 12989 2261 13001 2264
rect 13035 2261 13047 2295
rect 12989 2255 13047 2261
rect 15013 2295 15071 2301
rect 15013 2261 15025 2295
rect 15059 2261 15071 2295
rect 18046 2292 18052 2304
rect 18007 2264 18052 2292
rect 15013 2255 15071 2261
rect 18046 2252 18052 2264
rect 18104 2252 18110 2304
rect 1104 2202 18860 2224
rect 1104 2150 5398 2202
rect 5450 2150 5462 2202
rect 5514 2150 5526 2202
rect 5578 2150 5590 2202
rect 5642 2150 5654 2202
rect 5706 2150 9846 2202
rect 9898 2150 9910 2202
rect 9962 2150 9974 2202
rect 10026 2150 10038 2202
rect 10090 2150 10102 2202
rect 10154 2150 14294 2202
rect 14346 2150 14358 2202
rect 14410 2150 14422 2202
rect 14474 2150 14486 2202
rect 14538 2150 14550 2202
rect 14602 2150 18860 2202
rect 1104 2128 18860 2150
rect 2774 1708 2780 1760
rect 2832 1748 2838 1760
rect 3050 1748 3056 1760
rect 2832 1720 3056 1748
rect 2832 1708 2838 1720
rect 3050 1708 3056 1720
rect 3108 1708 3114 1760
<< via1 >>
rect 11704 15172 11756 15224
rect 15476 15172 15528 15224
rect 4436 14900 4488 14952
rect 11244 14900 11296 14952
rect 8852 14832 8904 14884
rect 17040 14832 17092 14884
rect 3516 14764 3568 14816
rect 13360 14764 13412 14816
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 3302 14662 3354 14714
rect 3366 14662 3418 14714
rect 3430 14662 3482 14714
rect 7622 14662 7674 14714
rect 7686 14662 7738 14714
rect 7750 14662 7802 14714
rect 7814 14662 7866 14714
rect 7878 14662 7930 14714
rect 12070 14662 12122 14714
rect 12134 14662 12186 14714
rect 12198 14662 12250 14714
rect 12262 14662 12314 14714
rect 12326 14662 12378 14714
rect 16518 14662 16570 14714
rect 16582 14662 16634 14714
rect 16646 14662 16698 14714
rect 16710 14662 16762 14714
rect 16774 14662 16826 14714
rect 2964 14560 3016 14612
rect 13636 14560 13688 14612
rect 2228 14424 2280 14476
rect 11152 14492 11204 14544
rect 11244 14492 11296 14544
rect 15844 14492 15896 14544
rect 7748 14424 7800 14476
rect 17316 14424 17368 14476
rect 1216 14356 1268 14408
rect 8576 14356 8628 14408
rect 9128 14356 9180 14408
rect 16396 14356 16448 14408
rect 2872 14288 2924 14340
rect 9772 14288 9824 14340
rect 12440 14288 12492 14340
rect 12992 14288 13044 14340
rect 18328 14288 18380 14340
rect 4804 14220 4856 14272
rect 13728 14220 13780 14272
rect 5398 14118 5450 14170
rect 5462 14118 5514 14170
rect 5526 14118 5578 14170
rect 5590 14118 5642 14170
rect 5654 14118 5706 14170
rect 9846 14118 9898 14170
rect 9910 14118 9962 14170
rect 9974 14118 10026 14170
rect 10038 14118 10090 14170
rect 10102 14118 10154 14170
rect 14294 14118 14346 14170
rect 14358 14118 14410 14170
rect 14422 14118 14474 14170
rect 14486 14118 14538 14170
rect 14550 14118 14602 14170
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 6736 14016 6788 14068
rect 7748 14059 7800 14068
rect 7748 14025 7757 14059
rect 7757 14025 7791 14059
rect 7791 14025 7800 14059
rect 7748 14016 7800 14025
rect 8576 14059 8628 14068
rect 5540 13948 5592 14000
rect 8576 14025 8585 14059
rect 8585 14025 8619 14059
rect 8619 14025 8628 14059
rect 8576 14016 8628 14025
rect 8852 14059 8904 14068
rect 8852 14025 8861 14059
rect 8861 14025 8895 14059
rect 8895 14025 8904 14059
rect 8852 14016 8904 14025
rect 9128 14059 9180 14068
rect 9128 14025 9137 14059
rect 9137 14025 9171 14059
rect 9171 14025 9180 14059
rect 9128 14016 9180 14025
rect 9772 14016 9824 14068
rect 11152 14059 11204 14068
rect 11152 14025 11161 14059
rect 11161 14025 11195 14059
rect 11195 14025 11204 14059
rect 11152 14016 11204 14025
rect 12624 14059 12676 14068
rect 12624 14025 12633 14059
rect 12633 14025 12667 14059
rect 12667 14025 12676 14059
rect 12624 14016 12676 14025
rect 13360 14059 13412 14068
rect 13360 14025 13369 14059
rect 13369 14025 13403 14059
rect 13403 14025 13412 14059
rect 13360 14016 13412 14025
rect 13728 14059 13780 14068
rect 13728 14025 13737 14059
rect 13737 14025 13771 14059
rect 13771 14025 13780 14059
rect 13728 14016 13780 14025
rect 14096 14059 14148 14068
rect 14096 14025 14105 14059
rect 14105 14025 14139 14059
rect 14139 14025 14148 14059
rect 14096 14016 14148 14025
rect 14924 14016 14976 14068
rect 19616 14016 19668 14068
rect 6000 13812 6052 13864
rect 6460 13880 6512 13932
rect 7748 13880 7800 13932
rect 8852 13880 8904 13932
rect 12440 13948 12492 14000
rect 14004 13948 14056 14000
rect 13912 13923 13964 13932
rect 13176 13812 13228 13864
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 15108 13880 15160 13932
rect 15476 13880 15528 13932
rect 15752 13880 15804 13932
rect 14096 13812 14148 13864
rect 1584 13744 1636 13796
rect 296 13676 348 13728
rect 5540 13676 5592 13728
rect 6368 13676 6420 13728
rect 11612 13719 11664 13728
rect 11612 13685 11621 13719
rect 11621 13685 11655 13719
rect 11655 13685 11664 13719
rect 11612 13676 11664 13685
rect 15016 13719 15068 13728
rect 15016 13685 15025 13719
rect 15025 13685 15059 13719
rect 15059 13685 15068 13719
rect 15016 13676 15068 13685
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 3302 13574 3354 13626
rect 3366 13574 3418 13626
rect 3430 13574 3482 13626
rect 7622 13574 7674 13626
rect 7686 13574 7738 13626
rect 7750 13574 7802 13626
rect 7814 13574 7866 13626
rect 7878 13574 7930 13626
rect 12070 13574 12122 13626
rect 12134 13574 12186 13626
rect 12198 13574 12250 13626
rect 12262 13574 12314 13626
rect 12326 13574 12378 13626
rect 16518 13574 16570 13626
rect 16582 13574 16634 13626
rect 16646 13574 16698 13626
rect 16710 13574 16762 13626
rect 16774 13574 16826 13626
rect 11612 13472 11664 13524
rect 12164 13472 12216 13524
rect 5908 13336 5960 13388
rect 6828 13404 6880 13456
rect 8208 13336 8260 13388
rect 9404 13336 9456 13388
rect 11980 13336 12032 13388
rect 12440 13379 12492 13388
rect 12440 13345 12449 13379
rect 12449 13345 12483 13379
rect 12483 13345 12492 13379
rect 12440 13336 12492 13345
rect 2872 13268 2924 13320
rect 12072 13268 12124 13320
rect 12164 13311 12216 13320
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 13268 13336 13320 13388
rect 15292 13336 15344 13388
rect 12164 13268 12216 13277
rect 15200 13268 15252 13320
rect 3976 13200 4028 13252
rect 5264 13200 5316 13252
rect 5172 13175 5224 13184
rect 5172 13141 5181 13175
rect 5181 13141 5215 13175
rect 5215 13141 5224 13175
rect 5172 13132 5224 13141
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 7012 13200 7064 13252
rect 16028 13200 16080 13252
rect 7196 13175 7248 13184
rect 7196 13141 7205 13175
rect 7205 13141 7239 13175
rect 7239 13141 7248 13175
rect 7196 13132 7248 13141
rect 8300 13132 8352 13184
rect 9588 13175 9640 13184
rect 9588 13141 9597 13175
rect 9597 13141 9631 13175
rect 9631 13141 9640 13175
rect 9588 13132 9640 13141
rect 11152 13132 11204 13184
rect 11336 13175 11388 13184
rect 11336 13141 11345 13175
rect 11345 13141 11379 13175
rect 11379 13141 11388 13175
rect 11336 13132 11388 13141
rect 12624 13175 12676 13184
rect 12624 13141 12633 13175
rect 12633 13141 12667 13175
rect 12667 13141 12676 13175
rect 12624 13132 12676 13141
rect 13820 13175 13872 13184
rect 13820 13141 13829 13175
rect 13829 13141 13863 13175
rect 13863 13141 13872 13175
rect 13820 13132 13872 13141
rect 5398 13030 5450 13082
rect 5462 13030 5514 13082
rect 5526 13030 5578 13082
rect 5590 13030 5642 13082
rect 5654 13030 5706 13082
rect 9846 13030 9898 13082
rect 9910 13030 9962 13082
rect 9974 13030 10026 13082
rect 10038 13030 10090 13082
rect 10102 13030 10154 13082
rect 14294 13030 14346 13082
rect 14358 13030 14410 13082
rect 14422 13030 14474 13082
rect 14486 13030 14538 13082
rect 14550 13030 14602 13082
rect 2872 12928 2924 12980
rect 3056 12928 3108 12980
rect 3884 12971 3936 12980
rect 3884 12937 3893 12971
rect 3893 12937 3927 12971
rect 3927 12937 3936 12971
rect 3884 12928 3936 12937
rect 4436 12971 4488 12980
rect 2964 12860 3016 12912
rect 4436 12937 4445 12971
rect 4445 12937 4479 12971
rect 4479 12937 4488 12971
rect 4436 12928 4488 12937
rect 5172 12971 5224 12980
rect 5172 12937 5181 12971
rect 5181 12937 5215 12971
rect 5215 12937 5224 12971
rect 5172 12928 5224 12937
rect 5264 12928 5316 12980
rect 6368 12928 6420 12980
rect 7196 12928 7248 12980
rect 10232 12928 10284 12980
rect 11152 12928 11204 12980
rect 11336 12928 11388 12980
rect 12624 12928 12676 12980
rect 4068 12860 4120 12912
rect 6276 12860 6328 12912
rect 12072 12903 12124 12912
rect 6644 12792 6696 12844
rect 7196 12792 7248 12844
rect 9680 12792 9732 12844
rect 12072 12869 12081 12903
rect 12081 12869 12115 12903
rect 12115 12869 12124 12903
rect 12072 12860 12124 12869
rect 13268 12860 13320 12912
rect 13820 12860 13872 12912
rect 15660 12860 15712 12912
rect 2872 12656 2924 12708
rect 4068 12767 4120 12776
rect 4068 12733 4077 12767
rect 4077 12733 4111 12767
rect 4111 12733 4120 12767
rect 4068 12724 4120 12733
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 6368 12724 6420 12776
rect 6828 12724 6880 12776
rect 8208 12724 8260 12776
rect 9496 12724 9548 12776
rect 10232 12767 10284 12776
rect 10232 12733 10241 12767
rect 10241 12733 10275 12767
rect 10275 12733 10284 12767
rect 10232 12724 10284 12733
rect 14096 12792 14148 12844
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 12440 12724 12492 12776
rect 13360 12724 13412 12776
rect 14464 12767 14516 12776
rect 14464 12733 14473 12767
rect 14473 12733 14507 12767
rect 14507 12733 14516 12767
rect 14464 12724 14516 12733
rect 7012 12656 7064 12708
rect 7104 12656 7156 12708
rect 10508 12699 10560 12708
rect 10508 12665 10517 12699
rect 10517 12665 10551 12699
rect 10551 12665 10560 12699
rect 10508 12656 10560 12665
rect 12164 12656 12216 12708
rect 17868 12656 17920 12708
rect 2044 12588 2096 12640
rect 3516 12631 3568 12640
rect 3516 12597 3525 12631
rect 3525 12597 3559 12631
rect 3559 12597 3568 12631
rect 3516 12588 3568 12597
rect 4804 12631 4856 12640
rect 4804 12597 4813 12631
rect 4813 12597 4847 12631
rect 4847 12597 4856 12631
rect 4804 12588 4856 12597
rect 11796 12588 11848 12640
rect 12624 12631 12676 12640
rect 12624 12597 12633 12631
rect 12633 12597 12667 12631
rect 12667 12597 12676 12631
rect 12624 12588 12676 12597
rect 13084 12631 13136 12640
rect 13084 12597 13093 12631
rect 13093 12597 13127 12631
rect 13127 12597 13136 12631
rect 13084 12588 13136 12597
rect 14280 12588 14332 12640
rect 16396 12588 16448 12640
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 3302 12486 3354 12538
rect 3366 12486 3418 12538
rect 3430 12486 3482 12538
rect 7622 12486 7674 12538
rect 7686 12486 7738 12538
rect 7750 12486 7802 12538
rect 7814 12486 7866 12538
rect 7878 12486 7930 12538
rect 12070 12486 12122 12538
rect 12134 12486 12186 12538
rect 12198 12486 12250 12538
rect 12262 12486 12314 12538
rect 12326 12486 12378 12538
rect 16518 12486 16570 12538
rect 16582 12486 16634 12538
rect 16646 12486 16698 12538
rect 16710 12486 16762 12538
rect 16774 12486 16826 12538
rect 2964 12384 3016 12436
rect 7288 12384 7340 12436
rect 9496 12384 9548 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 11704 12384 11756 12436
rect 12440 12384 12492 12436
rect 14096 12427 14148 12436
rect 2688 12316 2740 12368
rect 3148 12316 3200 12368
rect 12716 12316 12768 12368
rect 13636 12316 13688 12368
rect 4068 12248 4120 12300
rect 6552 12248 6604 12300
rect 7380 12248 7432 12300
rect 9588 12291 9640 12300
rect 9588 12257 9597 12291
rect 9597 12257 9631 12291
rect 9631 12257 9640 12291
rect 9588 12248 9640 12257
rect 10232 12291 10284 12300
rect 10232 12257 10241 12291
rect 10241 12257 10275 12291
rect 10275 12257 10284 12291
rect 10232 12248 10284 12257
rect 11612 12248 11664 12300
rect 11704 12248 11756 12300
rect 11980 12248 12032 12300
rect 12624 12248 12676 12300
rect 13360 12291 13412 12300
rect 3700 12180 3752 12232
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 7564 12180 7616 12232
rect 10416 12180 10468 12232
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 13084 12180 13136 12232
rect 13360 12257 13369 12291
rect 13369 12257 13403 12291
rect 13403 12257 13412 12291
rect 13360 12248 13412 12257
rect 13544 12180 13596 12232
rect 14096 12393 14105 12427
rect 14105 12393 14139 12427
rect 14139 12393 14148 12427
rect 14096 12384 14148 12393
rect 14648 12291 14700 12300
rect 14648 12257 14657 12291
rect 14657 12257 14691 12291
rect 14691 12257 14700 12291
rect 14648 12248 14700 12257
rect 15200 12291 15252 12300
rect 15200 12257 15209 12291
rect 15209 12257 15243 12291
rect 15243 12257 15252 12291
rect 15200 12248 15252 12257
rect 15844 12248 15896 12300
rect 16120 12248 16172 12300
rect 16764 12180 16816 12232
rect 3148 12155 3200 12164
rect 3148 12121 3157 12155
rect 3157 12121 3191 12155
rect 3191 12121 3200 12155
rect 3148 12112 3200 12121
rect 4160 12112 4212 12164
rect 5172 12112 5224 12164
rect 3332 12044 3384 12096
rect 4344 12044 4396 12096
rect 4896 12087 4948 12096
rect 4896 12053 4905 12087
rect 4905 12053 4939 12087
rect 4939 12053 4948 12087
rect 6092 12087 6144 12096
rect 4896 12044 4948 12053
rect 6092 12053 6101 12087
rect 6101 12053 6135 12087
rect 6135 12053 6144 12087
rect 6092 12044 6144 12053
rect 7196 12044 7248 12096
rect 9404 12112 9456 12164
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 10508 12087 10560 12096
rect 10508 12053 10517 12087
rect 10517 12053 10551 12087
rect 10551 12053 10560 12087
rect 10508 12044 10560 12053
rect 10876 12087 10928 12096
rect 10876 12053 10885 12087
rect 10885 12053 10919 12087
rect 10919 12053 10928 12087
rect 10876 12044 10928 12053
rect 12716 12044 12768 12096
rect 12900 12112 12952 12164
rect 13268 12087 13320 12096
rect 13268 12053 13277 12087
rect 13277 12053 13311 12087
rect 13311 12053 13320 12087
rect 13268 12044 13320 12053
rect 14096 12044 14148 12096
rect 15844 12044 15896 12096
rect 18604 12044 18656 12096
rect 5398 11942 5450 11994
rect 5462 11942 5514 11994
rect 5526 11942 5578 11994
rect 5590 11942 5642 11994
rect 5654 11942 5706 11994
rect 9846 11942 9898 11994
rect 9910 11942 9962 11994
rect 9974 11942 10026 11994
rect 10038 11942 10090 11994
rect 10102 11942 10154 11994
rect 14294 11942 14346 11994
rect 14358 11942 14410 11994
rect 14422 11942 14474 11994
rect 14486 11942 14538 11994
rect 14550 11942 14602 11994
rect 2688 11883 2740 11892
rect 2688 11849 2697 11883
rect 2697 11849 2731 11883
rect 2731 11849 2740 11883
rect 2688 11840 2740 11849
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 3332 11883 3384 11892
rect 3332 11849 3341 11883
rect 3341 11849 3375 11883
rect 3375 11849 3384 11883
rect 3332 11840 3384 11849
rect 3516 11840 3568 11892
rect 4344 11883 4396 11892
rect 4344 11849 4353 11883
rect 4353 11849 4387 11883
rect 4387 11849 4396 11883
rect 4344 11840 4396 11849
rect 4896 11840 4948 11892
rect 6460 11840 6512 11892
rect 6644 11883 6696 11892
rect 6644 11849 6653 11883
rect 6653 11849 6687 11883
rect 6687 11849 6696 11883
rect 6644 11840 6696 11849
rect 7104 11883 7156 11892
rect 7104 11849 7113 11883
rect 7113 11849 7147 11883
rect 7147 11849 7156 11883
rect 7104 11840 7156 11849
rect 8300 11883 8352 11892
rect 8300 11849 8309 11883
rect 8309 11849 8343 11883
rect 8343 11849 8352 11883
rect 8300 11840 8352 11849
rect 6092 11772 6144 11824
rect 10416 11840 10468 11892
rect 12440 11840 12492 11892
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 2872 11704 2924 11756
rect 3792 11704 3844 11756
rect 4068 11704 4120 11756
rect 12900 11840 12952 11892
rect 13268 11840 13320 11892
rect 15200 11840 15252 11892
rect 16764 11883 16816 11892
rect 16764 11849 16773 11883
rect 16773 11849 16807 11883
rect 16807 11849 16816 11883
rect 16764 11840 16816 11849
rect 17408 11840 17460 11892
rect 13544 11772 13596 11824
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 6920 11704 6972 11756
rect 8576 11704 8628 11756
rect 10416 11747 10468 11756
rect 10416 11713 10425 11747
rect 10425 11713 10459 11747
rect 10459 11713 10468 11747
rect 10416 11704 10468 11713
rect 12808 11704 12860 11756
rect 14188 11704 14240 11756
rect 2780 11568 2832 11620
rect 2872 11568 2924 11620
rect 6276 11636 6328 11688
rect 7288 11636 7340 11688
rect 7380 11568 7432 11620
rect 8392 11568 8444 11620
rect 8668 11636 8720 11688
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 10048 11679 10100 11688
rect 10048 11645 10057 11679
rect 10057 11645 10091 11679
rect 10091 11645 10100 11679
rect 10048 11636 10100 11645
rect 10232 11679 10284 11688
rect 10232 11645 10241 11679
rect 10241 11645 10275 11679
rect 10275 11645 10284 11679
rect 10232 11636 10284 11645
rect 12624 11636 12676 11688
rect 14648 11636 14700 11688
rect 15108 11747 15160 11756
rect 15108 11713 15117 11747
rect 15117 11713 15151 11747
rect 15151 11713 15160 11747
rect 15108 11704 15160 11713
rect 15752 11704 15804 11756
rect 16028 11679 16080 11688
rect 9772 11568 9824 11620
rect 10508 11568 10560 11620
rect 14096 11568 14148 11620
rect 14832 11568 14884 11620
rect 16028 11645 16037 11679
rect 16037 11645 16071 11679
rect 16071 11645 16080 11679
rect 16028 11636 16080 11645
rect 3056 11500 3108 11552
rect 5908 11500 5960 11552
rect 6276 11500 6328 11552
rect 6460 11543 6512 11552
rect 6460 11509 6469 11543
rect 6469 11509 6503 11543
rect 6503 11509 6512 11543
rect 6460 11500 6512 11509
rect 6920 11500 6972 11552
rect 7564 11543 7616 11552
rect 7564 11509 7573 11543
rect 7573 11509 7607 11543
rect 7607 11509 7616 11543
rect 7564 11500 7616 11509
rect 9312 11500 9364 11552
rect 9496 11500 9548 11552
rect 9680 11500 9732 11552
rect 11796 11500 11848 11552
rect 13820 11500 13872 11552
rect 15108 11500 15160 11552
rect 15384 11500 15436 11552
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 16028 11500 16080 11552
rect 16212 11500 16264 11552
rect 18236 11500 18288 11552
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 3302 11398 3354 11450
rect 3366 11398 3418 11450
rect 3430 11398 3482 11450
rect 7622 11398 7674 11450
rect 7686 11398 7738 11450
rect 7750 11398 7802 11450
rect 7814 11398 7866 11450
rect 7878 11398 7930 11450
rect 12070 11398 12122 11450
rect 12134 11398 12186 11450
rect 12198 11398 12250 11450
rect 12262 11398 12314 11450
rect 12326 11398 12378 11450
rect 16518 11398 16570 11450
rect 16582 11398 16634 11450
rect 16646 11398 16698 11450
rect 16710 11398 16762 11450
rect 16774 11398 16826 11450
rect 2504 11296 2556 11348
rect 6368 11296 6420 11348
rect 6828 11296 6880 11348
rect 3056 11203 3108 11212
rect 3056 11169 3065 11203
rect 3065 11169 3099 11203
rect 3099 11169 3108 11203
rect 3056 11160 3108 11169
rect 7012 11228 7064 11280
rect 9404 11296 9456 11348
rect 9588 11296 9640 11348
rect 9772 11339 9824 11348
rect 9772 11305 9781 11339
rect 9781 11305 9815 11339
rect 9815 11305 9824 11339
rect 9772 11296 9824 11305
rect 4712 11160 4764 11212
rect 6368 11160 6420 11212
rect 7288 11160 7340 11212
rect 9496 11228 9548 11280
rect 12716 11228 12768 11280
rect 13084 11271 13136 11280
rect 13084 11237 13093 11271
rect 13093 11237 13127 11271
rect 13127 11237 13136 11271
rect 15752 11296 15804 11348
rect 15844 11296 15896 11348
rect 13084 11228 13136 11237
rect 8300 11203 8352 11212
rect 8300 11169 8309 11203
rect 8309 11169 8343 11203
rect 8343 11169 8352 11203
rect 8576 11203 8628 11212
rect 8300 11160 8352 11169
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 9588 11203 9640 11212
rect 9588 11169 9597 11203
rect 9597 11169 9631 11203
rect 9631 11169 9640 11203
rect 9588 11160 9640 11169
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 15384 11203 15436 11212
rect 15384 11169 15393 11203
rect 15393 11169 15427 11203
rect 15427 11169 15436 11203
rect 15384 11160 15436 11169
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 4528 11092 4580 11144
rect 5816 11092 5868 11144
rect 6184 11092 6236 11144
rect 9312 11135 9364 11144
rect 6276 11024 6328 11076
rect 8668 11024 8720 11076
rect 9312 11101 9321 11135
rect 9321 11101 9355 11135
rect 9355 11101 9364 11135
rect 9312 11092 9364 11101
rect 9588 11024 9640 11076
rect 2596 10999 2648 11008
rect 2596 10965 2605 10999
rect 2605 10965 2639 10999
rect 2639 10965 2648 10999
rect 2596 10956 2648 10965
rect 4068 10956 4120 11008
rect 10048 11024 10100 11076
rect 10968 11024 11020 11076
rect 11520 11092 11572 11144
rect 11336 11024 11388 11076
rect 14648 11024 14700 11076
rect 15568 11092 15620 11144
rect 15752 11160 15804 11212
rect 15844 11092 15896 11144
rect 17408 11203 17460 11212
rect 17408 11169 17417 11203
rect 17417 11169 17451 11203
rect 17451 11169 17460 11203
rect 17408 11160 17460 11169
rect 17224 11024 17276 11076
rect 18144 11228 18196 11280
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 18512 11067 18564 11076
rect 14924 10999 14976 11008
rect 14924 10965 14933 10999
rect 14933 10965 14967 10999
rect 14967 10965 14976 10999
rect 14924 10956 14976 10965
rect 16856 10956 16908 11008
rect 18512 11033 18521 11067
rect 18521 11033 18555 11067
rect 18555 11033 18564 11067
rect 18512 11024 18564 11033
rect 5398 10854 5450 10906
rect 5462 10854 5514 10906
rect 5526 10854 5578 10906
rect 5590 10854 5642 10906
rect 5654 10854 5706 10906
rect 9846 10854 9898 10906
rect 9910 10854 9962 10906
rect 9974 10854 10026 10906
rect 10038 10854 10090 10906
rect 10102 10854 10154 10906
rect 14294 10854 14346 10906
rect 14358 10854 14410 10906
rect 14422 10854 14474 10906
rect 14486 10854 14538 10906
rect 14550 10854 14602 10906
rect 2688 10752 2740 10804
rect 4068 10752 4120 10804
rect 6920 10752 6972 10804
rect 1952 10684 2004 10736
rect 4160 10684 4212 10736
rect 5908 10727 5960 10736
rect 5908 10693 5926 10727
rect 5926 10693 5960 10727
rect 5908 10684 5960 10693
rect 6828 10684 6880 10736
rect 3056 10616 3108 10668
rect 9404 10752 9456 10804
rect 8392 10684 8444 10736
rect 11704 10752 11756 10804
rect 14648 10795 14700 10804
rect 14648 10761 14657 10795
rect 14657 10761 14691 10795
rect 14691 10761 14700 10795
rect 14648 10752 14700 10761
rect 13360 10684 13412 10736
rect 16488 10684 16540 10736
rect 17500 10727 17552 10736
rect 17500 10693 17509 10727
rect 17509 10693 17543 10727
rect 17543 10693 17552 10727
rect 17500 10684 17552 10693
rect 8208 10616 8260 10668
rect 11704 10616 11756 10668
rect 12624 10659 12676 10668
rect 12624 10625 12642 10659
rect 12642 10625 12676 10659
rect 12624 10616 12676 10625
rect 2228 10548 2280 10600
rect 2872 10591 2924 10600
rect 2872 10557 2881 10591
rect 2881 10557 2915 10591
rect 2915 10557 2924 10591
rect 2872 10548 2924 10557
rect 4988 10548 5040 10600
rect 9680 10591 9732 10600
rect 2504 10412 2556 10464
rect 2688 10412 2740 10464
rect 4160 10455 4212 10464
rect 4160 10421 4169 10455
rect 4169 10421 4203 10455
rect 4203 10421 4212 10455
rect 4160 10412 4212 10421
rect 4896 10412 4948 10464
rect 5264 10412 5316 10464
rect 5816 10412 5868 10464
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 16948 10616 17000 10668
rect 14464 10548 14516 10557
rect 15752 10548 15804 10600
rect 6828 10412 6880 10464
rect 10968 10480 11020 10532
rect 11612 10412 11664 10464
rect 17224 10591 17276 10600
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 15752 10412 15804 10464
rect 15936 10412 15988 10464
rect 18328 10412 18380 10464
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 3430 10310 3482 10362
rect 7622 10310 7674 10362
rect 7686 10310 7738 10362
rect 7750 10310 7802 10362
rect 7814 10310 7866 10362
rect 7878 10310 7930 10362
rect 12070 10310 12122 10362
rect 12134 10310 12186 10362
rect 12198 10310 12250 10362
rect 12262 10310 12314 10362
rect 12326 10310 12378 10362
rect 16518 10310 16570 10362
rect 16582 10310 16634 10362
rect 16646 10310 16698 10362
rect 16710 10310 16762 10362
rect 16774 10310 16826 10362
rect 6552 10251 6604 10260
rect 6552 10217 6561 10251
rect 6561 10217 6595 10251
rect 6595 10217 6604 10251
rect 6552 10208 6604 10217
rect 8208 10208 8260 10260
rect 2412 10140 2464 10192
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 8392 10140 8444 10192
rect 14740 10208 14792 10260
rect 15660 10208 15712 10260
rect 3056 10115 3108 10124
rect 3056 10081 3065 10115
rect 3065 10081 3099 10115
rect 3099 10081 3108 10115
rect 3056 10072 3108 10081
rect 16856 10208 16908 10260
rect 17408 10208 17460 10260
rect 17040 10115 17092 10124
rect 17040 10081 17049 10115
rect 17049 10081 17083 10115
rect 17083 10081 17092 10115
rect 17040 10072 17092 10081
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 1952 10047 2004 10056
rect 1952 10013 1961 10047
rect 1961 10013 1995 10047
rect 1995 10013 2004 10047
rect 1952 10004 2004 10013
rect 2688 10004 2740 10056
rect 4436 10004 4488 10056
rect 4712 9936 4764 9988
rect 6828 10004 6880 10056
rect 10140 10047 10192 10056
rect 10140 10013 10158 10047
rect 10158 10013 10192 10047
rect 10416 10047 10468 10056
rect 10140 10004 10192 10013
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 11520 10004 11572 10056
rect 12900 10004 12952 10056
rect 1400 9868 1452 9920
rect 1860 9868 1912 9920
rect 2872 9868 2924 9920
rect 5908 9911 5960 9920
rect 5908 9877 5917 9911
rect 5917 9877 5951 9911
rect 5951 9877 5960 9911
rect 5908 9868 5960 9877
rect 7380 9936 7432 9988
rect 13084 9936 13136 9988
rect 14188 9868 14240 9920
rect 16396 9868 16448 9920
rect 17500 9911 17552 9920
rect 17500 9877 17509 9911
rect 17509 9877 17543 9911
rect 17543 9877 17552 9911
rect 17500 9868 17552 9877
rect 18512 9868 18564 9920
rect 5398 9766 5450 9818
rect 5462 9766 5514 9818
rect 5526 9766 5578 9818
rect 5590 9766 5642 9818
rect 5654 9766 5706 9818
rect 9846 9766 9898 9818
rect 9910 9766 9962 9818
rect 9974 9766 10026 9818
rect 10038 9766 10090 9818
rect 10102 9766 10154 9818
rect 14294 9766 14346 9818
rect 14358 9766 14410 9818
rect 14422 9766 14474 9818
rect 14486 9766 14538 9818
rect 14550 9766 14602 9818
rect 4160 9664 4212 9716
rect 16028 9664 16080 9716
rect 2688 9596 2740 9648
rect 1952 9528 2004 9580
rect 2228 9528 2280 9580
rect 2504 9528 2556 9580
rect 2320 9460 2372 9512
rect 6552 9596 6604 9648
rect 4068 9528 4120 9580
rect 7104 9528 7156 9580
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 8024 9528 8076 9580
rect 5816 9503 5868 9512
rect 2872 9392 2924 9444
rect 4528 9392 4580 9444
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 5816 9460 5868 9469
rect 6828 9460 6880 9512
rect 9588 9596 9640 9648
rect 10416 9596 10468 9648
rect 11520 9596 11572 9648
rect 14832 9596 14884 9648
rect 8668 9528 8720 9580
rect 6092 9324 6144 9376
rect 6184 9324 6236 9376
rect 16120 9528 16172 9580
rect 17684 9571 17736 9580
rect 17684 9537 17693 9571
rect 17693 9537 17727 9571
rect 17727 9537 17736 9571
rect 17684 9528 17736 9537
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 13820 9460 13872 9512
rect 17960 9460 18012 9512
rect 9680 9392 9732 9444
rect 9772 9324 9824 9376
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 14648 9324 14700 9376
rect 16856 9324 16908 9376
rect 18052 9367 18104 9376
rect 18052 9333 18061 9367
rect 18061 9333 18095 9367
rect 18095 9333 18104 9367
rect 18052 9324 18104 9333
rect 18420 9367 18472 9376
rect 18420 9333 18429 9367
rect 18429 9333 18463 9367
rect 18463 9333 18472 9367
rect 18420 9324 18472 9333
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 3430 9222 3482 9274
rect 7622 9222 7674 9274
rect 7686 9222 7738 9274
rect 7750 9222 7802 9274
rect 7814 9222 7866 9274
rect 7878 9222 7930 9274
rect 12070 9222 12122 9274
rect 12134 9222 12186 9274
rect 12198 9222 12250 9274
rect 12262 9222 12314 9274
rect 12326 9222 12378 9274
rect 16518 9222 16570 9274
rect 16582 9222 16634 9274
rect 16646 9222 16698 9274
rect 16710 9222 16762 9274
rect 16774 9222 16826 9274
rect 1952 9120 2004 9172
rect 2504 9163 2556 9172
rect 2504 9129 2513 9163
rect 2513 9129 2547 9163
rect 2547 9129 2556 9163
rect 2504 9120 2556 9129
rect 4252 9120 4304 9172
rect 6184 9120 6236 9172
rect 7380 9120 7432 9172
rect 7564 9120 7616 9172
rect 9680 9120 9732 9172
rect 10232 9120 10284 9172
rect 3148 9052 3200 9104
rect 3976 9052 4028 9104
rect 11336 9120 11388 9172
rect 12624 9120 12676 9172
rect 14740 9120 14792 9172
rect 16212 9120 16264 9172
rect 16396 9163 16448 9172
rect 16396 9129 16405 9163
rect 16405 9129 16439 9163
rect 16439 9129 16448 9163
rect 16396 9120 16448 9129
rect 17960 9120 18012 9172
rect 16120 9052 16172 9104
rect 17132 9052 17184 9104
rect 2504 8984 2556 9036
rect 11520 9027 11572 9036
rect 3608 8916 3660 8968
rect 3976 8916 4028 8968
rect 4436 8848 4488 8900
rect 4988 8848 5040 8900
rect 5724 8891 5776 8900
rect 5724 8857 5758 8891
rect 5758 8857 5776 8891
rect 5724 8848 5776 8857
rect 5816 8848 5868 8900
rect 6828 8916 6880 8968
rect 11520 8993 11529 9027
rect 11529 8993 11563 9027
rect 11563 8993 11572 9027
rect 11520 8984 11572 8993
rect 16028 9027 16080 9036
rect 16028 8993 16037 9027
rect 16037 8993 16071 9027
rect 16071 8993 16080 9027
rect 16028 8984 16080 8993
rect 2964 8823 3016 8832
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 4160 8780 4212 8832
rect 5172 8780 5224 8832
rect 7104 8848 7156 8900
rect 9772 8916 9824 8968
rect 13268 8916 13320 8968
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 16856 8916 16908 8968
rect 6092 8780 6144 8832
rect 8668 8780 8720 8832
rect 13452 8848 13504 8900
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 15108 8780 15160 8789
rect 15476 8823 15528 8832
rect 15476 8789 15485 8823
rect 15485 8789 15519 8823
rect 15519 8789 15528 8823
rect 15476 8780 15528 8789
rect 16120 8780 16172 8832
rect 16396 8780 16448 8832
rect 17776 8780 17828 8832
rect 5398 8678 5450 8730
rect 5462 8678 5514 8730
rect 5526 8678 5578 8730
rect 5590 8678 5642 8730
rect 5654 8678 5706 8730
rect 9846 8678 9898 8730
rect 9910 8678 9962 8730
rect 9974 8678 10026 8730
rect 10038 8678 10090 8730
rect 10102 8678 10154 8730
rect 14294 8678 14346 8730
rect 14358 8678 14410 8730
rect 14422 8678 14474 8730
rect 14486 8678 14538 8730
rect 14550 8678 14602 8730
rect 2228 8576 2280 8628
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 1952 8415 2004 8424
rect 1952 8381 1961 8415
rect 1961 8381 1995 8415
rect 1995 8381 2004 8415
rect 1952 8372 2004 8381
rect 9772 8576 9824 8628
rect 4252 8508 4304 8560
rect 4896 8508 4948 8560
rect 3148 8440 3200 8492
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 2780 8372 2832 8424
rect 3608 8415 3660 8424
rect 1768 8304 1820 8356
rect 2228 8304 2280 8356
rect 2504 8304 2556 8356
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 5816 8440 5868 8492
rect 6828 8508 6880 8560
rect 9404 8508 9456 8560
rect 14832 8576 14884 8628
rect 16304 8619 16356 8628
rect 16304 8585 16313 8619
rect 16313 8585 16347 8619
rect 16347 8585 16356 8619
rect 16304 8576 16356 8585
rect 17040 8576 17092 8628
rect 11520 8483 11572 8492
rect 11520 8449 11529 8483
rect 11529 8449 11563 8483
rect 11563 8449 11572 8483
rect 11520 8440 11572 8449
rect 11612 8440 11664 8492
rect 16028 8508 16080 8560
rect 4436 8372 4488 8424
rect 14556 8372 14608 8424
rect 14740 8372 14792 8424
rect 16028 8415 16080 8424
rect 6092 8347 6144 8356
rect 6092 8313 6101 8347
rect 6101 8313 6135 8347
rect 6135 8313 6144 8347
rect 6092 8304 6144 8313
rect 15200 8347 15252 8356
rect 2964 8236 3016 8288
rect 5724 8236 5776 8288
rect 8576 8236 8628 8288
rect 10416 8279 10468 8288
rect 10416 8245 10425 8279
rect 10425 8245 10459 8279
rect 10459 8245 10468 8279
rect 10416 8236 10468 8245
rect 15200 8313 15209 8347
rect 15209 8313 15243 8347
rect 15243 8313 15252 8347
rect 16028 8381 16037 8415
rect 16037 8381 16071 8415
rect 16071 8381 16080 8415
rect 16028 8372 16080 8381
rect 15200 8304 15252 8313
rect 17684 8304 17736 8356
rect 14740 8236 14792 8288
rect 15384 8279 15436 8288
rect 15384 8245 15393 8279
rect 15393 8245 15427 8279
rect 15427 8245 15436 8279
rect 15384 8236 15436 8245
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 3430 8134 3482 8186
rect 7622 8134 7674 8186
rect 7686 8134 7738 8186
rect 7750 8134 7802 8186
rect 7814 8134 7866 8186
rect 7878 8134 7930 8186
rect 12070 8134 12122 8186
rect 12134 8134 12186 8186
rect 12198 8134 12250 8186
rect 12262 8134 12314 8186
rect 12326 8134 12378 8186
rect 16518 8134 16570 8186
rect 16582 8134 16634 8186
rect 16646 8134 16698 8186
rect 16710 8134 16762 8186
rect 16774 8134 16826 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 1584 8032 1636 8084
rect 1952 8032 2004 8084
rect 14740 8032 14792 8084
rect 18052 8032 18104 8084
rect 1676 7964 1728 8016
rect 1492 7896 1544 7948
rect 4528 7964 4580 8016
rect 16948 8007 17000 8016
rect 16948 7973 16957 8007
rect 16957 7973 16991 8007
rect 16991 7973 17000 8007
rect 16948 7964 17000 7973
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 14832 7896 14884 7948
rect 15384 7896 15436 7948
rect 2964 7828 3016 7880
rect 4436 7828 4488 7880
rect 8300 7828 8352 7880
rect 10600 7828 10652 7880
rect 2412 7760 2464 7812
rect 2688 7760 2740 7812
rect 4160 7760 4212 7812
rect 7472 7760 7524 7812
rect 10416 7760 10468 7812
rect 13268 7760 13320 7812
rect 15476 7828 15528 7880
rect 16120 7760 16172 7812
rect 2136 7692 2188 7744
rect 2780 7692 2832 7744
rect 3884 7692 3936 7744
rect 5632 7692 5684 7744
rect 6092 7692 6144 7744
rect 8484 7692 8536 7744
rect 9312 7692 9364 7744
rect 12256 7692 12308 7744
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 14556 7692 14608 7744
rect 14740 7692 14792 7744
rect 15384 7692 15436 7744
rect 17224 7735 17276 7744
rect 17224 7701 17233 7735
rect 17233 7701 17267 7735
rect 17267 7701 17276 7735
rect 17224 7692 17276 7701
rect 5398 7590 5450 7642
rect 5462 7590 5514 7642
rect 5526 7590 5578 7642
rect 5590 7590 5642 7642
rect 5654 7590 5706 7642
rect 9846 7590 9898 7642
rect 9910 7590 9962 7642
rect 9974 7590 10026 7642
rect 10038 7590 10090 7642
rect 10102 7590 10154 7642
rect 14294 7590 14346 7642
rect 14358 7590 14410 7642
rect 14422 7590 14474 7642
rect 14486 7590 14538 7642
rect 14550 7590 14602 7642
rect 1492 7488 1544 7540
rect 2136 7531 2188 7540
rect 2136 7497 2145 7531
rect 2145 7497 2179 7531
rect 2179 7497 2188 7531
rect 2136 7488 2188 7497
rect 2780 7488 2832 7540
rect 3608 7488 3660 7540
rect 3792 7488 3844 7540
rect 3976 7488 4028 7540
rect 4528 7488 4580 7540
rect 14188 7488 14240 7540
rect 15384 7531 15436 7540
rect 15384 7497 15393 7531
rect 15393 7497 15427 7531
rect 15427 7497 15436 7531
rect 15384 7488 15436 7497
rect 17132 7531 17184 7540
rect 17132 7497 17141 7531
rect 17141 7497 17175 7531
rect 17175 7497 17184 7531
rect 17132 7488 17184 7497
rect 1676 7420 1728 7472
rect 2228 7352 2280 7404
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 4436 7420 4488 7472
rect 2780 7148 2832 7200
rect 3608 7352 3660 7404
rect 5172 7352 5224 7404
rect 5632 7395 5684 7404
rect 6460 7420 6512 7472
rect 6736 7420 6788 7472
rect 11888 7420 11940 7472
rect 5632 7361 5650 7395
rect 5650 7361 5684 7395
rect 5632 7352 5684 7361
rect 8024 7352 8076 7404
rect 9312 7352 9364 7404
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 11980 7352 12032 7404
rect 14924 7352 14976 7404
rect 15476 7352 15528 7404
rect 4436 7327 4488 7336
rect 4436 7293 4445 7327
rect 4445 7293 4479 7327
rect 4479 7293 4488 7327
rect 4436 7284 4488 7293
rect 8300 7284 8352 7336
rect 15844 7284 15896 7336
rect 16396 7327 16448 7336
rect 16396 7293 16405 7327
rect 16405 7293 16439 7327
rect 16439 7293 16448 7327
rect 18052 7352 18104 7404
rect 16396 7284 16448 7293
rect 4160 7148 4212 7200
rect 4988 7148 5040 7200
rect 5172 7148 5224 7200
rect 7472 7148 7524 7200
rect 9404 7148 9456 7200
rect 10232 7148 10284 7200
rect 16212 7216 16264 7268
rect 13820 7148 13872 7200
rect 17132 7148 17184 7200
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 18052 7148 18104 7157
rect 18420 7191 18472 7200
rect 18420 7157 18429 7191
rect 18429 7157 18463 7191
rect 18463 7157 18472 7191
rect 18420 7148 18472 7157
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 3430 7046 3482 7098
rect 7622 7046 7674 7098
rect 7686 7046 7738 7098
rect 7750 7046 7802 7098
rect 7814 7046 7866 7098
rect 7878 7046 7930 7098
rect 12070 7046 12122 7098
rect 12134 7046 12186 7098
rect 12198 7046 12250 7098
rect 12262 7046 12314 7098
rect 12326 7046 12378 7098
rect 16518 7046 16570 7098
rect 16582 7046 16634 7098
rect 16646 7046 16698 7098
rect 16710 7046 16762 7098
rect 16774 7046 16826 7098
rect 1676 6944 1728 6996
rect 2228 6944 2280 6996
rect 5816 6987 5868 6996
rect 1492 6876 1544 6928
rect 5816 6953 5825 6987
rect 5825 6953 5859 6987
rect 5859 6953 5868 6987
rect 5816 6944 5868 6953
rect 11980 6944 12032 6996
rect 1952 6740 2004 6792
rect 2964 6808 3016 6860
rect 3976 6808 4028 6860
rect 6276 6876 6328 6928
rect 4252 6740 4304 6792
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 6828 6740 6880 6792
rect 8392 6740 8444 6792
rect 9404 6740 9456 6792
rect 3608 6672 3660 6724
rect 6184 6672 6236 6724
rect 11336 6740 11388 6792
rect 1584 6604 1636 6656
rect 2964 6604 3016 6656
rect 3148 6604 3200 6656
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 4344 6604 4396 6656
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 10416 6604 10468 6656
rect 10784 6604 10836 6656
rect 11980 6672 12032 6724
rect 15476 6944 15528 6996
rect 18144 6987 18196 6996
rect 18144 6953 18153 6987
rect 18153 6953 18187 6987
rect 18187 6953 18196 6987
rect 18144 6944 18196 6953
rect 14832 6876 14884 6928
rect 15108 6808 15160 6860
rect 16212 6851 16264 6860
rect 16212 6817 16221 6851
rect 16221 6817 16255 6851
rect 16255 6817 16264 6851
rect 16212 6808 16264 6817
rect 17132 6851 17184 6860
rect 15476 6740 15528 6792
rect 17132 6817 17141 6851
rect 17141 6817 17175 6851
rect 17175 6817 17184 6851
rect 17132 6808 17184 6817
rect 17040 6783 17092 6792
rect 17040 6749 17049 6783
rect 17049 6749 17083 6783
rect 17083 6749 17092 6783
rect 17040 6740 17092 6749
rect 17316 6740 17368 6792
rect 13084 6604 13136 6656
rect 16028 6672 16080 6724
rect 14096 6604 14148 6656
rect 14832 6604 14884 6656
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 5398 6502 5450 6554
rect 5462 6502 5514 6554
rect 5526 6502 5578 6554
rect 5590 6502 5642 6554
rect 5654 6502 5706 6554
rect 9846 6502 9898 6554
rect 9910 6502 9962 6554
rect 9974 6502 10026 6554
rect 10038 6502 10090 6554
rect 10102 6502 10154 6554
rect 14294 6502 14346 6554
rect 14358 6502 14410 6554
rect 14422 6502 14474 6554
rect 14486 6502 14538 6554
rect 14550 6502 14602 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 4252 6443 4304 6452
rect 4252 6409 4261 6443
rect 4261 6409 4295 6443
rect 4295 6409 4304 6443
rect 4252 6400 4304 6409
rect 6552 6400 6604 6452
rect 6736 6400 6788 6452
rect 13084 6400 13136 6452
rect 13268 6443 13320 6452
rect 13268 6409 13277 6443
rect 13277 6409 13311 6443
rect 13311 6409 13320 6443
rect 13268 6400 13320 6409
rect 16028 6400 16080 6452
rect 16948 6443 17000 6452
rect 4436 6332 4488 6384
rect 2228 6307 2280 6316
rect 2228 6273 2237 6307
rect 2237 6273 2271 6307
rect 2271 6273 2280 6307
rect 2228 6264 2280 6273
rect 3792 6264 3844 6316
rect 4068 6264 4120 6316
rect 2412 6196 2464 6248
rect 2688 6196 2740 6248
rect 2780 6196 2832 6248
rect 3516 6239 3568 6248
rect 3516 6205 3525 6239
rect 3525 6205 3559 6239
rect 3559 6205 3568 6239
rect 3516 6196 3568 6205
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 4160 6196 4212 6248
rect 4344 6239 4396 6248
rect 4344 6205 4353 6239
rect 4353 6205 4387 6239
rect 4387 6205 4396 6239
rect 4344 6196 4396 6205
rect 5632 6264 5684 6316
rect 5908 6307 5960 6316
rect 5908 6273 5926 6307
rect 5926 6273 5960 6307
rect 5908 6264 5960 6273
rect 8300 6332 8352 6384
rect 2964 6128 3016 6180
rect 4068 6128 4120 6180
rect 6552 6196 6604 6248
rect 10140 6264 10192 6316
rect 12348 6332 12400 6384
rect 13176 6264 13228 6316
rect 15752 6332 15804 6384
rect 16948 6409 16957 6443
rect 16957 6409 16991 6443
rect 16991 6409 17000 6443
rect 16948 6400 17000 6409
rect 16856 6332 16908 6384
rect 1952 6060 2004 6112
rect 2780 6103 2832 6112
rect 2780 6069 2789 6103
rect 2789 6069 2823 6103
rect 2823 6069 2832 6103
rect 2780 6060 2832 6069
rect 3148 6060 3200 6112
rect 4344 6060 4396 6112
rect 4712 6060 4764 6112
rect 5816 6060 5868 6112
rect 6736 6128 6788 6180
rect 13452 6196 13504 6248
rect 15108 6264 15160 6316
rect 16396 6264 16448 6316
rect 15476 6196 15528 6248
rect 15660 6239 15712 6248
rect 15660 6205 15669 6239
rect 15669 6205 15703 6239
rect 15703 6205 15712 6239
rect 15660 6196 15712 6205
rect 15752 6239 15804 6248
rect 15752 6205 15761 6239
rect 15761 6205 15795 6239
rect 15795 6205 15804 6239
rect 15752 6196 15804 6205
rect 17132 6196 17184 6248
rect 13084 6128 13136 6180
rect 14832 6128 14884 6180
rect 18144 6128 18196 6180
rect 8024 6060 8076 6112
rect 8852 6103 8904 6112
rect 8852 6069 8861 6103
rect 8861 6069 8895 6103
rect 8895 6069 8904 6103
rect 8852 6060 8904 6069
rect 12992 6060 13044 6112
rect 15200 6060 15252 6112
rect 16028 6103 16080 6112
rect 16028 6069 16037 6103
rect 16037 6069 16071 6103
rect 16071 6069 16080 6103
rect 16028 6060 16080 6069
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 3430 5958 3482 6010
rect 7622 5958 7674 6010
rect 7686 5958 7738 6010
rect 7750 5958 7802 6010
rect 7814 5958 7866 6010
rect 7878 5958 7930 6010
rect 12070 5958 12122 6010
rect 12134 5958 12186 6010
rect 12198 5958 12250 6010
rect 12262 5958 12314 6010
rect 12326 5958 12378 6010
rect 16518 5958 16570 6010
rect 16582 5958 16634 6010
rect 16646 5958 16698 6010
rect 16710 5958 16762 6010
rect 16774 5958 16826 6010
rect 2964 5788 3016 5840
rect 3148 5788 3200 5840
rect 3516 5856 3568 5908
rect 3700 5856 3752 5908
rect 3884 5856 3936 5908
rect 3792 5788 3844 5840
rect 5724 5856 5776 5908
rect 6184 5856 6236 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 15108 5899 15160 5908
rect 15108 5865 15117 5899
rect 15117 5865 15151 5899
rect 15151 5865 15160 5899
rect 15108 5856 15160 5865
rect 15660 5856 15712 5908
rect 16396 5899 16448 5908
rect 16396 5865 16405 5899
rect 16405 5865 16439 5899
rect 16439 5865 16448 5899
rect 16396 5856 16448 5865
rect 17500 5899 17552 5908
rect 17500 5865 17509 5899
rect 17509 5865 17543 5899
rect 17543 5865 17552 5899
rect 17500 5856 17552 5865
rect 18052 5899 18104 5908
rect 18052 5865 18061 5899
rect 18061 5865 18095 5899
rect 18095 5865 18104 5899
rect 18052 5856 18104 5865
rect 6276 5788 6328 5840
rect 7380 5788 7432 5840
rect 8116 5788 8168 5840
rect 1952 5763 2004 5772
rect 1952 5729 1961 5763
rect 1961 5729 1995 5763
rect 1995 5729 2004 5763
rect 1952 5720 2004 5729
rect 1860 5695 1912 5704
rect 1860 5661 1869 5695
rect 1869 5661 1903 5695
rect 1903 5661 1912 5695
rect 1860 5652 1912 5661
rect 4068 5720 4120 5772
rect 4436 5720 4488 5772
rect 5908 5720 5960 5772
rect 12992 5788 13044 5840
rect 13176 5788 13228 5840
rect 6092 5652 6144 5704
rect 12808 5720 12860 5772
rect 15752 5788 15804 5840
rect 16304 5788 16356 5840
rect 15292 5720 15344 5772
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 7472 5695 7524 5704
rect 3148 5627 3200 5636
rect 3148 5593 3157 5627
rect 3157 5593 3191 5627
rect 3191 5593 3200 5627
rect 3148 5584 3200 5593
rect 1676 5516 1728 5568
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 3700 5516 3752 5568
rect 4344 5516 4396 5568
rect 4712 5584 4764 5636
rect 7472 5661 7481 5695
rect 7481 5661 7515 5695
rect 7515 5661 7524 5695
rect 7472 5652 7524 5661
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 11980 5652 12032 5704
rect 14188 5652 14240 5704
rect 14740 5695 14792 5704
rect 14740 5661 14749 5695
rect 14749 5661 14783 5695
rect 14783 5661 14792 5695
rect 14740 5652 14792 5661
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 16856 5695 16908 5704
rect 16856 5661 16865 5695
rect 16865 5661 16899 5695
rect 16899 5661 16908 5695
rect 16856 5652 16908 5661
rect 17500 5652 17552 5704
rect 6184 5559 6236 5568
rect 6184 5525 6193 5559
rect 6193 5525 6227 5559
rect 6227 5525 6236 5559
rect 6184 5516 6236 5525
rect 6276 5516 6328 5568
rect 7380 5559 7432 5568
rect 7380 5525 7389 5559
rect 7389 5525 7423 5559
rect 7423 5525 7432 5559
rect 7380 5516 7432 5525
rect 9220 5559 9272 5568
rect 9220 5525 9229 5559
rect 9229 5525 9263 5559
rect 9263 5525 9272 5559
rect 9220 5516 9272 5525
rect 11244 5584 11296 5636
rect 12624 5627 12676 5636
rect 12624 5593 12633 5627
rect 12633 5593 12667 5627
rect 12667 5593 12676 5627
rect 12624 5584 12676 5593
rect 13360 5584 13412 5636
rect 16304 5584 16356 5636
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 17500 5516 17552 5568
rect 18144 5652 18196 5704
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 5398 5414 5450 5466
rect 5462 5414 5514 5466
rect 5526 5414 5578 5466
rect 5590 5414 5642 5466
rect 5654 5414 5706 5466
rect 9846 5414 9898 5466
rect 9910 5414 9962 5466
rect 9974 5414 10026 5466
rect 10038 5414 10090 5466
rect 10102 5414 10154 5466
rect 14294 5414 14346 5466
rect 14358 5414 14410 5466
rect 14422 5414 14474 5466
rect 14486 5414 14538 5466
rect 14550 5414 14602 5466
rect 1860 5312 1912 5364
rect 2136 5312 2188 5364
rect 2228 5312 2280 5364
rect 3884 5312 3936 5364
rect 2320 5176 2372 5228
rect 3792 5176 3844 5228
rect 6184 5244 6236 5296
rect 6552 5312 6604 5364
rect 6828 5312 6880 5364
rect 7104 5244 7156 5296
rect 3608 5108 3660 5160
rect 1952 5015 2004 5024
rect 1952 4981 1961 5015
rect 1961 4981 1995 5015
rect 1995 4981 2004 5015
rect 1952 4972 2004 4981
rect 7472 5176 7524 5228
rect 4068 5151 4120 5160
rect 4068 5117 4077 5151
rect 4077 5117 4111 5151
rect 4111 5117 4120 5151
rect 4712 5151 4764 5160
rect 4068 5108 4120 5117
rect 4712 5117 4721 5151
rect 4721 5117 4755 5151
rect 4755 5117 4764 5151
rect 4712 5108 4764 5117
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 6092 5108 6144 5160
rect 6644 5108 6696 5160
rect 7104 5108 7156 5160
rect 8116 5219 8168 5228
rect 8116 5185 8125 5219
rect 8125 5185 8159 5219
rect 8159 5185 8168 5219
rect 8116 5176 8168 5185
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 9404 5219 9456 5228
rect 9404 5185 9413 5219
rect 9413 5185 9447 5219
rect 9447 5185 9456 5219
rect 9404 5176 9456 5185
rect 9588 5108 9640 5160
rect 9680 5151 9732 5160
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 9772 5040 9824 5092
rect 11152 5312 11204 5364
rect 12624 5312 12676 5364
rect 13728 5312 13780 5364
rect 14372 5312 14424 5364
rect 11796 5244 11848 5296
rect 15200 5312 15252 5364
rect 15292 5355 15344 5364
rect 15292 5321 15301 5355
rect 15301 5321 15335 5355
rect 15335 5321 15344 5355
rect 17592 5355 17644 5364
rect 15292 5312 15344 5321
rect 17592 5321 17601 5355
rect 17601 5321 17635 5355
rect 17635 5321 17644 5355
rect 17592 5312 17644 5321
rect 15384 5244 15436 5296
rect 16028 5244 16080 5296
rect 10416 5219 10468 5228
rect 10416 5185 10425 5219
rect 10425 5185 10459 5219
rect 10459 5185 10468 5219
rect 10416 5176 10468 5185
rect 11060 5176 11112 5228
rect 11888 5108 11940 5160
rect 4436 5015 4488 5024
rect 4436 4981 4445 5015
rect 4445 4981 4479 5015
rect 4479 4981 4488 5015
rect 4436 4972 4488 4981
rect 5724 4972 5776 5024
rect 6736 4972 6788 5024
rect 6920 4972 6972 5024
rect 11336 4972 11388 5024
rect 14188 5151 14240 5160
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 15936 5176 15988 5228
rect 16212 5176 16264 5228
rect 16856 5176 16908 5228
rect 14832 5040 14884 5092
rect 16028 5108 16080 5160
rect 13544 4972 13596 5024
rect 15752 5040 15804 5092
rect 16304 5015 16356 5024
rect 16304 4981 16313 5015
rect 16313 4981 16347 5015
rect 16347 4981 16356 5015
rect 16304 4972 16356 4981
rect 16856 5015 16908 5024
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 17960 5015 18012 5024
rect 17960 4981 17969 5015
rect 17969 4981 18003 5015
rect 18003 4981 18012 5015
rect 17960 4972 18012 4981
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 3430 4870 3482 4922
rect 7622 4870 7674 4922
rect 7686 4870 7738 4922
rect 7750 4870 7802 4922
rect 7814 4870 7866 4922
rect 7878 4870 7930 4922
rect 12070 4870 12122 4922
rect 12134 4870 12186 4922
rect 12198 4870 12250 4922
rect 12262 4870 12314 4922
rect 12326 4870 12378 4922
rect 16518 4870 16570 4922
rect 16582 4870 16634 4922
rect 16646 4870 16698 4922
rect 16710 4870 16762 4922
rect 16774 4870 16826 4922
rect 2228 4743 2280 4752
rect 2228 4709 2237 4743
rect 2237 4709 2271 4743
rect 2271 4709 2280 4743
rect 2228 4700 2280 4709
rect 1860 4564 1912 4616
rect 5816 4768 5868 4820
rect 7104 4768 7156 4820
rect 3792 4700 3844 4752
rect 4436 4700 4488 4752
rect 13544 4768 13596 4820
rect 13636 4768 13688 4820
rect 14280 4811 14332 4820
rect 14280 4777 14289 4811
rect 14289 4777 14323 4811
rect 14323 4777 14332 4811
rect 14280 4768 14332 4777
rect 14464 4768 14516 4820
rect 14740 4768 14792 4820
rect 15752 4768 15804 4820
rect 16212 4768 16264 4820
rect 3700 4632 3752 4684
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 5724 4675 5776 4684
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 14096 4700 14148 4752
rect 15384 4700 15436 4752
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 1584 4428 1636 4480
rect 3884 4564 3936 4616
rect 4712 4564 4764 4616
rect 7472 4632 7524 4684
rect 8024 4632 8076 4684
rect 9220 4564 9272 4616
rect 9772 4632 9824 4684
rect 10232 4564 10284 4616
rect 10784 4632 10836 4684
rect 10968 4675 11020 4684
rect 10968 4641 10977 4675
rect 10977 4641 11011 4675
rect 11011 4641 11020 4675
rect 10968 4632 11020 4641
rect 12072 4632 12124 4684
rect 12532 4632 12584 4684
rect 11888 4564 11940 4616
rect 17408 4632 17460 4684
rect 6092 4428 6144 4480
rect 8116 4496 8168 4548
rect 10784 4539 10836 4548
rect 6644 4471 6696 4480
rect 6644 4437 6653 4471
rect 6653 4437 6687 4471
rect 6687 4437 6696 4471
rect 6644 4428 6696 4437
rect 6828 4428 6880 4480
rect 8208 4428 8260 4480
rect 9128 4428 9180 4480
rect 10784 4505 10793 4539
rect 10793 4505 10827 4539
rect 10827 4505 10836 4539
rect 10784 4496 10836 4505
rect 11060 4539 11112 4548
rect 11060 4505 11069 4539
rect 11069 4505 11103 4539
rect 11103 4505 11112 4539
rect 11060 4496 11112 4505
rect 14280 4564 14332 4616
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 11152 4428 11204 4480
rect 11796 4428 11848 4480
rect 13728 4428 13780 4480
rect 14924 4539 14976 4548
rect 14924 4505 14933 4539
rect 14933 4505 14967 4539
rect 14967 4505 14976 4539
rect 14924 4496 14976 4505
rect 17132 4496 17184 4548
rect 16028 4428 16080 4480
rect 17776 4428 17828 4480
rect 5398 4326 5450 4378
rect 5462 4326 5514 4378
rect 5526 4326 5578 4378
rect 5590 4326 5642 4378
rect 5654 4326 5706 4378
rect 9846 4326 9898 4378
rect 9910 4326 9962 4378
rect 9974 4326 10026 4378
rect 10038 4326 10090 4378
rect 10102 4326 10154 4378
rect 14294 4326 14346 4378
rect 14358 4326 14410 4378
rect 14422 4326 14474 4378
rect 14486 4326 14538 4378
rect 14550 4326 14602 4378
rect 5908 4224 5960 4276
rect 6552 4224 6604 4276
rect 8116 4224 8168 4276
rect 8208 4224 8260 4276
rect 11060 4224 11112 4276
rect 6644 4156 6696 4208
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 3056 4131 3108 4140
rect 1860 4063 1912 4072
rect 1860 4029 1869 4063
rect 1869 4029 1903 4063
rect 1903 4029 1912 4063
rect 1860 4020 1912 4029
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 9128 4199 9180 4208
rect 9128 4165 9137 4199
rect 9137 4165 9171 4199
rect 9171 4165 9180 4199
rect 9128 4156 9180 4165
rect 9588 4156 9640 4208
rect 14556 4224 14608 4276
rect 14648 4224 14700 4276
rect 11704 4156 11756 4208
rect 12532 4199 12584 4208
rect 8116 4063 8168 4072
rect 8116 4029 8125 4063
rect 8125 4029 8159 4063
rect 8159 4029 8168 4063
rect 8116 4020 8168 4029
rect 8852 4088 8904 4140
rect 9036 4063 9088 4072
rect 2320 3995 2372 4004
rect 2320 3961 2329 3995
rect 2329 3961 2363 3995
rect 2363 3961 2372 3995
rect 2320 3952 2372 3961
rect 5724 3952 5776 4004
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 10048 4063 10100 4072
rect 10048 4029 10057 4063
rect 10057 4029 10091 4063
rect 10091 4029 10100 4063
rect 10048 4020 10100 4029
rect 10324 4020 10376 4072
rect 11704 4020 11756 4072
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 12532 4165 12541 4199
rect 12541 4165 12575 4199
rect 12575 4165 12584 4199
rect 12532 4156 12584 4165
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 2872 3884 2924 3936
rect 10232 3884 10284 3936
rect 10784 3952 10836 4004
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 14464 3884 14516 3936
rect 14740 3884 14792 3936
rect 17960 3927 18012 3936
rect 17960 3893 17969 3927
rect 17969 3893 18003 3927
rect 18003 3893 18012 3927
rect 17960 3884 18012 3893
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 3430 3782 3482 3834
rect 7622 3782 7674 3834
rect 7686 3782 7738 3834
rect 7750 3782 7802 3834
rect 7814 3782 7866 3834
rect 7878 3782 7930 3834
rect 12070 3782 12122 3834
rect 12134 3782 12186 3834
rect 12198 3782 12250 3834
rect 12262 3782 12314 3834
rect 12326 3782 12378 3834
rect 16518 3782 16570 3834
rect 16582 3782 16634 3834
rect 16646 3782 16698 3834
rect 16710 3782 16762 3834
rect 16774 3782 16826 3834
rect 3424 3680 3476 3732
rect 8208 3680 8260 3732
rect 8944 3723 8996 3732
rect 8944 3689 8953 3723
rect 8953 3689 8987 3723
rect 8987 3689 8996 3723
rect 8944 3680 8996 3689
rect 9036 3680 9088 3732
rect 14096 3680 14148 3732
rect 14924 3680 14976 3732
rect 15752 3723 15804 3732
rect 15752 3689 15761 3723
rect 15761 3689 15795 3723
rect 15795 3689 15804 3723
rect 15752 3680 15804 3689
rect 7288 3544 7340 3596
rect 10048 3612 10100 3664
rect 15476 3612 15528 3664
rect 12992 3544 13044 3596
rect 13360 3544 13412 3596
rect 15016 3587 15068 3596
rect 15016 3553 15025 3587
rect 15025 3553 15059 3587
rect 15059 3553 15068 3587
rect 15016 3544 15068 3553
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 6920 3476 6972 3528
rect 2872 3408 2924 3460
rect 3056 3408 3108 3460
rect 9128 3519 9180 3528
rect 9128 3485 9172 3519
rect 9172 3485 9180 3519
rect 9128 3476 9180 3485
rect 9588 3476 9640 3528
rect 11244 3476 11296 3528
rect 11888 3476 11940 3528
rect 12532 3476 12584 3528
rect 1400 3340 1452 3392
rect 7564 3340 7616 3392
rect 8116 3408 8168 3460
rect 11612 3408 11664 3460
rect 9772 3340 9824 3392
rect 11980 3340 12032 3392
rect 13360 3340 13412 3392
rect 14464 3408 14516 3460
rect 17868 3408 17920 3460
rect 5398 3238 5450 3290
rect 5462 3238 5514 3290
rect 5526 3238 5578 3290
rect 5590 3238 5642 3290
rect 5654 3238 5706 3290
rect 9846 3238 9898 3290
rect 9910 3238 9962 3290
rect 9974 3238 10026 3290
rect 10038 3238 10090 3290
rect 10102 3238 10154 3290
rect 14294 3238 14346 3290
rect 14358 3238 14410 3290
rect 14422 3238 14474 3290
rect 14486 3238 14538 3290
rect 14550 3238 14602 3290
rect 3608 3136 3660 3188
rect 3700 3068 3752 3120
rect 1768 3000 1820 3052
rect 2596 3000 2648 3052
rect 3424 3043 3476 3052
rect 3424 3009 3433 3043
rect 3433 3009 3467 3043
rect 3467 3009 3476 3043
rect 3424 3000 3476 3009
rect 5080 3000 5132 3052
rect 940 2932 992 2984
rect 2320 2932 2372 2984
rect 4620 2975 4672 2984
rect 4620 2941 4629 2975
rect 4629 2941 4663 2975
rect 4663 2941 4672 2975
rect 4620 2932 4672 2941
rect 2780 2796 2832 2848
rect 3516 2796 3568 2848
rect 8116 3136 8168 3188
rect 8668 3136 8720 3188
rect 11796 3136 11848 3188
rect 11888 3136 11940 3188
rect 7564 3068 7616 3120
rect 8760 3111 8812 3120
rect 8760 3077 8769 3111
rect 8769 3077 8803 3111
rect 8803 3077 8812 3111
rect 8760 3068 8812 3077
rect 9312 3111 9364 3120
rect 9312 3077 9321 3111
rect 9321 3077 9355 3111
rect 9355 3077 9364 3111
rect 9312 3068 9364 3077
rect 9772 3068 9824 3120
rect 11244 3068 11296 3120
rect 11704 3111 11756 3120
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 12072 3068 12124 3120
rect 7012 3000 7064 3052
rect 7380 3000 7432 3052
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 10784 3000 10836 3009
rect 12624 3111 12676 3120
rect 12624 3077 12633 3111
rect 12633 3077 12667 3111
rect 12667 3077 12676 3111
rect 12624 3068 12676 3077
rect 13452 3136 13504 3188
rect 14096 3068 14148 3120
rect 14188 3068 14240 3120
rect 14556 3068 14608 3120
rect 14648 3068 14700 3120
rect 15476 3043 15528 3052
rect 15476 3009 15485 3043
rect 15485 3009 15519 3043
rect 15519 3009 15528 3043
rect 15476 3000 15528 3009
rect 16120 3000 16172 3052
rect 17132 3068 17184 3120
rect 17408 3043 17460 3052
rect 17408 3009 17417 3043
rect 17417 3009 17451 3043
rect 17451 3009 17460 3043
rect 17408 3000 17460 3009
rect 17868 3043 17920 3052
rect 17868 3009 17877 3043
rect 17877 3009 17911 3043
rect 17911 3009 17920 3043
rect 17868 3000 17920 3009
rect 9404 2932 9456 2984
rect 11612 2975 11664 2984
rect 11612 2941 11621 2975
rect 11621 2941 11655 2975
rect 11655 2941 11664 2975
rect 11612 2932 11664 2941
rect 11888 2932 11940 2984
rect 14004 2975 14056 2984
rect 6368 2796 6420 2848
rect 6920 2796 6972 2848
rect 7472 2839 7524 2848
rect 7472 2805 7481 2839
rect 7481 2805 7515 2839
rect 7515 2805 7524 2839
rect 7472 2796 7524 2805
rect 10232 2864 10284 2916
rect 11520 2864 11572 2916
rect 11796 2864 11848 2916
rect 13084 2864 13136 2916
rect 8668 2796 8720 2848
rect 8760 2796 8812 2848
rect 10600 2839 10652 2848
rect 10600 2805 10609 2839
rect 10609 2805 10643 2839
rect 10643 2805 10652 2839
rect 10600 2796 10652 2805
rect 14004 2941 14013 2975
rect 14013 2941 14047 2975
rect 14047 2941 14056 2975
rect 14004 2932 14056 2941
rect 13912 2864 13964 2916
rect 14372 2864 14424 2916
rect 15476 2864 15528 2916
rect 13820 2796 13872 2848
rect 18880 2864 18932 2916
rect 15752 2796 15804 2848
rect 16396 2796 16448 2848
rect 17040 2796 17092 2848
rect 17500 2796 17552 2848
rect 17960 2796 18012 2848
rect 18420 2839 18472 2848
rect 18420 2805 18429 2839
rect 18429 2805 18463 2839
rect 18463 2805 18472 2839
rect 18420 2796 18472 2805
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 3430 2694 3482 2746
rect 7622 2694 7674 2746
rect 7686 2694 7738 2746
rect 7750 2694 7802 2746
rect 7814 2694 7866 2746
rect 7878 2694 7930 2746
rect 12070 2694 12122 2746
rect 12134 2694 12186 2746
rect 12198 2694 12250 2746
rect 12262 2694 12314 2746
rect 12326 2694 12378 2746
rect 16518 2694 16570 2746
rect 16582 2694 16634 2746
rect 16646 2694 16698 2746
rect 16710 2694 16762 2746
rect 16774 2694 16826 2746
rect 11704 2592 11756 2644
rect 14464 2592 14516 2644
rect 15476 2635 15528 2644
rect 15476 2601 15485 2635
rect 15485 2601 15519 2635
rect 15519 2601 15528 2635
rect 15476 2592 15528 2601
rect 9680 2524 9732 2576
rect 10876 2524 10928 2576
rect 11060 2524 11112 2576
rect 4896 2388 4948 2440
rect 9128 2388 9180 2440
rect 9496 2388 9548 2440
rect 9772 2388 9824 2440
rect 11704 2456 11756 2508
rect 12900 2499 12952 2508
rect 12900 2465 12909 2499
rect 12909 2465 12943 2499
rect 12943 2465 12952 2499
rect 12900 2456 12952 2465
rect 12992 2456 13044 2508
rect 15200 2524 15252 2576
rect 11152 2431 11204 2440
rect 11152 2397 11170 2431
rect 11170 2397 11204 2431
rect 11152 2388 11204 2397
rect 14096 2388 14148 2440
rect 14832 2431 14884 2440
rect 14832 2397 14841 2431
rect 14841 2397 14875 2431
rect 14875 2397 14884 2431
rect 14832 2388 14884 2397
rect 1400 2320 1452 2372
rect 4160 2320 4212 2372
rect 9404 2363 9456 2372
rect 9404 2329 9413 2363
rect 9413 2329 9447 2363
rect 9447 2329 9456 2363
rect 9404 2320 9456 2329
rect 7380 2252 7432 2304
rect 8300 2252 8352 2304
rect 9496 2252 9548 2304
rect 11060 2252 11112 2304
rect 11980 2363 12032 2372
rect 11980 2329 11989 2363
rect 11989 2329 12023 2363
rect 12023 2329 12032 2363
rect 11980 2320 12032 2329
rect 12440 2252 12492 2304
rect 16120 2320 16172 2372
rect 18052 2295 18104 2304
rect 18052 2261 18061 2295
rect 18061 2261 18095 2295
rect 18095 2261 18104 2295
rect 18052 2252 18104 2261
rect 5398 2150 5450 2202
rect 5462 2150 5514 2202
rect 5526 2150 5578 2202
rect 5590 2150 5642 2202
rect 5654 2150 5706 2202
rect 9846 2150 9898 2202
rect 9910 2150 9962 2202
rect 9974 2150 10026 2202
rect 10038 2150 10090 2202
rect 10102 2150 10154 2202
rect 14294 2150 14346 2202
rect 14358 2150 14410 2202
rect 14422 2150 14474 2202
rect 14486 2150 14538 2202
rect 14550 2150 14602 2202
rect 2780 1708 2832 1760
rect 3056 1708 3108 1760
<< metal2 >>
rect 294 16400 350 17200
rect 938 16538 994 17200
rect 938 16510 1256 16538
rect 938 16400 994 16510
rect 308 13734 336 16400
rect 1228 14414 1256 16510
rect 1582 16400 1638 17200
rect 2226 16400 2282 17200
rect 2870 16400 2926 17200
rect 3054 16416 3110 16425
rect 1216 14408 1268 14414
rect 1216 14350 1268 14356
rect 1596 13802 1624 16400
rect 2240 14482 2268 16400
rect 2778 16280 2834 16289
rect 2778 16215 2834 16224
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2134 13832 2190 13841
rect 1584 13796 1636 13802
rect 2134 13767 2190 13776
rect 1584 13738 1636 13744
rect 296 13728 348 13734
rect 296 13670 348 13676
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 1582 10568 1638 10577
rect 1582 10503 1638 10512
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1412 8129 1440 9862
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1398 8120 1454 8129
rect 1504 8090 1532 8191
rect 1596 8090 1624 10503
rect 1964 10062 1992 10678
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1674 8936 1730 8945
rect 1674 8871 1730 8880
rect 1398 8055 1454 8064
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1504 7954 1532 8026
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1504 7546 1532 7890
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1596 7426 1624 8026
rect 1688 8022 1716 8871
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 1688 7478 1716 7958
rect 1504 7398 1624 7426
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1504 6934 1532 7398
rect 1676 7336 1728 7342
rect 1582 7304 1638 7313
rect 1676 7278 1728 7284
rect 1582 7239 1638 7248
rect 1492 6928 1544 6934
rect 1492 6870 1544 6876
rect 1596 6662 1624 7239
rect 1688 7002 1716 7278
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1582 6488 1638 6497
rect 1582 6423 1584 6432
rect 1636 6423 1638 6432
rect 1584 6394 1636 6400
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1492 4480 1544 4486
rect 1490 4448 1492 4457
rect 1584 4480 1636 4486
rect 1544 4448 1546 4457
rect 1584 4422 1636 4428
rect 1490 4383 1546 4392
rect 1596 3641 1624 4422
rect 1688 4146 1716 5510
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1582 3632 1638 3641
rect 1582 3567 1638 3576
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 940 2984 992 2990
rect 940 2926 992 2932
rect 952 800 980 2926
rect 1412 2825 1440 3334
rect 1780 3058 1808 8298
rect 1872 5710 1900 9862
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1964 9178 1992 9522
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 8090 1992 8366
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2056 6905 2084 12582
rect 2148 8514 2176 13767
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2700 11898 2728 12310
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2504 11756 2556 11762
rect 2792 11744 2820 16215
rect 2884 14346 2912 16400
rect 3514 16400 3570 17200
rect 4158 16400 4214 17200
rect 4802 16400 4858 17200
rect 5446 16538 5502 17200
rect 5276 16510 5502 16538
rect 3054 16351 3110 16360
rect 2962 14648 3018 14657
rect 2962 14583 2964 14592
rect 3016 14583 3018 14592
rect 2964 14554 3016 14560
rect 2872 14340 2924 14346
rect 2872 14282 2924 14288
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2884 12986 2912 13262
rect 3068 12986 3096 16351
rect 3528 14822 3556 16400
rect 3974 15872 4030 15881
rect 3974 15807 4030 15816
rect 3790 15464 3846 15473
rect 3790 15399 3846 15408
rect 3606 15056 3662 15065
rect 3606 14991 3662 15000
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3174 14716 3482 14725
rect 3174 14714 3180 14716
rect 3236 14714 3260 14716
rect 3316 14714 3340 14716
rect 3396 14714 3420 14716
rect 3476 14714 3482 14716
rect 3236 14662 3238 14714
rect 3418 14662 3420 14714
rect 3174 14660 3180 14662
rect 3236 14660 3260 14662
rect 3316 14660 3340 14662
rect 3396 14660 3420 14662
rect 3476 14660 3482 14662
rect 3174 14651 3482 14660
rect 3174 13628 3482 13637
rect 3174 13626 3180 13628
rect 3236 13626 3260 13628
rect 3316 13626 3340 13628
rect 3396 13626 3420 13628
rect 3476 13626 3482 13628
rect 3236 13574 3238 13626
rect 3418 13574 3420 13626
rect 3174 13572 3180 13574
rect 3236 13572 3260 13574
rect 3316 13572 3340 13574
rect 3396 13572 3420 13574
rect 3476 13572 3482 13574
rect 3174 13563 3482 13572
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2884 11762 2912 12650
rect 2976 12442 3004 12854
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3174 12540 3482 12549
rect 3174 12538 3180 12540
rect 3236 12538 3260 12540
rect 3316 12538 3340 12540
rect 3396 12538 3420 12540
rect 3476 12538 3482 12540
rect 3236 12486 3238 12538
rect 3418 12486 3420 12538
rect 3174 12484 3180 12486
rect 3236 12484 3260 12486
rect 3316 12484 3340 12486
rect 3396 12484 3420 12486
rect 3476 12484 3482 12486
rect 3174 12475 3482 12484
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 3148 12368 3200 12374
rect 3148 12310 3200 12316
rect 3160 12170 3188 12310
rect 3148 12164 3200 12170
rect 3148 12106 3200 12112
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3344 11898 3372 12038
rect 3528 11898 3556 12582
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 2504 11698 2556 11704
rect 2700 11716 2820 11744
rect 2872 11756 2924 11762
rect 2516 11354 2544 11698
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2240 9586 2268 10542
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2412 10192 2464 10198
rect 2412 10134 2464 10140
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 8634 2268 9318
rect 2332 8634 2360 9454
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2148 8486 2360 8514
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2148 7546 2176 7686
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2240 7410 2268 8298
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2042 6896 2098 6905
rect 2042 6831 2098 6840
rect 1952 6792 2004 6798
rect 1950 6760 1952 6769
rect 2004 6760 2006 6769
rect 1950 6695 2006 6704
rect 2240 6474 2268 6938
rect 2148 6446 2268 6474
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1964 5778 1992 6054
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 2148 5370 2176 6446
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2240 5370 2268 6258
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 1872 4622 1900 5306
rect 2332 5234 2360 8486
rect 2424 7818 2452 10134
rect 2516 10130 2544 10406
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2516 9178 2544 9522
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2516 8362 2544 8978
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 2412 7812 2464 7818
rect 2412 7754 2464 7760
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2424 5574 2452 6190
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2424 5273 2452 5510
rect 2410 5264 2466 5273
rect 2320 5228 2372 5234
rect 2410 5199 2466 5208
rect 2320 5170 2372 5176
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 1400 2372 1452 2378
rect 1400 2314 1452 2320
rect 1412 800 1440 2314
rect 1872 800 1900 4014
rect 1964 1601 1992 4966
rect 2228 4752 2280 4758
rect 2228 4694 2280 4700
rect 2240 3233 2268 4694
rect 2318 4040 2374 4049
rect 2318 3975 2320 3984
rect 2372 3975 2374 3984
rect 2320 3946 2372 3952
rect 2226 3224 2282 3233
rect 2226 3159 2282 3168
rect 2608 3058 2636 10950
rect 2700 10810 2728 11716
rect 2872 11698 2924 11704
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2700 10713 2728 10746
rect 2686 10704 2742 10713
rect 2686 10639 2742 10648
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2700 10062 2728 10406
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2700 7954 2728 9590
rect 2792 8537 2820 11562
rect 2884 10690 2912 11562
rect 2976 11150 3004 11834
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 3068 11218 3096 11494
rect 3174 11452 3482 11461
rect 3174 11450 3180 11452
rect 3236 11450 3260 11452
rect 3316 11450 3340 11452
rect 3396 11450 3420 11452
rect 3476 11450 3482 11452
rect 3236 11398 3238 11450
rect 3418 11398 3420 11450
rect 3174 11396 3180 11398
rect 3236 11396 3260 11398
rect 3316 11396 3340 11398
rect 3396 11396 3420 11398
rect 3476 11396 3482 11398
rect 3174 11387 3482 11396
rect 3620 11257 3648 14991
rect 3698 12744 3754 12753
rect 3698 12679 3754 12688
rect 3712 12322 3740 12679
rect 3804 12434 3832 15399
rect 3988 13258 4016 15807
rect 4172 14385 4200 16400
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4158 14376 4214 14385
rect 4158 14311 4214 14320
rect 4066 14240 4122 14249
rect 4122 14198 4200 14226
rect 4066 14175 4122 14184
rect 4066 13424 4122 13433
rect 4066 13359 4122 13368
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3896 12889 3924 12922
rect 4080 12918 4108 13359
rect 4068 12912 4120 12918
rect 3882 12880 3938 12889
rect 4068 12854 4120 12860
rect 3882 12815 3938 12824
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 3804 12406 4016 12434
rect 3712 12294 3924 12322
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3606 11248 3662 11257
rect 3056 11212 3108 11218
rect 3606 11183 3662 11192
rect 3056 11154 3108 11160
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 3606 11112 3662 11121
rect 3606 11047 3662 11056
rect 2884 10662 3004 10690
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2884 9926 2912 10542
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2778 8528 2834 8537
rect 2778 8463 2834 8472
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2792 7857 2820 8366
rect 2778 7848 2834 7857
rect 2688 7812 2740 7818
rect 2778 7783 2834 7792
rect 2688 7754 2740 7760
rect 2700 6254 2728 7754
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2792 7546 2820 7686
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 6254 2820 7142
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 4865 2820 6054
rect 2884 5681 2912 9386
rect 2976 8922 3004 10662
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 3068 10130 3096 10610
rect 3174 10364 3482 10373
rect 3174 10362 3180 10364
rect 3236 10362 3260 10364
rect 3316 10362 3340 10364
rect 3396 10362 3420 10364
rect 3476 10362 3482 10364
rect 3236 10310 3238 10362
rect 3418 10310 3420 10362
rect 3174 10308 3180 10310
rect 3236 10308 3260 10310
rect 3316 10308 3340 10310
rect 3396 10308 3420 10310
rect 3476 10308 3482 10310
rect 3174 10299 3482 10308
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 3174 9276 3482 9285
rect 3174 9274 3180 9276
rect 3236 9274 3260 9276
rect 3316 9274 3340 9276
rect 3396 9274 3420 9276
rect 3476 9274 3482 9276
rect 3236 9222 3238 9274
rect 3418 9222 3420 9274
rect 3174 9220 3180 9222
rect 3236 9220 3260 9222
rect 3316 9220 3340 9222
rect 3396 9220 3420 9222
rect 3476 9220 3482 9222
rect 3174 9211 3482 9220
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 2976 8894 3096 8922
rect 2964 8832 3016 8838
rect 2962 8800 2964 8809
rect 3016 8800 3018 8809
rect 2962 8735 3018 8744
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 7886 3004 8230
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2976 6662 3004 6802
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2976 5846 3004 6122
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 2870 5672 2926 5681
rect 2870 5607 2926 5616
rect 3068 5409 3096 8894
rect 3160 8498 3188 9046
rect 3620 8974 3648 11047
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3174 8188 3482 8197
rect 3174 8186 3180 8188
rect 3236 8186 3260 8188
rect 3316 8186 3340 8188
rect 3396 8186 3420 8188
rect 3476 8186 3482 8188
rect 3236 8134 3238 8186
rect 3418 8134 3420 8186
rect 3174 8132 3180 8134
rect 3236 8132 3260 8134
rect 3316 8132 3340 8134
rect 3396 8132 3420 8134
rect 3476 8132 3482 8134
rect 3174 8123 3482 8132
rect 3174 7100 3482 7109
rect 3174 7098 3180 7100
rect 3236 7098 3260 7100
rect 3316 7098 3340 7100
rect 3396 7098 3420 7100
rect 3476 7098 3482 7100
rect 3236 7046 3238 7098
rect 3418 7046 3420 7098
rect 3174 7044 3180 7046
rect 3236 7044 3260 7046
rect 3316 7044 3340 7046
rect 3396 7044 3420 7046
rect 3476 7044 3482 7046
rect 3174 7035 3482 7044
rect 3528 6662 3556 8434
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3620 7546 3648 8366
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3620 6730 3648 7346
rect 3608 6724 3660 6730
rect 3608 6666 3660 6672
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3160 6118 3188 6598
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3608 6248 3660 6254
rect 3712 6225 3740 12174
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3804 7721 3832 11698
rect 3896 10577 3924 12294
rect 3882 10568 3938 10577
rect 3882 10503 3938 10512
rect 3988 9110 4016 12406
rect 4080 12306 4108 12718
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4172 12170 4200 14198
rect 4448 12986 4476 14894
rect 4816 14278 4844 16400
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 5276 13433 5304 16510
rect 5446 16400 5502 16510
rect 6090 16538 6146 17200
rect 6734 16538 6790 17200
rect 6090 16510 6500 16538
rect 6090 16400 6146 16510
rect 5398 14172 5706 14181
rect 5398 14170 5404 14172
rect 5460 14170 5484 14172
rect 5540 14170 5564 14172
rect 5620 14170 5644 14172
rect 5700 14170 5706 14172
rect 5460 14118 5462 14170
rect 5642 14118 5644 14170
rect 5398 14116 5404 14118
rect 5460 14116 5484 14118
rect 5540 14116 5564 14118
rect 5620 14116 5644 14118
rect 5700 14116 5706 14118
rect 5398 14107 5706 14116
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5552 13734 5580 13942
rect 6472 13938 6500 16510
rect 6564 16510 6790 16538
rect 6564 14074 6592 16510
rect 6734 16400 6790 16510
rect 7378 16400 7434 17200
rect 8022 16400 8078 17200
rect 8666 16538 8722 17200
rect 9310 16538 9366 17200
rect 8666 16510 8984 16538
rect 8666 16400 8722 16510
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5262 13424 5318 13433
rect 5262 13359 5318 13368
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5184 12986 5212 13126
rect 5276 12986 5304 13194
rect 5398 13084 5706 13093
rect 5398 13082 5404 13084
rect 5460 13082 5484 13084
rect 5540 13082 5564 13084
rect 5620 13082 5644 13084
rect 5700 13082 5706 13084
rect 5460 13030 5462 13082
rect 5642 13030 5644 13082
rect 5398 13028 5404 13030
rect 5460 13028 5484 13030
rect 5540 13028 5564 13030
rect 5620 13028 5644 13030
rect 5700 13028 5706 13030
rect 5398 13019 5706 13028
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 11898 4384 12038
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4066 11792 4122 11801
rect 4066 11727 4068 11736
rect 4120 11727 4122 11736
rect 4068 11698 4120 11704
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4540 11150 4568 11630
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4068 11008 4120 11014
rect 4066 10976 4068 10985
rect 4120 10976 4122 10985
rect 4066 10911 4122 10920
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4080 10169 4108 10746
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4172 10470 4200 10678
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4066 10160 4122 10169
rect 4066 10095 4122 10104
rect 4172 9722 4200 10406
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4342 9752 4398 9761
rect 4160 9716 4212 9722
rect 4342 9687 4398 9696
rect 4160 9658 4212 9664
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4080 9489 4108 9522
rect 4066 9480 4122 9489
rect 4066 9415 4122 9424
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3884 7744 3936 7750
rect 3790 7712 3846 7721
rect 3884 7686 3936 7692
rect 3790 7647 3846 7656
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3804 6497 3832 7482
rect 3790 6488 3846 6497
rect 3790 6423 3846 6432
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3608 6190 3660 6196
rect 3698 6216 3754 6225
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3174 6012 3482 6021
rect 3174 6010 3180 6012
rect 3236 6010 3260 6012
rect 3316 6010 3340 6012
rect 3396 6010 3420 6012
rect 3476 6010 3482 6012
rect 3236 5958 3238 6010
rect 3418 5958 3420 6010
rect 3174 5956 3180 5958
rect 3236 5956 3260 5958
rect 3316 5956 3340 5958
rect 3396 5956 3420 5958
rect 3476 5956 3482 5958
rect 3174 5947 3482 5956
rect 3528 5914 3556 6190
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3148 5840 3200 5846
rect 3148 5782 3200 5788
rect 3160 5642 3188 5782
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3054 5400 3110 5409
rect 3054 5335 3110 5344
rect 3620 5166 3648 6190
rect 3698 6151 3754 6160
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3712 5574 3740 5850
rect 3804 5846 3832 6258
rect 3896 5914 3924 7686
rect 3988 7546 4016 8910
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 7818 4200 8774
rect 4264 8566 4292 9114
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 4264 7290 4292 8502
rect 4080 7262 4292 7290
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3988 6662 4016 6802
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3882 5808 3938 5817
rect 3882 5743 3938 5752
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3174 4924 3482 4933
rect 3174 4922 3180 4924
rect 3236 4922 3260 4924
rect 3316 4922 3340 4924
rect 3396 4922 3420 4924
rect 3476 4922 3482 4924
rect 3236 4870 3238 4922
rect 3418 4870 3420 4922
rect 3174 4868 3180 4870
rect 3236 4868 3260 4870
rect 3316 4868 3340 4870
rect 3396 4868 3420 4870
rect 3476 4868 3482 4870
rect 2778 4856 2834 4865
rect 3174 4859 3482 4868
rect 2778 4791 2834 4800
rect 3054 4720 3110 4729
rect 3712 4690 3740 5510
rect 3896 5370 3924 5743
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3804 5137 3832 5170
rect 3790 5128 3846 5137
rect 3790 5063 3846 5072
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3054 4655 3110 4664
rect 3700 4684 3752 4690
rect 3068 4146 3096 4655
rect 3700 4626 3752 4632
rect 3238 4176 3294 4185
rect 3056 4140 3108 4146
rect 3238 4111 3240 4120
rect 3056 4082 3108 4088
rect 3292 4111 3294 4120
rect 3240 4082 3292 4088
rect 2872 3936 2924 3942
rect 2924 3884 3004 3890
rect 2872 3878 3004 3884
rect 2884 3862 3004 3878
rect 2688 3528 2740 3534
rect 2686 3496 2688 3505
rect 2740 3496 2742 3505
rect 2686 3431 2742 3440
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 1950 1592 2006 1601
rect 1950 1527 2006 1536
rect 2332 800 2360 2926
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2792 2009 2820 2790
rect 2778 2000 2834 2009
rect 2778 1935 2834 1944
rect 2780 1760 2832 1766
rect 2780 1702 2832 1708
rect 2792 800 2820 1702
rect 938 0 994 800
rect 1398 0 1454 800
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 2884 377 2912 3402
rect 2976 2417 3004 3862
rect 3174 3836 3482 3845
rect 3174 3834 3180 3836
rect 3236 3834 3260 3836
rect 3316 3834 3340 3836
rect 3396 3834 3420 3836
rect 3476 3834 3482 3836
rect 3236 3782 3238 3834
rect 3418 3782 3420 3834
rect 3174 3780 3180 3782
rect 3236 3780 3260 3782
rect 3316 3780 3340 3782
rect 3396 3780 3420 3782
rect 3476 3780 3482 3782
rect 3174 3771 3482 3780
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 2962 2408 3018 2417
rect 2962 2343 3018 2352
rect 3068 1766 3096 3402
rect 3436 3058 3464 3674
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3174 2748 3482 2757
rect 3174 2746 3180 2748
rect 3236 2746 3260 2748
rect 3316 2746 3340 2748
rect 3396 2746 3420 2748
rect 3476 2746 3482 2748
rect 3236 2694 3238 2746
rect 3418 2694 3420 2746
rect 3174 2692 3180 2694
rect 3236 2692 3260 2694
rect 3316 2692 3340 2694
rect 3396 2692 3420 2694
rect 3476 2692 3482 2694
rect 3174 2683 3482 2692
rect 3056 1760 3108 1766
rect 3056 1702 3108 1708
rect 3528 1193 3556 2790
rect 3514 1184 3570 1193
rect 3514 1119 3570 1128
rect 3252 870 3372 898
rect 3252 800 3280 870
rect 2870 368 2926 377
rect 2870 303 2926 312
rect 3238 0 3294 800
rect 3344 762 3372 870
rect 3620 762 3648 3130
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 3712 800 3740 3062
rect 3804 921 3832 4694
rect 3896 4622 3924 5306
rect 3988 4729 4016 6598
rect 4080 6322 4108 7262
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4172 6254 4200 7142
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4264 6458 4292 6734
rect 4356 6662 4384 9687
rect 4448 8906 4476 9998
rect 4540 9450 4568 11086
rect 4724 9994 4752 11154
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4448 8430 4476 8842
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4448 7886 4476 8366
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4448 7478 4476 7822
rect 4540 7546 4568 7958
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 4448 7342 4476 7414
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4448 6798 4476 7278
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4356 6254 4384 6598
rect 4448 6390 4476 6734
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 5778 4108 6122
rect 4356 6118 4384 6190
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 5166 4108 5714
rect 4356 5574 4384 6054
rect 4448 5778 4476 6326
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4724 5642 4752 6054
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4724 5166 4752 5578
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4448 4758 4476 4966
rect 4436 4752 4488 4758
rect 3974 4720 4030 4729
rect 4436 4694 4488 4700
rect 3974 4655 4030 4664
rect 4724 4622 4752 5102
rect 3884 4616 3936 4622
rect 3882 4584 3884 4593
rect 4712 4616 4764 4622
rect 3936 4584 3938 4593
rect 4712 4558 4764 4564
rect 3882 4519 3938 4528
rect 3896 4493 3924 4519
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 3790 912 3846 921
rect 3790 847 3846 856
rect 4172 800 4200 2314
rect 4632 800 4660 2926
rect 4816 2774 4844 12582
rect 5368 12434 5396 12718
rect 5276 12406 5396 12434
rect 5172 12164 5224 12170
rect 5172 12106 5224 12112
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4908 11898 4936 12038
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 8566 4936 10406
rect 5000 8906 5028 10542
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 5000 7206 5028 8842
rect 5184 8838 5212 12106
rect 5276 10470 5304 12406
rect 5398 11996 5706 12005
rect 5398 11994 5404 11996
rect 5460 11994 5484 11996
rect 5540 11994 5564 11996
rect 5620 11994 5644 11996
rect 5700 11994 5706 11996
rect 5460 11942 5462 11994
rect 5642 11942 5644 11994
rect 5398 11940 5404 11942
rect 5460 11940 5484 11942
rect 5540 11940 5564 11942
rect 5620 11940 5644 11942
rect 5700 11940 5706 11942
rect 5398 11931 5706 11940
rect 5920 11558 5948 13330
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5398 10908 5706 10917
rect 5398 10906 5404 10908
rect 5460 10906 5484 10908
rect 5540 10906 5564 10908
rect 5620 10906 5644 10908
rect 5700 10906 5706 10908
rect 5460 10854 5462 10906
rect 5642 10854 5644 10906
rect 5398 10852 5404 10854
rect 5460 10852 5484 10854
rect 5540 10852 5564 10854
rect 5620 10852 5644 10854
rect 5700 10852 5706 10854
rect 5398 10843 5706 10852
rect 5828 10470 5856 11086
rect 5920 10742 5948 11494
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5398 9820 5706 9829
rect 5398 9818 5404 9820
rect 5460 9818 5484 9820
rect 5540 9818 5564 9820
rect 5620 9818 5644 9820
rect 5700 9818 5706 9820
rect 5460 9766 5462 9818
rect 5642 9766 5644 9818
rect 5398 9764 5404 9766
rect 5460 9764 5484 9766
rect 5540 9764 5564 9766
rect 5620 9764 5644 9766
rect 5700 9764 5706 9766
rect 5398 9755 5706 9764
rect 5828 9518 5856 10406
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5828 8906 5856 9454
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5398 8732 5706 8741
rect 5398 8730 5404 8732
rect 5460 8730 5484 8732
rect 5540 8730 5564 8732
rect 5620 8730 5644 8732
rect 5700 8730 5706 8732
rect 5460 8678 5462 8730
rect 5642 8678 5644 8730
rect 5398 8676 5404 8678
rect 5460 8676 5484 8678
rect 5540 8676 5564 8678
rect 5620 8676 5644 8678
rect 5700 8676 5706 8678
rect 5398 8667 5706 8676
rect 5736 8616 5764 8842
rect 5644 8588 5764 8616
rect 5644 7750 5672 8588
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5398 7644 5706 7653
rect 5398 7642 5404 7644
rect 5460 7642 5484 7644
rect 5540 7642 5564 7644
rect 5620 7642 5644 7644
rect 5700 7642 5706 7644
rect 5460 7590 5462 7642
rect 5642 7590 5644 7642
rect 5398 7588 5404 7590
rect 5460 7588 5484 7590
rect 5540 7588 5564 7590
rect 5620 7588 5644 7590
rect 5700 7588 5706 7590
rect 5398 7579 5706 7588
rect 5736 7426 5764 8230
rect 5644 7410 5764 7426
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5632 7404 5764 7410
rect 5684 7398 5764 7404
rect 5632 7346 5684 7352
rect 5184 7206 5212 7346
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5078 3088 5134 3097
rect 5078 3023 5080 3032
rect 5132 3023 5134 3032
rect 5080 2994 5132 3000
rect 5184 2774 5212 7142
rect 5398 6556 5706 6565
rect 5398 6554 5404 6556
rect 5460 6554 5484 6556
rect 5540 6554 5564 6556
rect 5620 6554 5644 6556
rect 5700 6554 5706 6556
rect 5460 6502 5462 6554
rect 5642 6502 5644 6554
rect 5398 6500 5404 6502
rect 5460 6500 5484 6502
rect 5540 6500 5564 6502
rect 5620 6500 5644 6502
rect 5700 6500 5706 6502
rect 5398 6491 5706 6500
rect 5736 6338 5764 7398
rect 5828 7002 5856 8434
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5644 6322 5764 6338
rect 5920 6322 5948 9862
rect 5632 6316 5764 6322
rect 5684 6310 5764 6316
rect 5908 6316 5960 6322
rect 5632 6258 5684 6264
rect 5908 6258 5960 6264
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5398 5468 5706 5477
rect 5398 5466 5404 5468
rect 5460 5466 5484 5468
rect 5540 5466 5564 5468
rect 5620 5466 5644 5468
rect 5700 5466 5706 5468
rect 5460 5414 5462 5466
rect 5642 5414 5644 5466
rect 5398 5412 5404 5414
rect 5460 5412 5484 5414
rect 5540 5412 5564 5414
rect 5620 5412 5644 5414
rect 5700 5412 5706 5414
rect 5398 5403 5706 5412
rect 5736 5352 5764 5850
rect 5552 5324 5764 5352
rect 5552 4690 5580 5324
rect 5828 5166 5856 6054
rect 5920 5778 5948 6258
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5920 5166 5948 5714
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4690 5764 4966
rect 5828 4826 5856 5102
rect 5906 4856 5962 4865
rect 5816 4820 5868 4826
rect 5906 4791 5962 4800
rect 5816 4762 5868 4768
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5398 4380 5706 4389
rect 5398 4378 5404 4380
rect 5460 4378 5484 4380
rect 5540 4378 5564 4380
rect 5620 4378 5644 4380
rect 5700 4378 5706 4380
rect 5460 4326 5462 4378
rect 5642 4326 5644 4378
rect 5398 4324 5404 4326
rect 5460 4324 5484 4326
rect 5540 4324 5564 4326
rect 5620 4324 5644 4326
rect 5700 4324 5706 4326
rect 5398 4315 5706 4324
rect 5920 4282 5948 4791
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5398 3292 5706 3301
rect 5398 3290 5404 3292
rect 5460 3290 5484 3292
rect 5540 3290 5564 3292
rect 5620 3290 5644 3292
rect 5700 3290 5706 3292
rect 5460 3238 5462 3290
rect 5642 3238 5644 3290
rect 5398 3236 5404 3238
rect 5460 3236 5484 3238
rect 5540 3236 5564 3238
rect 5620 3236 5644 3238
rect 5700 3236 5706 3238
rect 5398 3227 5706 3236
rect 4816 2746 4936 2774
rect 4908 2446 4936 2746
rect 5092 2746 5212 2774
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5092 800 5120 2746
rect 5398 2204 5706 2213
rect 5398 2202 5404 2204
rect 5460 2202 5484 2204
rect 5540 2202 5564 2204
rect 5620 2202 5644 2204
rect 5700 2202 5706 2204
rect 5460 2150 5462 2202
rect 5642 2150 5644 2202
rect 5398 2148 5404 2150
rect 5460 2148 5484 2150
rect 5540 2148 5564 2150
rect 5620 2148 5644 2150
rect 5700 2148 5706 2150
rect 5398 2139 5706 2148
rect 5736 1850 5764 3946
rect 5552 1822 5764 1850
rect 5552 800 5580 1822
rect 6012 800 6040 13806
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 13190 6408 13670
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6380 12986 6408 13126
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6288 12434 6316 12854
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6196 12406 6316 12434
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6104 11830 6132 12038
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 6196 11150 6224 12406
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6288 11558 6316 11630
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6380 11354 6408 12718
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6472 11665 6500 11834
rect 6458 11656 6514 11665
rect 6458 11591 6514 11600
rect 6472 11558 6500 11591
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6104 8838 6132 9318
rect 6196 9178 6224 9318
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6104 8362 6132 8774
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 5710 6132 7686
rect 6288 6934 6316 11018
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 6196 5914 6224 6666
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6288 5574 6316 5782
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6196 5302 6224 5510
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6104 4486 6132 5102
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6380 2854 6408 11154
rect 6472 7698 6500 11494
rect 6564 10266 6592 12242
rect 6656 11898 6684 12786
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6564 9654 6592 10202
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6472 7670 6684 7698
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6472 800 6500 7414
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6564 6254 6592 6394
rect 6552 6248 6604 6254
rect 6550 6216 6552 6225
rect 6604 6216 6606 6225
rect 6550 6151 6606 6160
rect 6564 5370 6592 6151
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6564 4282 6592 5306
rect 6656 5166 6684 7670
rect 6748 7478 6776 14010
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6840 12782 6868 13398
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 7024 12714 7052 13194
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7208 12986 7236 13126
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7116 11898 7144 12650
rect 7208 12102 7236 12786
rect 7288 12436 7340 12442
rect 7392 12434 7420 16400
rect 7622 14716 7930 14725
rect 7622 14714 7628 14716
rect 7684 14714 7708 14716
rect 7764 14714 7788 14716
rect 7844 14714 7868 14716
rect 7924 14714 7930 14716
rect 7684 14662 7686 14714
rect 7866 14662 7868 14714
rect 7622 14660 7628 14662
rect 7684 14660 7708 14662
rect 7764 14660 7788 14662
rect 7844 14660 7868 14662
rect 7924 14660 7930 14662
rect 7622 14651 7930 14660
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7760 14074 7788 14418
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7760 13938 7788 14010
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7622 13628 7930 13637
rect 7622 13626 7628 13628
rect 7684 13626 7708 13628
rect 7764 13626 7788 13628
rect 7844 13626 7868 13628
rect 7924 13626 7930 13628
rect 7684 13574 7686 13626
rect 7866 13574 7868 13626
rect 7622 13572 7628 13574
rect 7684 13572 7708 13574
rect 7764 13572 7788 13574
rect 7844 13572 7868 13574
rect 7924 13572 7930 13574
rect 7622 13563 7930 13572
rect 7622 12540 7930 12549
rect 7622 12538 7628 12540
rect 7684 12538 7708 12540
rect 7764 12538 7788 12540
rect 7844 12538 7868 12540
rect 7924 12538 7930 12540
rect 7684 12486 7686 12538
rect 7866 12486 7868 12538
rect 7622 12484 7628 12486
rect 7684 12484 7708 12486
rect 7764 12484 7788 12486
rect 7844 12484 7868 12486
rect 7924 12484 7930 12486
rect 7622 12475 7930 12484
rect 7392 12406 7512 12434
rect 7288 12378 7340 12384
rect 7300 12238 7328 12378
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 6920 11756 6972 11762
rect 6840 11716 6920 11744
rect 6840 11354 6868 11716
rect 6920 11698 6972 11704
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6932 10810 6960 11494
rect 7012 11280 7064 11286
rect 7208 11268 7236 12038
rect 7300 11694 7328 12174
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7012 11222 7064 11228
rect 7116 11240 7236 11268
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6840 10470 6868 10678
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6840 9518 6868 9998
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 8974 6868 9454
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6840 8566 6868 8910
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6748 6186 6776 6394
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6840 5370 6868 6734
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 4690 6776 4966
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6840 4486 6868 5306
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6656 4214 6684 4422
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6932 3534 6960 4966
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 7024 3058 7052 11222
rect 7116 9586 7144 11240
rect 7300 11218 7328 11630
rect 7392 11626 7420 12242
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7392 9994 7420 11562
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7116 6662 7144 8842
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 5302 7144 6598
rect 7104 5296 7156 5302
rect 7104 5238 7156 5244
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7116 4826 7144 5102
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7300 3602 7328 9522
rect 7392 9178 7420 9930
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7484 7936 7512 12406
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7576 11558 7604 12174
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7622 11452 7930 11461
rect 7622 11450 7628 11452
rect 7684 11450 7708 11452
rect 7764 11450 7788 11452
rect 7844 11450 7868 11452
rect 7924 11450 7930 11452
rect 7684 11398 7686 11450
rect 7866 11398 7868 11450
rect 7622 11396 7628 11398
rect 7684 11396 7708 11398
rect 7764 11396 7788 11398
rect 7844 11396 7868 11398
rect 7924 11396 7930 11398
rect 7622 11387 7930 11396
rect 7622 10364 7930 10373
rect 7622 10362 7628 10364
rect 7684 10362 7708 10364
rect 7764 10362 7788 10364
rect 7844 10362 7868 10364
rect 7924 10362 7930 10364
rect 7684 10310 7686 10362
rect 7866 10310 7868 10362
rect 7622 10308 7628 10310
rect 7684 10308 7708 10310
rect 7764 10308 7788 10310
rect 7844 10308 7868 10310
rect 7924 10308 7930 10310
rect 7622 10299 7930 10308
rect 8036 9586 8064 16400
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8588 14074 8616 14350
rect 8864 14074 8892 14826
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8864 13977 8892 14010
rect 8850 13968 8906 13977
rect 8850 13903 8852 13912
rect 8904 13903 8906 13912
rect 8852 13874 8904 13880
rect 8864 13843 8892 13874
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8220 12782 8248 13330
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8128 9466 8156 12038
rect 8220 11234 8248 12718
rect 8312 11898 8340 13126
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8220 11218 8340 11234
rect 8220 11212 8352 11218
rect 8220 11206 8300 11212
rect 8220 10674 8248 11206
rect 8300 11154 8352 11160
rect 8404 10742 8432 11562
rect 8588 11257 8616 11698
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8574 11248 8630 11257
rect 8574 11183 8576 11192
rect 8628 11183 8630 11192
rect 8576 11154 8628 11160
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8220 10266 8248 10610
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8404 10198 8432 10678
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8128 9438 8248 9466
rect 7622 9276 7930 9285
rect 7622 9274 7628 9276
rect 7684 9274 7708 9276
rect 7764 9274 7788 9276
rect 7844 9274 7868 9276
rect 7924 9274 7930 9276
rect 7684 9222 7686 9274
rect 7866 9222 7868 9274
rect 7622 9220 7628 9222
rect 7684 9220 7708 9222
rect 7764 9220 7788 9222
rect 7844 9220 7868 9222
rect 7924 9220 7930 9222
rect 7622 9211 7930 9220
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7576 9081 7604 9114
rect 7562 9072 7618 9081
rect 7562 9007 7618 9016
rect 7622 8188 7930 8197
rect 7622 8186 7628 8188
rect 7684 8186 7708 8188
rect 7764 8186 7788 8188
rect 7844 8186 7868 8188
rect 7924 8186 7930 8188
rect 7684 8134 7686 8186
rect 7866 8134 7868 8186
rect 7622 8132 7628 8134
rect 7684 8132 7708 8134
rect 7764 8132 7788 8134
rect 7844 8132 7868 8134
rect 7924 8132 7930 8134
rect 7622 8123 7930 8132
rect 7392 7908 7512 7936
rect 7392 5846 7420 7908
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 7484 7206 7512 7754
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7484 5710 7512 7142
rect 7622 7100 7930 7109
rect 7622 7098 7628 7100
rect 7684 7098 7708 7100
rect 7764 7098 7788 7100
rect 7844 7098 7868 7100
rect 7924 7098 7930 7100
rect 7684 7046 7686 7098
rect 7866 7046 7868 7098
rect 7622 7044 7628 7046
rect 7684 7044 7708 7046
rect 7764 7044 7788 7046
rect 7844 7044 7868 7046
rect 7924 7044 7930 7046
rect 7622 7035 7930 7044
rect 8036 6118 8064 7346
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7622 6012 7930 6021
rect 7622 6010 7628 6012
rect 7684 6010 7708 6012
rect 7764 6010 7788 6012
rect 7844 6010 7868 6012
rect 7924 6010 7930 6012
rect 7684 5958 7686 6010
rect 7866 5958 7868 6010
rect 7622 5956 7628 5958
rect 7684 5956 7708 5958
rect 7764 5956 7788 5958
rect 7844 5956 7868 5958
rect 7924 5956 7930 5958
rect 7622 5947 7930 5956
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7392 3058 7420 5510
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 4729 7512 5170
rect 7622 4924 7930 4933
rect 7622 4922 7628 4924
rect 7684 4922 7708 4924
rect 7764 4922 7788 4924
rect 7844 4922 7868 4924
rect 7924 4922 7930 4924
rect 7684 4870 7686 4922
rect 7866 4870 7868 4922
rect 7622 4868 7628 4870
rect 7684 4868 7708 4870
rect 7764 4868 7788 4870
rect 7844 4868 7868 4870
rect 7924 4868 7930 4870
rect 7622 4859 7930 4868
rect 7470 4720 7526 4729
rect 8036 4690 8064 6054
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8128 5234 8156 5782
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7470 4655 7472 4664
rect 7524 4655 7526 4664
rect 8024 4684 8076 4690
rect 7472 4626 7524 4632
rect 8024 4626 8076 4632
rect 8128 4554 8156 5170
rect 8220 4570 8248 9438
rect 8588 8294 8616 11154
rect 8680 11082 8708 11630
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8680 8838 8708 9522
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8312 7342 8340 7822
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8312 6746 8340 7278
rect 8392 6792 8444 6798
rect 8312 6740 8392 6746
rect 8312 6734 8444 6740
rect 8312 6718 8432 6734
rect 8312 6390 8340 6718
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8496 5234 8524 7686
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8116 4548 8168 4554
rect 8220 4542 8340 4570
rect 8116 4490 8168 4496
rect 8128 4282 8156 4490
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8220 4282 8248 4422
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8312 4162 8340 4542
rect 8220 4134 8340 4162
rect 8864 4146 8892 6054
rect 8852 4140 8904 4146
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 7622 3836 7930 3845
rect 7622 3834 7628 3836
rect 7684 3834 7708 3836
rect 7764 3834 7788 3836
rect 7844 3834 7868 3836
rect 7924 3834 7930 3836
rect 7684 3782 7686 3834
rect 7866 3782 7868 3834
rect 7622 3780 7628 3782
rect 7684 3780 7708 3782
rect 7764 3780 7788 3782
rect 7844 3780 7868 3782
rect 7924 3780 7930 3782
rect 7622 3771 7930 3780
rect 8128 3466 8156 4014
rect 8220 3738 8248 4134
rect 8852 4082 8904 4088
rect 8758 4040 8814 4049
rect 8758 3975 8814 3984
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7576 3126 7604 3334
rect 8128 3194 8156 3402
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 7564 3120 7616 3126
rect 7564 3062 7616 3068
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7392 2961 7420 2994
rect 7378 2952 7434 2961
rect 7378 2887 7434 2896
rect 8680 2854 8708 3130
rect 8772 3126 8800 3975
rect 8956 3738 8984 16510
rect 9048 16510 9366 16538
rect 9048 4078 9076 16510
rect 9310 16400 9366 16510
rect 9954 16538 10010 17200
rect 10598 16538 10654 17200
rect 11242 16538 11298 17200
rect 9954 16510 10272 16538
rect 9954 16400 10010 16510
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9140 14074 9168 14350
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9784 14074 9812 14282
rect 9846 14172 10154 14181
rect 9846 14170 9852 14172
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 10148 14170 10154 14172
rect 9908 14118 9910 14170
rect 10090 14118 10092 14170
rect 9846 14116 9852 14118
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 10148 14116 10154 14118
rect 9846 14107 10154 14116
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9140 13841 9168 14010
rect 9126 13832 9182 13841
rect 9126 13767 9182 13776
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9416 12170 9444 13330
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9508 12442 9536 12718
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9600 12306 9628 13126
rect 9846 13084 10154 13093
rect 9846 13082 9852 13084
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 10148 13082 10154 13084
rect 9908 13030 9910 13082
rect 10090 13030 10092 13082
rect 9846 13028 9852 13030
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 10148 13028 10154 13030
rect 9846 13019 10154 13028
rect 10244 12986 10272 16510
rect 10336 16510 10654 16538
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9692 12442 9720 12786
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9770 12336 9826 12345
rect 9588 12300 9640 12306
rect 10244 12306 10272 12718
rect 9770 12271 9826 12280
rect 10232 12300 10284 12306
rect 9588 12242 9640 12248
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9416 11694 9444 12106
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9784 11626 9812 12271
rect 10232 12242 10284 12248
rect 9846 11996 10154 12005
rect 9846 11994 9852 11996
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 10148 11994 10154 11996
rect 9908 11942 9910 11994
rect 10090 11942 10092 11994
rect 9846 11940 9852 11942
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 10148 11940 10154 11942
rect 9846 11931 10154 11940
rect 10244 11694 10272 12242
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9324 11150 9352 11494
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9416 10810 9444 11290
rect 9508 11286 9536 11494
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9600 11218 9628 11290
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9692 11098 9720 11494
rect 9784 11354 9812 11562
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9600 11082 9720 11098
rect 10060 11082 10088 11630
rect 9588 11076 9720 11082
rect 9640 11070 9720 11076
rect 10048 11076 10100 11082
rect 9588 11018 9640 11024
rect 10048 11018 10100 11024
rect 9846 10908 10154 10917
rect 9846 10906 9852 10908
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 10148 10906 10154 10908
rect 9908 10854 9910 10906
rect 10090 10854 10092 10906
rect 9846 10852 9852 10854
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 10148 10852 10154 10854
rect 9846 10843 10154 10852
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9416 8566 9444 10746
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9588 9648 9640 9654
rect 9692 9636 9720 10542
rect 10140 10056 10192 10062
rect 10244 10044 10272 11630
rect 10192 10016 10272 10044
rect 10140 9998 10192 10004
rect 9846 9820 10154 9829
rect 9846 9818 9852 9820
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 10148 9818 10154 9820
rect 9908 9766 9910 9818
rect 10090 9766 10092 9818
rect 9846 9764 9852 9766
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 10148 9764 10154 9766
rect 9846 9755 10154 9764
rect 9640 9608 9720 9636
rect 9588 9590 9640 9596
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9692 9178 9720 9386
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9784 8974 9812 9318
rect 10244 9178 10272 10016
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9784 8634 9812 8910
rect 9846 8732 10154 8741
rect 9846 8730 9852 8732
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 10148 8730 10154 8732
rect 9908 8678 9910 8730
rect 10090 8678 10092 8730
rect 9846 8676 9852 8678
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 10148 8676 10154 8678
rect 9846 8667 10154 8676
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7410 9352 7686
rect 9846 7644 10154 7653
rect 9846 7642 9852 7644
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 10148 7642 10154 7644
rect 9908 7590 9910 7642
rect 10090 7590 10092 7642
rect 9846 7588 9852 7590
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 10148 7588 10154 7590
rect 9846 7579 10154 7588
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9324 5710 9352 7346
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 9416 6798 9444 7142
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9232 4622 9260 5510
rect 9416 5234 9444 6734
rect 9846 6556 10154 6565
rect 9846 6554 9852 6556
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 10148 6554 10154 6556
rect 9908 6502 9910 6554
rect 10090 6502 10092 6554
rect 9846 6500 9852 6502
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 10148 6500 10154 6502
rect 9846 6491 10154 6500
rect 10244 6338 10272 7142
rect 10152 6322 10272 6338
rect 10140 6316 10272 6322
rect 10192 6310 10272 6316
rect 10140 6258 10192 6264
rect 9846 5468 10154 5477
rect 9846 5466 9852 5468
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 10148 5466 10154 5468
rect 9908 5414 9910 5466
rect 10090 5414 10092 5466
rect 9846 5412 9852 5414
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 10148 5412 10154 5414
rect 9846 5403 10154 5412
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4214 9168 4422
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9048 3738 9076 4014
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9140 3534 9168 4150
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 6932 800 6960 2790
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7392 800 7420 2246
rect 3344 734 3648 762
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6918 0 6974 800
rect 7378 0 7434 800
rect 7484 762 7512 2790
rect 7622 2748 7930 2757
rect 7622 2746 7628 2748
rect 7684 2746 7708 2748
rect 7764 2746 7788 2748
rect 7844 2746 7868 2748
rect 7924 2746 7930 2748
rect 7684 2694 7686 2746
rect 7866 2694 7868 2746
rect 7622 2692 7628 2694
rect 7684 2692 7708 2694
rect 7764 2692 7788 2694
rect 7844 2692 7868 2694
rect 7924 2692 7930 2694
rect 7622 2683 7930 2692
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 7760 870 7880 898
rect 7760 762 7788 870
rect 7852 800 7880 870
rect 8312 800 8340 2246
rect 8772 800 8800 2790
rect 9140 2446 9168 3470
rect 9232 3058 9260 4558
rect 9600 4214 9628 5102
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9310 4040 9366 4049
rect 9310 3975 9366 3984
rect 9324 3126 9352 3975
rect 9600 3534 9628 4150
rect 9692 4049 9720 5102
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9784 4690 9812 5034
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 9846 4380 10154 4389
rect 9846 4378 9852 4380
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 10148 4378 10154 4380
rect 9908 4326 9910 4378
rect 10090 4326 10092 4378
rect 9846 4324 9852 4326
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 10148 4324 10154 4326
rect 9846 4315 10154 4324
rect 10048 4072 10100 4078
rect 9678 4040 9734 4049
rect 10048 4014 10100 4020
rect 9678 3975 9734 3984
rect 9588 3528 9640 3534
rect 9508 3488 9588 3516
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9416 2378 9444 2926
rect 9508 2446 9536 3488
rect 9588 3470 9640 3476
rect 9692 2666 9720 3975
rect 10060 3670 10088 4014
rect 10244 3942 10272 4558
rect 10336 4078 10364 16510
rect 10598 16400 10654 16510
rect 11072 16510 11298 16538
rect 10506 12744 10562 12753
rect 10506 12679 10508 12688
rect 10560 12679 10562 12688
rect 10508 12650 10560 12656
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10428 11898 10456 12174
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10428 11506 10456 11698
rect 10520 11626 10548 12038
rect 10508 11620 10560 11626
rect 10508 11562 10560 11568
rect 10428 11478 10548 11506
rect 10520 11121 10548 11478
rect 10506 11112 10562 11121
rect 10506 11047 10562 11056
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10428 9654 10456 9998
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10428 7818 10456 8230
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 5234 10456 6598
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 10520 3505 10548 11047
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10612 7410 10640 7822
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 4690 10824 6598
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10796 4010 10824 4490
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10506 3496 10562 3505
rect 10506 3431 10562 3440
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9784 3126 9812 3334
rect 9846 3292 10154 3301
rect 9846 3290 9852 3292
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 10148 3290 10154 3292
rect 9908 3238 9910 3290
rect 10090 3238 10092 3290
rect 9846 3236 9852 3238
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 10148 3236 10154 3238
rect 9846 3227 10154 3236
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 10796 3058 10824 3946
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10232 2916 10284 2922
rect 10232 2858 10284 2864
rect 9692 2638 9812 2666
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9232 870 9352 898
rect 9232 800 9260 870
rect 7484 734 7788 762
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9324 762 9352 870
rect 9508 762 9536 2246
rect 9692 800 9720 2518
rect 9784 2446 9812 2638
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9846 2204 10154 2213
rect 9846 2202 9852 2204
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 10148 2202 10154 2204
rect 9908 2150 9910 2202
rect 10090 2150 10092 2202
rect 9846 2148 9852 2150
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 10148 2148 10154 2150
rect 9846 2139 10154 2148
rect 10244 1442 10272 2858
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10152 1414 10272 1442
rect 10152 800 10180 1414
rect 10612 800 10640 2790
rect 10888 2582 10916 12038
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10980 10538 11008 11018
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 11072 5352 11100 16510
rect 11242 16400 11298 16510
rect 11886 16400 11942 17200
rect 12530 16400 12586 17200
rect 13174 16538 13230 17200
rect 12728 16510 13230 16538
rect 11704 15224 11756 15230
rect 11704 15166 11756 15172
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11256 14550 11284 14894
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 11164 14074 11192 14486
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11624 13530 11652 13670
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11152 13184 11204 13190
rect 11336 13184 11388 13190
rect 11204 13144 11284 13172
rect 11152 13126 11204 13132
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11164 5370 11192 12922
rect 11256 12238 11284 13144
rect 11336 13126 11388 13132
rect 11348 12986 11376 13126
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11716 12442 11744 15166
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11348 9178 11376 11018
rect 11532 10062 11560 11086
rect 11624 10470 11652 12242
rect 11716 10810 11744 12242
rect 11808 11558 11836 12582
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11716 10674 11744 10746
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11532 9654 11560 9998
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11532 9042 11560 9590
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11532 8498 11560 8978
rect 11624 8498 11652 10406
rect 11900 9466 11928 16400
rect 12070 14716 12378 14725
rect 12070 14714 12076 14716
rect 12132 14714 12156 14716
rect 12212 14714 12236 14716
rect 12292 14714 12316 14716
rect 12372 14714 12378 14716
rect 12132 14662 12134 14714
rect 12314 14662 12316 14714
rect 12070 14660 12076 14662
rect 12132 14660 12156 14662
rect 12212 14660 12236 14662
rect 12292 14660 12316 14662
rect 12372 14660 12378 14662
rect 12070 14651 12378 14660
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12452 14006 12480 14282
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12070 13628 12378 13637
rect 12070 13626 12076 13628
rect 12132 13626 12156 13628
rect 12212 13626 12236 13628
rect 12292 13626 12316 13628
rect 12372 13626 12378 13628
rect 12132 13574 12134 13626
rect 12314 13574 12316 13626
rect 12070 13572 12076 13574
rect 12132 13572 12156 13574
rect 12212 13572 12236 13574
rect 12292 13572 12316 13574
rect 12372 13572 12378 13574
rect 12070 13563 12378 13572
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11992 12306 12020 13330
rect 12176 13326 12204 13466
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12084 12918 12112 13262
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12176 12714 12204 13262
rect 12452 12782 12480 13330
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 12070 12540 12378 12549
rect 12070 12538 12076 12540
rect 12132 12538 12156 12540
rect 12212 12538 12236 12540
rect 12292 12538 12316 12540
rect 12372 12538 12378 12540
rect 12132 12486 12134 12538
rect 12314 12486 12316 12538
rect 12070 12484 12076 12486
rect 12132 12484 12156 12486
rect 12212 12484 12236 12486
rect 12292 12484 12316 12486
rect 12372 12484 12378 12486
rect 12070 12475 12378 12484
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 12452 11898 12480 12378
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12070 11452 12378 11461
rect 12070 11450 12076 11452
rect 12132 11450 12156 11452
rect 12212 11450 12236 11452
rect 12292 11450 12316 11452
rect 12372 11450 12378 11452
rect 12132 11398 12134 11450
rect 12314 11398 12316 11450
rect 12070 11396 12076 11398
rect 12132 11396 12156 11398
rect 12212 11396 12236 11398
rect 12292 11396 12316 11398
rect 12372 11396 12378 11398
rect 12070 11387 12378 11396
rect 12070 10364 12378 10373
rect 12070 10362 12076 10364
rect 12132 10362 12156 10364
rect 12212 10362 12236 10364
rect 12292 10362 12316 10364
rect 12372 10362 12378 10364
rect 12132 10310 12134 10362
rect 12314 10310 12316 10362
rect 12070 10308 12076 10310
rect 12132 10308 12156 10310
rect 12212 10308 12236 10310
rect 12292 10308 12316 10310
rect 12372 10308 12378 10310
rect 12070 10299 12378 10308
rect 11716 9438 11928 9466
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 10980 5324 11100 5352
rect 11152 5364 11204 5370
rect 10980 4690 11008 5324
rect 11152 5306 11204 5312
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 11072 4554 11100 5170
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11072 2582 11100 4218
rect 11164 2961 11192 4422
rect 11256 3534 11284 5578
rect 11348 5030 11376 6734
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11716 4214 11744 9438
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 7478 11928 9318
rect 12070 9276 12378 9285
rect 12070 9274 12076 9276
rect 12132 9274 12156 9276
rect 12212 9274 12236 9276
rect 12292 9274 12316 9276
rect 12372 9274 12378 9276
rect 12132 9222 12134 9274
rect 12314 9222 12316 9274
rect 12070 9220 12076 9222
rect 12132 9220 12156 9222
rect 12212 9220 12236 9222
rect 12292 9220 12316 9222
rect 12372 9220 12378 9222
rect 12070 9211 12378 9220
rect 12070 8188 12378 8197
rect 12070 8186 12076 8188
rect 12132 8186 12156 8188
rect 12212 8186 12236 8188
rect 12292 8186 12316 8188
rect 12372 8186 12378 8188
rect 12132 8134 12134 8186
rect 12314 8134 12316 8186
rect 12070 8132 12076 8134
rect 12132 8132 12156 8134
rect 12212 8132 12236 8134
rect 12292 8132 12316 8134
rect 12372 8132 12378 8134
rect 12070 8123 12378 8132
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11992 7002 12020 7346
rect 12268 7290 12296 7686
rect 12268 7262 12480 7290
rect 12070 7100 12378 7109
rect 12070 7098 12076 7100
rect 12132 7098 12156 7100
rect 12212 7098 12236 7100
rect 12292 7098 12316 7100
rect 12372 7098 12378 7100
rect 12132 7046 12134 7098
rect 12314 7046 12316 7098
rect 12070 7044 12076 7046
rect 12132 7044 12156 7046
rect 12212 7044 12236 7046
rect 12292 7044 12316 7046
rect 12372 7044 12378 7046
rect 12070 7035 12378 7044
rect 11980 6996 12032 7002
rect 12452 6984 12480 7262
rect 11980 6938 12032 6944
rect 12360 6956 12480 6984
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 11992 5710 12020 6666
rect 12360 6390 12388 6956
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12070 6012 12378 6021
rect 12070 6010 12076 6012
rect 12132 6010 12156 6012
rect 12212 6010 12236 6012
rect 12292 6010 12316 6012
rect 12372 6010 12378 6012
rect 12132 5958 12134 6010
rect 12314 5958 12316 6010
rect 12070 5956 12076 5958
rect 12132 5956 12156 5958
rect 12212 5956 12236 5958
rect 12292 5956 12316 5958
rect 12372 5956 12378 5958
rect 12070 5947 12378 5956
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11808 4486 11836 5238
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11900 4622 11928 5102
rect 12070 4924 12378 4933
rect 12070 4922 12076 4924
rect 12132 4922 12156 4924
rect 12212 4922 12236 4924
rect 12292 4922 12316 4924
rect 12372 4922 12378 4924
rect 12132 4870 12134 4922
rect 12314 4870 12316 4922
rect 12070 4868 12076 4870
rect 12132 4868 12156 4870
rect 12212 4868 12236 4870
rect 12292 4868 12316 4870
rect 12372 4868 12378 4870
rect 12070 4859 12378 4868
rect 12544 4690 12572 16400
rect 12622 14376 12678 14385
rect 12622 14311 12678 14320
rect 12636 14074 12664 14311
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12636 12986 12664 13126
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 12306 12664 12582
rect 12728 12374 12756 16510
rect 13174 16400 13230 16510
rect 13818 16400 13874 17200
rect 14462 16538 14518 17200
rect 14016 16510 14518 16538
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12636 10674 12664 11630
rect 12728 11286 12756 12038
rect 12912 11898 12940 12106
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12820 11665 12848 11698
rect 12806 11656 12862 11665
rect 12806 11591 12862 11600
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12636 9178 12664 10610
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12912 10062 12940 10542
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 13004 7562 13032 14282
rect 13372 14074 13400 14758
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13096 12238 13124 12582
rect 13084 12232 13136 12238
rect 13188 12209 13216 13806
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13280 12918 13308 13330
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13372 12306 13400 12718
rect 13648 12434 13676 14554
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13740 14074 13768 14214
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13832 13705 13860 16400
rect 14016 14006 14044 16510
rect 14462 16400 14518 16510
rect 15106 16400 15162 17200
rect 15474 16552 15530 16561
rect 15474 16487 15530 16496
rect 14294 14172 14602 14181
rect 14294 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14516 14170 14540 14172
rect 14596 14170 14602 14172
rect 14356 14118 14358 14170
rect 14538 14118 14540 14170
rect 14294 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14516 14116 14540 14118
rect 14596 14116 14602 14118
rect 14294 14107 14602 14116
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13818 13696 13874 13705
rect 13818 13631 13874 13640
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12918 13860 13126
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13648 12406 13768 12434
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13084 12174 13136 12180
rect 13174 12200 13230 12209
rect 13174 12135 13230 12144
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 13096 9994 13124 11222
rect 13188 10146 13216 12135
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13280 11898 13308 12038
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13372 10742 13400 12242
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13556 11830 13584 12174
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13188 10118 13400 10146
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13280 8974 13308 9454
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 12912 7534 13032 7562
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 12636 5370 12664 5578
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 11716 4078 11744 4150
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11900 3618 11928 4558
rect 12084 4078 12112 4626
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12072 4072 12124 4078
rect 12544 4049 12572 4150
rect 12072 4014 12124 4020
rect 12530 4040 12586 4049
rect 12530 3975 12586 3984
rect 12070 3836 12378 3845
rect 12070 3834 12076 3836
rect 12132 3834 12156 3836
rect 12212 3834 12236 3836
rect 12292 3834 12316 3836
rect 12372 3834 12378 3836
rect 12132 3782 12134 3834
rect 12314 3782 12316 3834
rect 12070 3780 12076 3782
rect 12132 3780 12156 3782
rect 12212 3780 12236 3782
rect 12292 3780 12316 3782
rect 12372 3780 12378 3782
rect 12070 3771 12378 3780
rect 11900 3590 12112 3618
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11256 3126 11284 3470
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 11624 2990 11652 3402
rect 11900 3194 11928 3470
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11612 2984 11664 2990
rect 11150 2952 11206 2961
rect 11612 2926 11664 2932
rect 11150 2887 11206 2896
rect 11520 2916 11572 2922
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11164 2446 11192 2887
rect 11520 2858 11572 2864
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11072 800 11100 2246
rect 11532 800 11560 2858
rect 11716 2650 11744 3062
rect 11808 2922 11836 3130
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 11794 2816 11850 2825
rect 11794 2751 11850 2760
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11808 2530 11836 2751
rect 11716 2514 11836 2530
rect 11704 2508 11836 2514
rect 11756 2502 11836 2508
rect 11704 2450 11756 2456
rect 11900 2122 11928 2926
rect 11992 2378 12020 3334
rect 12084 3126 12112 3590
rect 12544 3534 12572 3975
rect 12622 3632 12678 3641
rect 12622 3567 12678 3576
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12636 3126 12664 3567
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12084 2961 12112 3062
rect 12070 2952 12126 2961
rect 12070 2887 12126 2896
rect 12070 2748 12378 2757
rect 12070 2746 12076 2748
rect 12132 2746 12156 2748
rect 12212 2746 12236 2748
rect 12292 2746 12316 2748
rect 12372 2746 12378 2748
rect 12132 2694 12134 2746
rect 12314 2694 12316 2746
rect 12070 2692 12076 2694
rect 12132 2692 12156 2694
rect 12212 2692 12236 2694
rect 12292 2692 12316 2694
rect 12372 2692 12378 2694
rect 12070 2683 12378 2692
rect 12820 2394 12848 5714
rect 12912 2514 12940 7534
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13096 6458 13124 6598
rect 13280 6458 13308 7754
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 13004 5846 13032 6054
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13004 2514 13032 3538
rect 13096 2922 13124 6122
rect 13188 5846 13216 6258
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 13372 5642 13400 10118
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 13464 7750 13492 8842
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 6254 13492 7686
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13542 5264 13598 5273
rect 13542 5199 13598 5208
rect 13556 5030 13584 5199
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13542 4856 13598 4865
rect 13648 4826 13676 12310
rect 13740 5370 13768 12406
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 10713 13860 11494
rect 13818 10704 13874 10713
rect 13818 10639 13874 10648
rect 13832 9518 13860 10639
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13740 5273 13768 5306
rect 13726 5264 13782 5273
rect 13726 5199 13782 5208
rect 13542 4791 13544 4800
rect 13596 4791 13598 4800
rect 13636 4820 13688 4826
rect 13544 4762 13596 4768
rect 13636 4762 13688 4768
rect 13740 4486 13768 5199
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13372 3398 13400 3538
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13084 2916 13136 2922
rect 13084 2858 13136 2864
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 11980 2372 12032 2378
rect 12820 2366 12940 2394
rect 11980 2314 12032 2320
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 11900 2094 12020 2122
rect 11992 800 12020 2094
rect 12452 800 12480 2246
rect 12912 800 12940 2366
rect 13372 800 13400 3334
rect 13464 3194 13492 4014
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13832 3097 13860 7142
rect 13818 3088 13874 3097
rect 13818 3023 13874 3032
rect 13924 2922 13952 13874
rect 14016 2990 14044 13942
rect 14108 13870 14136 14010
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14294 13084 14602 13093
rect 14294 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14516 13082 14540 13084
rect 14596 13082 14602 13084
rect 14356 13030 14358 13082
rect 14538 13030 14540 13082
rect 14294 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14516 13028 14540 13030
rect 14596 13028 14602 13030
rect 14294 13019 14602 13028
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14108 12442 14136 12786
rect 14292 12753 14320 12786
rect 14464 12776 14516 12782
rect 14278 12744 14334 12753
rect 14464 12718 14516 12724
rect 14278 12679 14334 12688
rect 14292 12646 14320 12679
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14096 12436 14148 12442
rect 14476 12434 14504 12718
rect 14476 12406 14688 12434
rect 14096 12378 14148 12384
rect 14660 12306 14688 12406
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14108 11626 14136 12038
rect 14294 11996 14602 12005
rect 14294 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14516 11994 14540 11996
rect 14596 11994 14602 11996
rect 14356 11942 14358 11994
rect 14538 11942 14540 11994
rect 14294 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14516 11940 14540 11942
rect 14596 11940 14602 11942
rect 14294 11931 14602 11940
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 14200 9926 14228 11698
rect 14660 11694 14688 12242
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14832 11620 14884 11626
rect 14832 11562 14884 11568
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14294 10908 14602 10917
rect 14294 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14516 10906 14540 10908
rect 14596 10906 14602 10908
rect 14356 10854 14358 10906
rect 14538 10854 14540 10906
rect 14294 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14516 10852 14540 10854
rect 14596 10852 14602 10854
rect 14294 10843 14602 10852
rect 14660 10810 14688 11018
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14464 10600 14516 10606
rect 14462 10568 14464 10577
rect 14516 10568 14518 10577
rect 14462 10503 14518 10512
rect 14752 10266 14780 11154
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14294 9820 14602 9829
rect 14294 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14516 9818 14540 9820
rect 14596 9818 14602 9820
rect 14356 9766 14358 9818
rect 14538 9766 14540 9818
rect 14294 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14516 9764 14540 9766
rect 14596 9764 14602 9766
rect 14294 9755 14602 9764
rect 14844 9654 14872 11562
rect 14936 11200 14964 14010
rect 15120 13938 15148 16400
rect 15290 15736 15346 15745
rect 15290 15671 15346 15680
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13433 15056 13670
rect 15014 13424 15070 13433
rect 15304 13394 15332 15671
rect 15488 15230 15516 16487
rect 15750 16400 15806 17200
rect 16394 16400 16450 17200
rect 17038 16400 17094 17200
rect 17682 16538 17738 17200
rect 17328 16510 17738 16538
rect 15476 15224 15528 15230
rect 15476 15166 15528 15172
rect 15764 13938 15792 16400
rect 16210 16144 16266 16153
rect 16210 16079 16266 16088
rect 16026 14920 16082 14929
rect 16026 14855 16082 14864
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 15856 14113 15884 14486
rect 15842 14104 15898 14113
rect 15842 14039 15898 14048
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15014 13359 15070 13368
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15200 13320 15252 13326
rect 15198 13288 15200 13297
rect 15252 13288 15254 13297
rect 15198 13223 15254 13232
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15212 11898 15240 12242
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15120 11558 15148 11698
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15290 11248 15346 11257
rect 14936 11172 15148 11200
rect 15396 11218 15424 11494
rect 15290 11183 15346 11192
rect 15384 11212 15436 11218
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14832 9648 14884 9654
rect 14832 9590 14884 9596
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14660 8838 14688 9318
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14752 8974 14780 9114
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14294 8732 14602 8741
rect 14294 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14516 8730 14540 8732
rect 14596 8730 14602 8732
rect 14356 8678 14358 8730
rect 14538 8678 14540 8730
rect 14294 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14516 8676 14540 8678
rect 14596 8676 14602 8678
rect 14294 8667 14602 8676
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14568 7750 14596 8366
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14294 7644 14602 7653
rect 14294 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14516 7642 14540 7644
rect 14596 7642 14602 7644
rect 14356 7590 14358 7642
rect 14538 7590 14540 7642
rect 14294 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14516 7588 14540 7590
rect 14596 7588 14602 7590
rect 14294 7579 14602 7588
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 5137 14136 6598
rect 14200 5914 14228 7482
rect 14294 6556 14602 6565
rect 14294 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14516 6554 14540 6556
rect 14596 6554 14602 6556
rect 14356 6502 14358 6554
rect 14538 6502 14540 6554
rect 14294 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14516 6500 14540 6502
rect 14596 6500 14602 6502
rect 14294 6491 14602 6500
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14200 5710 14228 5850
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14294 5468 14602 5477
rect 14294 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14516 5466 14540 5468
rect 14596 5466 14602 5468
rect 14356 5414 14358 5466
rect 14538 5414 14540 5466
rect 14294 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14516 5412 14540 5414
rect 14596 5412 14602 5414
rect 14294 5403 14602 5412
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14384 5250 14412 5306
rect 14384 5222 14504 5250
rect 14188 5160 14240 5166
rect 14094 5128 14150 5137
rect 14188 5102 14240 5108
rect 14094 5063 14150 5072
rect 14096 4752 14148 4758
rect 14200 4740 14228 5102
rect 14476 4826 14504 5222
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14148 4712 14228 4740
rect 14096 4694 14148 4700
rect 14292 4622 14320 4762
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14294 4380 14602 4389
rect 14294 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14516 4378 14540 4380
rect 14596 4378 14602 4380
rect 14356 4326 14358 4378
rect 14538 4326 14540 4378
rect 14294 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14516 4324 14540 4326
rect 14596 4324 14602 4326
rect 14294 4315 14602 4324
rect 14660 4282 14688 8774
rect 14752 8430 14780 8910
rect 14844 8634 14872 9590
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14752 8090 14780 8230
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14844 7954 14872 8570
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 5794 14780 7686
rect 14844 6934 14872 7890
rect 14936 7410 14964 10950
rect 15120 9674 15148 11172
rect 15028 9646 15148 9674
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14832 6928 14884 6934
rect 14832 6870 14884 6876
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14844 6186 14872 6598
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14752 5766 14872 5794
rect 14740 5704 14792 5710
rect 14738 5672 14740 5681
rect 14792 5672 14794 5681
rect 14738 5607 14794 5616
rect 14844 5386 14872 5766
rect 14752 5358 14872 5386
rect 14752 4826 14780 5358
rect 14832 5092 14884 5098
rect 14832 5034 14884 5040
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14108 3126 14136 3674
rect 14476 3466 14504 3878
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14568 3380 14596 4218
rect 14752 4185 14780 4762
rect 14738 4176 14794 4185
rect 14738 4111 14794 4120
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14568 3352 14688 3380
rect 14294 3292 14602 3301
rect 14294 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14516 3290 14540 3292
rect 14596 3290 14602 3292
rect 14356 3238 14358 3290
rect 14538 3238 14540 3290
rect 14294 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14516 3236 14540 3238
rect 14596 3236 14602 3238
rect 14294 3227 14602 3236
rect 14660 3126 14688 3352
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14188 3120 14240 3126
rect 14188 3062 14240 3068
rect 14556 3120 14608 3126
rect 14556 3062 14608 3068
rect 14648 3120 14700 3126
rect 14648 3062 14700 3068
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13832 800 13860 2790
rect 14108 2446 14136 3062
rect 14200 2774 14228 3062
rect 14372 2916 14424 2922
rect 14372 2858 14424 2864
rect 14384 2774 14412 2858
rect 14568 2774 14596 3062
rect 14200 2746 14412 2774
rect 14096 2440 14148 2446
rect 14384 2394 14412 2746
rect 14476 2746 14596 2774
rect 14476 2650 14504 2746
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14096 2382 14148 2388
rect 14200 2366 14412 2394
rect 14200 1986 14228 2366
rect 14294 2204 14602 2213
rect 14294 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14516 2202 14540 2204
rect 14596 2202 14602 2204
rect 14356 2150 14358 2202
rect 14538 2150 14540 2202
rect 14294 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14516 2148 14540 2150
rect 14596 2148 14602 2150
rect 14294 2139 14602 2148
rect 14200 1958 14320 1986
rect 14292 800 14320 1958
rect 14752 800 14780 3878
rect 14844 2446 14872 5034
rect 14924 4548 14976 4554
rect 14924 4490 14976 4496
rect 14936 3738 14964 4490
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 15028 3602 15056 9646
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15120 6866 15148 8774
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15120 5914 15148 6258
rect 15212 6118 15240 8298
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15304 5930 15332 11183
rect 15384 11154 15436 11160
rect 15488 10554 15516 13874
rect 15934 13424 15990 13433
rect 15934 13359 15990 13368
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15842 12880 15898 12889
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15580 11150 15608 11494
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15488 10526 15608 10554
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15396 7954 15424 8230
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 15488 7886 15516 8774
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15396 7546 15424 7686
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15488 7002 15516 7346
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15382 6896 15438 6905
rect 15382 6831 15438 6840
rect 15396 6225 15424 6831
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15488 6254 15516 6734
rect 15476 6248 15528 6254
rect 15382 6216 15438 6225
rect 15476 6190 15528 6196
rect 15382 6151 15438 6160
rect 15108 5908 15160 5914
rect 15304 5902 15424 5930
rect 15108 5850 15160 5856
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15212 5370 15240 5510
rect 15304 5370 15332 5714
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15396 5302 15424 5902
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 15396 4865 15424 5238
rect 15382 4856 15438 4865
rect 15382 4791 15438 4800
rect 15396 4758 15424 4791
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15580 4078 15608 10526
rect 15672 10266 15700 12854
rect 15842 12815 15898 12824
rect 15856 12306 15884 12815
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15948 12186 15976 13359
rect 16040 13258 16068 14855
rect 16118 14512 16174 14521
rect 16118 14447 16174 14456
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 16132 12434 16160 14447
rect 15764 12158 15976 12186
rect 16040 12406 16160 12434
rect 15764 11762 15792 12158
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15856 11354 15884 12038
rect 16040 11778 16068 12406
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 15948 11750 16068 11778
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15764 11218 15792 11290
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15764 10606 15792 11154
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15764 6746 15792 10406
rect 15856 7342 15884 11086
rect 15948 10470 15976 11750
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16040 11558 16068 11630
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15934 10160 15990 10169
rect 15934 10095 15990 10104
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15764 6718 15884 6746
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 6390 15792 6598
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15672 5914 15700 6190
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15764 5846 15792 6190
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 15856 5522 15884 6718
rect 15764 5494 15884 5522
rect 15764 5098 15792 5494
rect 15948 5386 15976 10095
rect 16040 9722 16068 11494
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16132 9586 16160 12242
rect 16224 11558 16252 16079
rect 16408 14414 16436 16400
rect 17052 14890 17080 16400
rect 17130 15328 17186 15337
rect 17130 15263 17186 15272
rect 17040 14884 17092 14890
rect 17040 14826 17092 14832
rect 16518 14716 16826 14725
rect 16518 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16740 14714 16764 14716
rect 16820 14714 16826 14716
rect 16580 14662 16582 14714
rect 16762 14662 16764 14714
rect 16518 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16740 14660 16764 14662
rect 16820 14660 16826 14662
rect 16518 14651 16826 14660
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16518 13628 16826 13637
rect 16518 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16740 13626 16764 13628
rect 16820 13626 16826 13628
rect 16580 13574 16582 13626
rect 16762 13574 16764 13626
rect 16518 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16740 13572 16764 13574
rect 16820 13572 16826 13574
rect 16518 13563 16826 13572
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16302 12064 16358 12073
rect 16302 11999 16358 12008
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16132 9110 16160 9522
rect 16316 9194 16344 11999
rect 16408 9926 16436 12582
rect 16518 12540 16826 12549
rect 16518 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16740 12538 16764 12540
rect 16820 12538 16826 12540
rect 16580 12486 16582 12538
rect 16762 12486 16764 12538
rect 16518 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16740 12484 16764 12486
rect 16820 12484 16826 12486
rect 16518 12475 16826 12484
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16776 11898 16804 12174
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16518 11452 16826 11461
rect 16518 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16740 11450 16764 11452
rect 16820 11450 16826 11452
rect 16580 11398 16582 11450
rect 16762 11398 16764 11450
rect 16518 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16740 11396 16764 11398
rect 16820 11396 16826 11398
rect 16518 11387 16826 11396
rect 16486 11112 16542 11121
rect 16486 11047 16542 11056
rect 16500 10742 16528 11047
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16518 10364 16826 10373
rect 16518 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16740 10362 16764 10364
rect 16820 10362 16826 10364
rect 16580 10310 16582 10362
rect 16762 10310 16764 10362
rect 16518 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16740 10308 16764 10310
rect 16820 10308 16826 10310
rect 16518 10299 16826 10308
rect 16868 10266 16896 10950
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16394 9480 16450 9489
rect 16394 9415 16450 9424
rect 16224 9178 16344 9194
rect 16408 9178 16436 9415
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16518 9276 16826 9285
rect 16518 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16740 9274 16764 9276
rect 16820 9274 16826 9276
rect 16580 9222 16582 9274
rect 16762 9222 16764 9274
rect 16518 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16740 9220 16764 9222
rect 16820 9220 16826 9222
rect 16518 9211 16826 9220
rect 16212 9172 16344 9178
rect 16264 9166 16344 9172
rect 16396 9172 16448 9178
rect 16212 9114 16264 9120
rect 16396 9114 16448 9120
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 16040 8566 16068 8978
rect 16408 8838 16436 9114
rect 16868 8974 16896 9318
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16120 8832 16172 8838
rect 16396 8832 16448 8838
rect 16120 8774 16172 8780
rect 16302 8800 16358 8809
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 16040 8430 16068 8502
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16132 7970 16160 8774
rect 16396 8774 16448 8780
rect 16302 8735 16358 8744
rect 16316 8634 16344 8735
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16040 7942 16160 7970
rect 16040 6905 16068 7942
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 16026 6896 16082 6905
rect 16026 6831 16082 6840
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 16040 6458 16068 6666
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16040 5710 16068 6054
rect 16132 5778 16160 7754
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 16224 6866 16252 7210
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16316 5846 16344 8570
rect 16518 8188 16826 8197
rect 16518 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16740 8186 16764 8188
rect 16820 8186 16826 8188
rect 16580 8134 16582 8186
rect 16762 8134 16764 8186
rect 16518 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16740 8132 16764 8134
rect 16820 8132 16826 8134
rect 16518 8123 16826 8132
rect 16396 7336 16448 7342
rect 16394 7304 16396 7313
rect 16448 7304 16450 7313
rect 16394 7239 16450 7248
rect 16518 7100 16826 7109
rect 16518 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16740 7098 16764 7100
rect 16820 7098 16826 7100
rect 16580 7046 16582 7098
rect 16762 7046 16764 7098
rect 16518 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16740 7044 16764 7046
rect 16820 7044 16826 7046
rect 16518 7035 16826 7044
rect 16868 6390 16896 8910
rect 16960 8022 16988 10610
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 17052 8634 17080 10066
rect 17144 9194 17172 15263
rect 17328 14482 17356 16510
rect 17682 16400 17738 16510
rect 18326 16400 18382 17200
rect 18970 16538 19026 17200
rect 18432 16510 19026 16538
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17224 11076 17276 11082
rect 17224 11018 17276 11024
rect 17236 10606 17264 11018
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17236 10130 17264 10542
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17328 9330 17356 14418
rect 18340 14346 18368 16400
rect 18328 14340 18380 14346
rect 18328 14282 18380 14288
rect 17868 12708 17920 12714
rect 17868 12650 17920 12656
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17420 11218 17448 11834
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17420 10266 17448 11154
rect 17880 11150 17908 12650
rect 18432 12209 18460 16510
rect 18970 16400 19026 16510
rect 19614 16400 19670 17200
rect 19628 14074 19656 16400
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 18418 12200 18474 12209
rect 18418 12135 18474 12144
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17498 10840 17554 10849
rect 17498 10775 17554 10784
rect 17512 10742 17540 10775
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17328 9302 17448 9330
rect 17144 9166 17356 9194
rect 17132 9104 17184 9110
rect 17132 9046 17184 9052
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 17144 7546 17172 9046
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17144 6866 17172 7142
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17040 6792 17092 6798
rect 17038 6760 17040 6769
rect 17092 6760 17094 6769
rect 17038 6695 17094 6704
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16960 6458 16988 6598
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16408 5914 16436 6258
rect 16518 6012 16826 6021
rect 16518 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16740 6010 16764 6012
rect 16820 6010 16826 6012
rect 16580 5958 16582 6010
rect 16762 5958 16764 6010
rect 16518 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16740 5956 16764 5958
rect 16820 5956 16826 5958
rect 16518 5947 16826 5956
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16304 5840 16356 5846
rect 16304 5782 16356 5788
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15856 5358 15976 5386
rect 15752 5092 15804 5098
rect 15752 5034 15804 5040
rect 15764 4826 15792 5034
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15856 4729 15884 5358
rect 16040 5302 16068 5646
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15842 4720 15898 4729
rect 15842 4655 15898 4664
rect 15948 4622 15976 5170
rect 16028 5160 16080 5166
rect 16132 5148 16160 5714
rect 16316 5642 16344 5782
rect 16868 5710 16896 6326
rect 17144 6254 17172 6802
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16868 5234 16896 5646
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16080 5120 16160 5148
rect 16028 5102 16080 5108
rect 16224 4826 16252 5170
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 15936 4616 15988 4622
rect 15934 4584 15936 4593
rect 15988 4584 15990 4593
rect 15934 4519 15990 4528
rect 16028 4480 16080 4486
rect 16080 4428 16160 4434
rect 16028 4422 16160 4428
rect 16040 4406 16160 4422
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15750 3768 15806 3777
rect 15750 3703 15752 3712
rect 15804 3703 15806 3712
rect 15752 3674 15804 3680
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15488 3058 15516 3606
rect 16132 3058 16160 4406
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 15476 2916 15528 2922
rect 15476 2858 15528 2864
rect 15488 2650 15516 2858
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 15212 800 15240 2518
rect 15764 1442 15792 2790
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 15672 1414 15792 1442
rect 15672 800 15700 1414
rect 16132 800 16160 2314
rect 9324 734 9536 762
rect 9678 0 9734 800
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16316 626 16344 4966
rect 16518 4924 16826 4933
rect 16518 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16740 4922 16764 4924
rect 16820 4922 16826 4924
rect 16580 4870 16582 4922
rect 16762 4870 16764 4922
rect 16518 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16740 4868 16764 4870
rect 16820 4868 16826 4870
rect 16518 4859 16826 4868
rect 16518 3836 16826 3845
rect 16518 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16740 3834 16764 3836
rect 16820 3834 16826 3836
rect 16580 3782 16582 3834
rect 16762 3782 16764 3834
rect 16518 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16740 3780 16764 3782
rect 16820 3780 16826 3782
rect 16518 3771 16826 3780
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16408 2632 16436 2790
rect 16518 2748 16826 2757
rect 16518 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16740 2746 16764 2748
rect 16820 2746 16826 2748
rect 16580 2694 16582 2746
rect 16762 2694 16764 2746
rect 16518 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16740 2692 16764 2694
rect 16820 2692 16826 2694
rect 16518 2683 16826 2692
rect 16408 2604 16620 2632
rect 16592 800 16620 2604
rect 16868 1465 16896 4966
rect 17132 4548 17184 4554
rect 17132 4490 17184 4496
rect 17144 3126 17172 4490
rect 17236 4321 17264 7686
rect 17328 6798 17356 9166
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17420 6610 17448 9302
rect 17512 9217 17540 9862
rect 17682 9616 17738 9625
rect 17682 9551 17684 9560
rect 17736 9551 17738 9560
rect 17684 9522 17736 9528
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17498 9208 17554 9217
rect 17972 9178 18000 9454
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 17498 9143 17554 9152
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17498 6896 17554 6905
rect 17498 6831 17554 6840
rect 17328 6582 17448 6610
rect 17222 4312 17278 4321
rect 17222 4247 17278 4256
rect 17328 3641 17356 6582
rect 17512 5914 17540 6831
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17512 5710 17540 5850
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17590 5672 17646 5681
rect 17590 5607 17646 5616
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17512 5273 17540 5510
rect 17604 5370 17632 5607
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17498 5264 17554 5273
rect 17498 5199 17554 5208
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17314 3632 17370 3641
rect 17314 3567 17370 3576
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 17420 3058 17448 4626
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 16854 1456 16910 1465
rect 16854 1391 16910 1400
rect 17052 800 17080 2790
rect 17512 800 17540 2790
rect 17696 1057 17724 8298
rect 17788 5953 17816 8774
rect 18064 8401 18092 9318
rect 18050 8392 18106 8401
rect 18050 8327 18106 8336
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18064 7410 18092 8026
rect 18156 7585 18184 11222
rect 18142 7576 18198 7585
rect 18142 7511 18198 7520
rect 18052 7404 18104 7410
rect 18104 7364 18184 7392
rect 18052 7346 18104 7352
rect 18052 7200 18104 7206
rect 18050 7168 18052 7177
rect 18104 7168 18106 7177
rect 18050 7103 18106 7112
rect 18156 7002 18184 7364
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18050 6352 18106 6361
rect 18050 6287 18106 6296
rect 17774 5944 17830 5953
rect 18064 5914 18092 6287
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 17774 5879 17830 5888
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18156 5710 18184 6122
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18248 5137 18276 11494
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18234 5128 18290 5137
rect 18234 5063 18290 5072
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17972 4729 18000 4966
rect 17958 4720 18014 4729
rect 17958 4655 18014 4664
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 3097 17816 4422
rect 17960 3936 18012 3942
rect 17958 3904 17960 3913
rect 18012 3904 18014 3913
rect 17958 3839 18014 3848
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17774 3088 17830 3097
rect 17880 3058 17908 3402
rect 17774 3023 17830 3032
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17682 1048 17738 1057
rect 17682 983 17738 992
rect 17972 800 18000 2790
rect 18340 2689 18368 10406
rect 18524 10033 18552 11018
rect 18510 10024 18566 10033
rect 18510 9959 18566 9968
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18432 7993 18460 9318
rect 18418 7984 18474 7993
rect 18418 7919 18474 7928
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18432 6769 18460 7142
rect 18418 6760 18474 6769
rect 18418 6695 18474 6704
rect 18420 5568 18472 5574
rect 18418 5536 18420 5545
rect 18472 5536 18474 5545
rect 18418 5471 18474 5480
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18326 2680 18382 2689
rect 18326 2615 18382 2624
rect 18052 2304 18104 2310
rect 18050 2272 18052 2281
rect 18104 2272 18106 2281
rect 18050 2207 18106 2216
rect 18432 800 18460 2790
rect 18524 1873 18552 9862
rect 18616 3505 18644 12038
rect 18602 3496 18658 3505
rect 18602 3431 18658 3440
rect 18880 2916 18932 2922
rect 18880 2858 18932 2864
rect 18510 1864 18566 1873
rect 18510 1799 18566 1808
rect 18892 800 18920 2858
rect 16394 640 16450 649
rect 16316 598 16394 626
rect 16394 575 16450 584
rect 16578 0 16634 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 18878 0 18934 800
<< via2 >>
rect 2778 16224 2834 16280
rect 2134 13776 2190 13832
rect 1582 10512 1638 10568
rect 1490 8200 1546 8256
rect 1398 8064 1454 8120
rect 1674 8880 1730 8936
rect 1582 7248 1638 7304
rect 1582 6452 1638 6488
rect 1582 6432 1584 6452
rect 1584 6432 1636 6452
rect 1636 6432 1638 6452
rect 1490 4428 1492 4448
rect 1492 4428 1544 4448
rect 1544 4428 1546 4448
rect 1490 4392 1546 4428
rect 1582 3576 1638 3632
rect 3054 16360 3110 16416
rect 2962 14612 3018 14648
rect 2962 14592 2964 14612
rect 2964 14592 3016 14612
rect 3016 14592 3018 14612
rect 3974 15816 4030 15872
rect 3790 15408 3846 15464
rect 3606 15000 3662 15056
rect 3180 14714 3236 14716
rect 3260 14714 3316 14716
rect 3340 14714 3396 14716
rect 3420 14714 3476 14716
rect 3180 14662 3226 14714
rect 3226 14662 3236 14714
rect 3260 14662 3290 14714
rect 3290 14662 3302 14714
rect 3302 14662 3316 14714
rect 3340 14662 3354 14714
rect 3354 14662 3366 14714
rect 3366 14662 3396 14714
rect 3420 14662 3430 14714
rect 3430 14662 3476 14714
rect 3180 14660 3236 14662
rect 3260 14660 3316 14662
rect 3340 14660 3396 14662
rect 3420 14660 3476 14662
rect 3180 13626 3236 13628
rect 3260 13626 3316 13628
rect 3340 13626 3396 13628
rect 3420 13626 3476 13628
rect 3180 13574 3226 13626
rect 3226 13574 3236 13626
rect 3260 13574 3290 13626
rect 3290 13574 3302 13626
rect 3302 13574 3316 13626
rect 3340 13574 3354 13626
rect 3354 13574 3366 13626
rect 3366 13574 3396 13626
rect 3420 13574 3430 13626
rect 3430 13574 3476 13626
rect 3180 13572 3236 13574
rect 3260 13572 3316 13574
rect 3340 13572 3396 13574
rect 3420 13572 3476 13574
rect 3180 12538 3236 12540
rect 3260 12538 3316 12540
rect 3340 12538 3396 12540
rect 3420 12538 3476 12540
rect 3180 12486 3226 12538
rect 3226 12486 3236 12538
rect 3260 12486 3290 12538
rect 3290 12486 3302 12538
rect 3302 12486 3316 12538
rect 3340 12486 3354 12538
rect 3354 12486 3366 12538
rect 3366 12486 3396 12538
rect 3420 12486 3430 12538
rect 3430 12486 3476 12538
rect 3180 12484 3236 12486
rect 3260 12484 3316 12486
rect 3340 12484 3396 12486
rect 3420 12484 3476 12486
rect 2042 6840 2098 6896
rect 1950 6740 1952 6760
rect 1952 6740 2004 6760
rect 2004 6740 2006 6760
rect 1950 6704 2006 6740
rect 2410 5208 2466 5264
rect 1398 2760 1454 2816
rect 2318 4004 2374 4040
rect 2318 3984 2320 4004
rect 2320 3984 2372 4004
rect 2372 3984 2374 4004
rect 2226 3168 2282 3224
rect 2686 10648 2742 10704
rect 3180 11450 3236 11452
rect 3260 11450 3316 11452
rect 3340 11450 3396 11452
rect 3420 11450 3476 11452
rect 3180 11398 3226 11450
rect 3226 11398 3236 11450
rect 3260 11398 3290 11450
rect 3290 11398 3302 11450
rect 3302 11398 3316 11450
rect 3340 11398 3354 11450
rect 3354 11398 3366 11450
rect 3366 11398 3396 11450
rect 3420 11398 3430 11450
rect 3430 11398 3476 11450
rect 3180 11396 3236 11398
rect 3260 11396 3316 11398
rect 3340 11396 3396 11398
rect 3420 11396 3476 11398
rect 3698 12688 3754 12744
rect 4158 14320 4214 14376
rect 4066 14184 4122 14240
rect 4066 13368 4122 13424
rect 3882 12824 3938 12880
rect 3606 11192 3662 11248
rect 3606 11056 3662 11112
rect 2778 8472 2834 8528
rect 2778 7792 2834 7848
rect 3180 10362 3236 10364
rect 3260 10362 3316 10364
rect 3340 10362 3396 10364
rect 3420 10362 3476 10364
rect 3180 10310 3226 10362
rect 3226 10310 3236 10362
rect 3260 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3316 10362
rect 3340 10310 3354 10362
rect 3354 10310 3366 10362
rect 3366 10310 3396 10362
rect 3420 10310 3430 10362
rect 3430 10310 3476 10362
rect 3180 10308 3236 10310
rect 3260 10308 3316 10310
rect 3340 10308 3396 10310
rect 3420 10308 3476 10310
rect 3180 9274 3236 9276
rect 3260 9274 3316 9276
rect 3340 9274 3396 9276
rect 3420 9274 3476 9276
rect 3180 9222 3226 9274
rect 3226 9222 3236 9274
rect 3260 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3316 9274
rect 3340 9222 3354 9274
rect 3354 9222 3366 9274
rect 3366 9222 3396 9274
rect 3420 9222 3430 9274
rect 3430 9222 3476 9274
rect 3180 9220 3236 9222
rect 3260 9220 3316 9222
rect 3340 9220 3396 9222
rect 3420 9220 3476 9222
rect 2962 8780 2964 8800
rect 2964 8780 3016 8800
rect 3016 8780 3018 8800
rect 2962 8744 3018 8780
rect 2870 5616 2926 5672
rect 3180 8186 3236 8188
rect 3260 8186 3316 8188
rect 3340 8186 3396 8188
rect 3420 8186 3476 8188
rect 3180 8134 3226 8186
rect 3226 8134 3236 8186
rect 3260 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3316 8186
rect 3340 8134 3354 8186
rect 3354 8134 3366 8186
rect 3366 8134 3396 8186
rect 3420 8134 3430 8186
rect 3430 8134 3476 8186
rect 3180 8132 3236 8134
rect 3260 8132 3316 8134
rect 3340 8132 3396 8134
rect 3420 8132 3476 8134
rect 3180 7098 3236 7100
rect 3260 7098 3316 7100
rect 3340 7098 3396 7100
rect 3420 7098 3476 7100
rect 3180 7046 3226 7098
rect 3226 7046 3236 7098
rect 3260 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3316 7098
rect 3340 7046 3354 7098
rect 3354 7046 3366 7098
rect 3366 7046 3396 7098
rect 3420 7046 3430 7098
rect 3430 7046 3476 7098
rect 3180 7044 3236 7046
rect 3260 7044 3316 7046
rect 3340 7044 3396 7046
rect 3420 7044 3476 7046
rect 3882 10512 3938 10568
rect 5404 14170 5460 14172
rect 5484 14170 5540 14172
rect 5564 14170 5620 14172
rect 5644 14170 5700 14172
rect 5404 14118 5450 14170
rect 5450 14118 5460 14170
rect 5484 14118 5514 14170
rect 5514 14118 5526 14170
rect 5526 14118 5540 14170
rect 5564 14118 5578 14170
rect 5578 14118 5590 14170
rect 5590 14118 5620 14170
rect 5644 14118 5654 14170
rect 5654 14118 5700 14170
rect 5404 14116 5460 14118
rect 5484 14116 5540 14118
rect 5564 14116 5620 14118
rect 5644 14116 5700 14118
rect 5262 13368 5318 13424
rect 5404 13082 5460 13084
rect 5484 13082 5540 13084
rect 5564 13082 5620 13084
rect 5644 13082 5700 13084
rect 5404 13030 5450 13082
rect 5450 13030 5460 13082
rect 5484 13030 5514 13082
rect 5514 13030 5526 13082
rect 5526 13030 5540 13082
rect 5564 13030 5578 13082
rect 5578 13030 5590 13082
rect 5590 13030 5620 13082
rect 5644 13030 5654 13082
rect 5654 13030 5700 13082
rect 5404 13028 5460 13030
rect 5484 13028 5540 13030
rect 5564 13028 5620 13030
rect 5644 13028 5700 13030
rect 4066 11756 4122 11792
rect 4066 11736 4068 11756
rect 4068 11736 4120 11756
rect 4120 11736 4122 11756
rect 4066 10956 4068 10976
rect 4068 10956 4120 10976
rect 4120 10956 4122 10976
rect 4066 10920 4122 10956
rect 4066 10104 4122 10160
rect 4342 9696 4398 9752
rect 4066 9424 4122 9480
rect 3790 7656 3846 7712
rect 3790 6432 3846 6488
rect 3180 6010 3236 6012
rect 3260 6010 3316 6012
rect 3340 6010 3396 6012
rect 3420 6010 3476 6012
rect 3180 5958 3226 6010
rect 3226 5958 3236 6010
rect 3260 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3316 6010
rect 3340 5958 3354 6010
rect 3354 5958 3366 6010
rect 3366 5958 3396 6010
rect 3420 5958 3430 6010
rect 3430 5958 3476 6010
rect 3180 5956 3236 5958
rect 3260 5956 3316 5958
rect 3340 5956 3396 5958
rect 3420 5956 3476 5958
rect 3054 5344 3110 5400
rect 3698 6160 3754 6216
rect 3882 5752 3938 5808
rect 3180 4922 3236 4924
rect 3260 4922 3316 4924
rect 3340 4922 3396 4924
rect 3420 4922 3476 4924
rect 3180 4870 3226 4922
rect 3226 4870 3236 4922
rect 3260 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3316 4922
rect 3340 4870 3354 4922
rect 3354 4870 3366 4922
rect 3366 4870 3396 4922
rect 3420 4870 3430 4922
rect 3430 4870 3476 4922
rect 3180 4868 3236 4870
rect 3260 4868 3316 4870
rect 3340 4868 3396 4870
rect 3420 4868 3476 4870
rect 2778 4800 2834 4856
rect 3054 4664 3110 4720
rect 3790 5072 3846 5128
rect 3238 4140 3294 4176
rect 3238 4120 3240 4140
rect 3240 4120 3292 4140
rect 3292 4120 3294 4140
rect 2686 3476 2688 3496
rect 2688 3476 2740 3496
rect 2740 3476 2742 3496
rect 2686 3440 2742 3476
rect 1950 1536 2006 1592
rect 2778 1944 2834 2000
rect 3180 3834 3236 3836
rect 3260 3834 3316 3836
rect 3340 3834 3396 3836
rect 3420 3834 3476 3836
rect 3180 3782 3226 3834
rect 3226 3782 3236 3834
rect 3260 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3316 3834
rect 3340 3782 3354 3834
rect 3354 3782 3366 3834
rect 3366 3782 3396 3834
rect 3420 3782 3430 3834
rect 3430 3782 3476 3834
rect 3180 3780 3236 3782
rect 3260 3780 3316 3782
rect 3340 3780 3396 3782
rect 3420 3780 3476 3782
rect 2962 2352 3018 2408
rect 3180 2746 3236 2748
rect 3260 2746 3316 2748
rect 3340 2746 3396 2748
rect 3420 2746 3476 2748
rect 3180 2694 3226 2746
rect 3226 2694 3236 2746
rect 3260 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3316 2746
rect 3340 2694 3354 2746
rect 3354 2694 3366 2746
rect 3366 2694 3396 2746
rect 3420 2694 3430 2746
rect 3430 2694 3476 2746
rect 3180 2692 3236 2694
rect 3260 2692 3316 2694
rect 3340 2692 3396 2694
rect 3420 2692 3476 2694
rect 3514 1128 3570 1184
rect 2870 312 2926 368
rect 3974 4664 4030 4720
rect 3882 4564 3884 4584
rect 3884 4564 3936 4584
rect 3936 4564 3938 4584
rect 3882 4528 3938 4564
rect 3790 856 3846 912
rect 5404 11994 5460 11996
rect 5484 11994 5540 11996
rect 5564 11994 5620 11996
rect 5644 11994 5700 11996
rect 5404 11942 5450 11994
rect 5450 11942 5460 11994
rect 5484 11942 5514 11994
rect 5514 11942 5526 11994
rect 5526 11942 5540 11994
rect 5564 11942 5578 11994
rect 5578 11942 5590 11994
rect 5590 11942 5620 11994
rect 5644 11942 5654 11994
rect 5654 11942 5700 11994
rect 5404 11940 5460 11942
rect 5484 11940 5540 11942
rect 5564 11940 5620 11942
rect 5644 11940 5700 11942
rect 5404 10906 5460 10908
rect 5484 10906 5540 10908
rect 5564 10906 5620 10908
rect 5644 10906 5700 10908
rect 5404 10854 5450 10906
rect 5450 10854 5460 10906
rect 5484 10854 5514 10906
rect 5514 10854 5526 10906
rect 5526 10854 5540 10906
rect 5564 10854 5578 10906
rect 5578 10854 5590 10906
rect 5590 10854 5620 10906
rect 5644 10854 5654 10906
rect 5654 10854 5700 10906
rect 5404 10852 5460 10854
rect 5484 10852 5540 10854
rect 5564 10852 5620 10854
rect 5644 10852 5700 10854
rect 5404 9818 5460 9820
rect 5484 9818 5540 9820
rect 5564 9818 5620 9820
rect 5644 9818 5700 9820
rect 5404 9766 5450 9818
rect 5450 9766 5460 9818
rect 5484 9766 5514 9818
rect 5514 9766 5526 9818
rect 5526 9766 5540 9818
rect 5564 9766 5578 9818
rect 5578 9766 5590 9818
rect 5590 9766 5620 9818
rect 5644 9766 5654 9818
rect 5654 9766 5700 9818
rect 5404 9764 5460 9766
rect 5484 9764 5540 9766
rect 5564 9764 5620 9766
rect 5644 9764 5700 9766
rect 5404 8730 5460 8732
rect 5484 8730 5540 8732
rect 5564 8730 5620 8732
rect 5644 8730 5700 8732
rect 5404 8678 5450 8730
rect 5450 8678 5460 8730
rect 5484 8678 5514 8730
rect 5514 8678 5526 8730
rect 5526 8678 5540 8730
rect 5564 8678 5578 8730
rect 5578 8678 5590 8730
rect 5590 8678 5620 8730
rect 5644 8678 5654 8730
rect 5654 8678 5700 8730
rect 5404 8676 5460 8678
rect 5484 8676 5540 8678
rect 5564 8676 5620 8678
rect 5644 8676 5700 8678
rect 5404 7642 5460 7644
rect 5484 7642 5540 7644
rect 5564 7642 5620 7644
rect 5644 7642 5700 7644
rect 5404 7590 5450 7642
rect 5450 7590 5460 7642
rect 5484 7590 5514 7642
rect 5514 7590 5526 7642
rect 5526 7590 5540 7642
rect 5564 7590 5578 7642
rect 5578 7590 5590 7642
rect 5590 7590 5620 7642
rect 5644 7590 5654 7642
rect 5654 7590 5700 7642
rect 5404 7588 5460 7590
rect 5484 7588 5540 7590
rect 5564 7588 5620 7590
rect 5644 7588 5700 7590
rect 5078 3052 5134 3088
rect 5078 3032 5080 3052
rect 5080 3032 5132 3052
rect 5132 3032 5134 3052
rect 5404 6554 5460 6556
rect 5484 6554 5540 6556
rect 5564 6554 5620 6556
rect 5644 6554 5700 6556
rect 5404 6502 5450 6554
rect 5450 6502 5460 6554
rect 5484 6502 5514 6554
rect 5514 6502 5526 6554
rect 5526 6502 5540 6554
rect 5564 6502 5578 6554
rect 5578 6502 5590 6554
rect 5590 6502 5620 6554
rect 5644 6502 5654 6554
rect 5654 6502 5700 6554
rect 5404 6500 5460 6502
rect 5484 6500 5540 6502
rect 5564 6500 5620 6502
rect 5644 6500 5700 6502
rect 5404 5466 5460 5468
rect 5484 5466 5540 5468
rect 5564 5466 5620 5468
rect 5644 5466 5700 5468
rect 5404 5414 5450 5466
rect 5450 5414 5460 5466
rect 5484 5414 5514 5466
rect 5514 5414 5526 5466
rect 5526 5414 5540 5466
rect 5564 5414 5578 5466
rect 5578 5414 5590 5466
rect 5590 5414 5620 5466
rect 5644 5414 5654 5466
rect 5654 5414 5700 5466
rect 5404 5412 5460 5414
rect 5484 5412 5540 5414
rect 5564 5412 5620 5414
rect 5644 5412 5700 5414
rect 5906 4800 5962 4856
rect 5404 4378 5460 4380
rect 5484 4378 5540 4380
rect 5564 4378 5620 4380
rect 5644 4378 5700 4380
rect 5404 4326 5450 4378
rect 5450 4326 5460 4378
rect 5484 4326 5514 4378
rect 5514 4326 5526 4378
rect 5526 4326 5540 4378
rect 5564 4326 5578 4378
rect 5578 4326 5590 4378
rect 5590 4326 5620 4378
rect 5644 4326 5654 4378
rect 5654 4326 5700 4378
rect 5404 4324 5460 4326
rect 5484 4324 5540 4326
rect 5564 4324 5620 4326
rect 5644 4324 5700 4326
rect 5404 3290 5460 3292
rect 5484 3290 5540 3292
rect 5564 3290 5620 3292
rect 5644 3290 5700 3292
rect 5404 3238 5450 3290
rect 5450 3238 5460 3290
rect 5484 3238 5514 3290
rect 5514 3238 5526 3290
rect 5526 3238 5540 3290
rect 5564 3238 5578 3290
rect 5578 3238 5590 3290
rect 5590 3238 5620 3290
rect 5644 3238 5654 3290
rect 5654 3238 5700 3290
rect 5404 3236 5460 3238
rect 5484 3236 5540 3238
rect 5564 3236 5620 3238
rect 5644 3236 5700 3238
rect 5404 2202 5460 2204
rect 5484 2202 5540 2204
rect 5564 2202 5620 2204
rect 5644 2202 5700 2204
rect 5404 2150 5450 2202
rect 5450 2150 5460 2202
rect 5484 2150 5514 2202
rect 5514 2150 5526 2202
rect 5526 2150 5540 2202
rect 5564 2150 5578 2202
rect 5578 2150 5590 2202
rect 5590 2150 5620 2202
rect 5644 2150 5654 2202
rect 5654 2150 5700 2202
rect 5404 2148 5460 2150
rect 5484 2148 5540 2150
rect 5564 2148 5620 2150
rect 5644 2148 5700 2150
rect 6458 11600 6514 11656
rect 6550 6196 6552 6216
rect 6552 6196 6604 6216
rect 6604 6196 6606 6216
rect 6550 6160 6606 6196
rect 7628 14714 7684 14716
rect 7708 14714 7764 14716
rect 7788 14714 7844 14716
rect 7868 14714 7924 14716
rect 7628 14662 7674 14714
rect 7674 14662 7684 14714
rect 7708 14662 7738 14714
rect 7738 14662 7750 14714
rect 7750 14662 7764 14714
rect 7788 14662 7802 14714
rect 7802 14662 7814 14714
rect 7814 14662 7844 14714
rect 7868 14662 7878 14714
rect 7878 14662 7924 14714
rect 7628 14660 7684 14662
rect 7708 14660 7764 14662
rect 7788 14660 7844 14662
rect 7868 14660 7924 14662
rect 7628 13626 7684 13628
rect 7708 13626 7764 13628
rect 7788 13626 7844 13628
rect 7868 13626 7924 13628
rect 7628 13574 7674 13626
rect 7674 13574 7684 13626
rect 7708 13574 7738 13626
rect 7738 13574 7750 13626
rect 7750 13574 7764 13626
rect 7788 13574 7802 13626
rect 7802 13574 7814 13626
rect 7814 13574 7844 13626
rect 7868 13574 7878 13626
rect 7878 13574 7924 13626
rect 7628 13572 7684 13574
rect 7708 13572 7764 13574
rect 7788 13572 7844 13574
rect 7868 13572 7924 13574
rect 7628 12538 7684 12540
rect 7708 12538 7764 12540
rect 7788 12538 7844 12540
rect 7868 12538 7924 12540
rect 7628 12486 7674 12538
rect 7674 12486 7684 12538
rect 7708 12486 7738 12538
rect 7738 12486 7750 12538
rect 7750 12486 7764 12538
rect 7788 12486 7802 12538
rect 7802 12486 7814 12538
rect 7814 12486 7844 12538
rect 7868 12486 7878 12538
rect 7878 12486 7924 12538
rect 7628 12484 7684 12486
rect 7708 12484 7764 12486
rect 7788 12484 7844 12486
rect 7868 12484 7924 12486
rect 7628 11450 7684 11452
rect 7708 11450 7764 11452
rect 7788 11450 7844 11452
rect 7868 11450 7924 11452
rect 7628 11398 7674 11450
rect 7674 11398 7684 11450
rect 7708 11398 7738 11450
rect 7738 11398 7750 11450
rect 7750 11398 7764 11450
rect 7788 11398 7802 11450
rect 7802 11398 7814 11450
rect 7814 11398 7844 11450
rect 7868 11398 7878 11450
rect 7878 11398 7924 11450
rect 7628 11396 7684 11398
rect 7708 11396 7764 11398
rect 7788 11396 7844 11398
rect 7868 11396 7924 11398
rect 7628 10362 7684 10364
rect 7708 10362 7764 10364
rect 7788 10362 7844 10364
rect 7868 10362 7924 10364
rect 7628 10310 7674 10362
rect 7674 10310 7684 10362
rect 7708 10310 7738 10362
rect 7738 10310 7750 10362
rect 7750 10310 7764 10362
rect 7788 10310 7802 10362
rect 7802 10310 7814 10362
rect 7814 10310 7844 10362
rect 7868 10310 7878 10362
rect 7878 10310 7924 10362
rect 7628 10308 7684 10310
rect 7708 10308 7764 10310
rect 7788 10308 7844 10310
rect 7868 10308 7924 10310
rect 8850 13932 8906 13968
rect 8850 13912 8852 13932
rect 8852 13912 8904 13932
rect 8904 13912 8906 13932
rect 8574 11212 8630 11248
rect 8574 11192 8576 11212
rect 8576 11192 8628 11212
rect 8628 11192 8630 11212
rect 7628 9274 7684 9276
rect 7708 9274 7764 9276
rect 7788 9274 7844 9276
rect 7868 9274 7924 9276
rect 7628 9222 7674 9274
rect 7674 9222 7684 9274
rect 7708 9222 7738 9274
rect 7738 9222 7750 9274
rect 7750 9222 7764 9274
rect 7788 9222 7802 9274
rect 7802 9222 7814 9274
rect 7814 9222 7844 9274
rect 7868 9222 7878 9274
rect 7878 9222 7924 9274
rect 7628 9220 7684 9222
rect 7708 9220 7764 9222
rect 7788 9220 7844 9222
rect 7868 9220 7924 9222
rect 7562 9016 7618 9072
rect 7628 8186 7684 8188
rect 7708 8186 7764 8188
rect 7788 8186 7844 8188
rect 7868 8186 7924 8188
rect 7628 8134 7674 8186
rect 7674 8134 7684 8186
rect 7708 8134 7738 8186
rect 7738 8134 7750 8186
rect 7750 8134 7764 8186
rect 7788 8134 7802 8186
rect 7802 8134 7814 8186
rect 7814 8134 7844 8186
rect 7868 8134 7878 8186
rect 7878 8134 7924 8186
rect 7628 8132 7684 8134
rect 7708 8132 7764 8134
rect 7788 8132 7844 8134
rect 7868 8132 7924 8134
rect 7628 7098 7684 7100
rect 7708 7098 7764 7100
rect 7788 7098 7844 7100
rect 7868 7098 7924 7100
rect 7628 7046 7674 7098
rect 7674 7046 7684 7098
rect 7708 7046 7738 7098
rect 7738 7046 7750 7098
rect 7750 7046 7764 7098
rect 7788 7046 7802 7098
rect 7802 7046 7814 7098
rect 7814 7046 7844 7098
rect 7868 7046 7878 7098
rect 7878 7046 7924 7098
rect 7628 7044 7684 7046
rect 7708 7044 7764 7046
rect 7788 7044 7844 7046
rect 7868 7044 7924 7046
rect 7628 6010 7684 6012
rect 7708 6010 7764 6012
rect 7788 6010 7844 6012
rect 7868 6010 7924 6012
rect 7628 5958 7674 6010
rect 7674 5958 7684 6010
rect 7708 5958 7738 6010
rect 7738 5958 7750 6010
rect 7750 5958 7764 6010
rect 7788 5958 7802 6010
rect 7802 5958 7814 6010
rect 7814 5958 7844 6010
rect 7868 5958 7878 6010
rect 7878 5958 7924 6010
rect 7628 5956 7684 5958
rect 7708 5956 7764 5958
rect 7788 5956 7844 5958
rect 7868 5956 7924 5958
rect 7628 4922 7684 4924
rect 7708 4922 7764 4924
rect 7788 4922 7844 4924
rect 7868 4922 7924 4924
rect 7628 4870 7674 4922
rect 7674 4870 7684 4922
rect 7708 4870 7738 4922
rect 7738 4870 7750 4922
rect 7750 4870 7764 4922
rect 7788 4870 7802 4922
rect 7802 4870 7814 4922
rect 7814 4870 7844 4922
rect 7868 4870 7878 4922
rect 7878 4870 7924 4922
rect 7628 4868 7684 4870
rect 7708 4868 7764 4870
rect 7788 4868 7844 4870
rect 7868 4868 7924 4870
rect 7470 4684 7526 4720
rect 7470 4664 7472 4684
rect 7472 4664 7524 4684
rect 7524 4664 7526 4684
rect 7628 3834 7684 3836
rect 7708 3834 7764 3836
rect 7788 3834 7844 3836
rect 7868 3834 7924 3836
rect 7628 3782 7674 3834
rect 7674 3782 7684 3834
rect 7708 3782 7738 3834
rect 7738 3782 7750 3834
rect 7750 3782 7764 3834
rect 7788 3782 7802 3834
rect 7802 3782 7814 3834
rect 7814 3782 7844 3834
rect 7868 3782 7878 3834
rect 7878 3782 7924 3834
rect 7628 3780 7684 3782
rect 7708 3780 7764 3782
rect 7788 3780 7844 3782
rect 7868 3780 7924 3782
rect 8758 3984 8814 4040
rect 7378 2896 7434 2952
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9898 14170
rect 9898 14118 9908 14170
rect 9932 14118 9962 14170
rect 9962 14118 9974 14170
rect 9974 14118 9988 14170
rect 10012 14118 10026 14170
rect 10026 14118 10038 14170
rect 10038 14118 10068 14170
rect 10092 14118 10102 14170
rect 10102 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9126 13776 9182 13832
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9898 13082
rect 9898 13030 9908 13082
rect 9932 13030 9962 13082
rect 9962 13030 9974 13082
rect 9974 13030 9988 13082
rect 10012 13030 10026 13082
rect 10026 13030 10038 13082
rect 10038 13030 10068 13082
rect 10092 13030 10102 13082
rect 10102 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9770 12280 9826 12336
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9898 11994
rect 9898 11942 9908 11994
rect 9932 11942 9962 11994
rect 9962 11942 9974 11994
rect 9974 11942 9988 11994
rect 10012 11942 10026 11994
rect 10026 11942 10038 11994
rect 10038 11942 10068 11994
rect 10092 11942 10102 11994
rect 10102 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9898 10906
rect 9898 10854 9908 10906
rect 9932 10854 9962 10906
rect 9962 10854 9974 10906
rect 9974 10854 9988 10906
rect 10012 10854 10026 10906
rect 10026 10854 10038 10906
rect 10038 10854 10068 10906
rect 10092 10854 10102 10906
rect 10102 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9898 9818
rect 9898 9766 9908 9818
rect 9932 9766 9962 9818
rect 9962 9766 9974 9818
rect 9974 9766 9988 9818
rect 10012 9766 10026 9818
rect 10026 9766 10038 9818
rect 10038 9766 10068 9818
rect 10092 9766 10102 9818
rect 10102 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9898 8730
rect 9898 8678 9908 8730
rect 9932 8678 9962 8730
rect 9962 8678 9974 8730
rect 9974 8678 9988 8730
rect 10012 8678 10026 8730
rect 10026 8678 10038 8730
rect 10038 8678 10068 8730
rect 10092 8678 10102 8730
rect 10102 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9898 7642
rect 9898 7590 9908 7642
rect 9932 7590 9962 7642
rect 9962 7590 9974 7642
rect 9974 7590 9988 7642
rect 10012 7590 10026 7642
rect 10026 7590 10038 7642
rect 10038 7590 10068 7642
rect 10092 7590 10102 7642
rect 10102 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9898 6554
rect 9898 6502 9908 6554
rect 9932 6502 9962 6554
rect 9962 6502 9974 6554
rect 9974 6502 9988 6554
rect 10012 6502 10026 6554
rect 10026 6502 10038 6554
rect 10038 6502 10068 6554
rect 10092 6502 10102 6554
rect 10102 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9898 5466
rect 9898 5414 9908 5466
rect 9932 5414 9962 5466
rect 9962 5414 9974 5466
rect 9974 5414 9988 5466
rect 10012 5414 10026 5466
rect 10026 5414 10038 5466
rect 10038 5414 10068 5466
rect 10092 5414 10102 5466
rect 10102 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 7628 2746 7684 2748
rect 7708 2746 7764 2748
rect 7788 2746 7844 2748
rect 7868 2746 7924 2748
rect 7628 2694 7674 2746
rect 7674 2694 7684 2746
rect 7708 2694 7738 2746
rect 7738 2694 7750 2746
rect 7750 2694 7764 2746
rect 7788 2694 7802 2746
rect 7802 2694 7814 2746
rect 7814 2694 7844 2746
rect 7868 2694 7878 2746
rect 7878 2694 7924 2746
rect 7628 2692 7684 2694
rect 7708 2692 7764 2694
rect 7788 2692 7844 2694
rect 7868 2692 7924 2694
rect 9310 3984 9366 4040
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9898 4378
rect 9898 4326 9908 4378
rect 9932 4326 9962 4378
rect 9962 4326 9974 4378
rect 9974 4326 9988 4378
rect 10012 4326 10026 4378
rect 10026 4326 10038 4378
rect 10038 4326 10068 4378
rect 10092 4326 10102 4378
rect 10102 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 9678 3984 9734 4040
rect 10506 12708 10562 12744
rect 10506 12688 10508 12708
rect 10508 12688 10560 12708
rect 10560 12688 10562 12708
rect 10506 11056 10562 11112
rect 10506 3440 10562 3496
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9898 3290
rect 9898 3238 9908 3290
rect 9932 3238 9962 3290
rect 9962 3238 9974 3290
rect 9974 3238 9988 3290
rect 10012 3238 10026 3290
rect 10026 3238 10038 3290
rect 10038 3238 10068 3290
rect 10092 3238 10102 3290
rect 10102 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9898 2202
rect 9898 2150 9908 2202
rect 9932 2150 9962 2202
rect 9962 2150 9974 2202
rect 9974 2150 9988 2202
rect 10012 2150 10026 2202
rect 10026 2150 10038 2202
rect 10038 2150 10068 2202
rect 10092 2150 10102 2202
rect 10102 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 12076 14714 12132 14716
rect 12156 14714 12212 14716
rect 12236 14714 12292 14716
rect 12316 14714 12372 14716
rect 12076 14662 12122 14714
rect 12122 14662 12132 14714
rect 12156 14662 12186 14714
rect 12186 14662 12198 14714
rect 12198 14662 12212 14714
rect 12236 14662 12250 14714
rect 12250 14662 12262 14714
rect 12262 14662 12292 14714
rect 12316 14662 12326 14714
rect 12326 14662 12372 14714
rect 12076 14660 12132 14662
rect 12156 14660 12212 14662
rect 12236 14660 12292 14662
rect 12316 14660 12372 14662
rect 12076 13626 12132 13628
rect 12156 13626 12212 13628
rect 12236 13626 12292 13628
rect 12316 13626 12372 13628
rect 12076 13574 12122 13626
rect 12122 13574 12132 13626
rect 12156 13574 12186 13626
rect 12186 13574 12198 13626
rect 12198 13574 12212 13626
rect 12236 13574 12250 13626
rect 12250 13574 12262 13626
rect 12262 13574 12292 13626
rect 12316 13574 12326 13626
rect 12326 13574 12372 13626
rect 12076 13572 12132 13574
rect 12156 13572 12212 13574
rect 12236 13572 12292 13574
rect 12316 13572 12372 13574
rect 12076 12538 12132 12540
rect 12156 12538 12212 12540
rect 12236 12538 12292 12540
rect 12316 12538 12372 12540
rect 12076 12486 12122 12538
rect 12122 12486 12132 12538
rect 12156 12486 12186 12538
rect 12186 12486 12198 12538
rect 12198 12486 12212 12538
rect 12236 12486 12250 12538
rect 12250 12486 12262 12538
rect 12262 12486 12292 12538
rect 12316 12486 12326 12538
rect 12326 12486 12372 12538
rect 12076 12484 12132 12486
rect 12156 12484 12212 12486
rect 12236 12484 12292 12486
rect 12316 12484 12372 12486
rect 12076 11450 12132 11452
rect 12156 11450 12212 11452
rect 12236 11450 12292 11452
rect 12316 11450 12372 11452
rect 12076 11398 12122 11450
rect 12122 11398 12132 11450
rect 12156 11398 12186 11450
rect 12186 11398 12198 11450
rect 12198 11398 12212 11450
rect 12236 11398 12250 11450
rect 12250 11398 12262 11450
rect 12262 11398 12292 11450
rect 12316 11398 12326 11450
rect 12326 11398 12372 11450
rect 12076 11396 12132 11398
rect 12156 11396 12212 11398
rect 12236 11396 12292 11398
rect 12316 11396 12372 11398
rect 12076 10362 12132 10364
rect 12156 10362 12212 10364
rect 12236 10362 12292 10364
rect 12316 10362 12372 10364
rect 12076 10310 12122 10362
rect 12122 10310 12132 10362
rect 12156 10310 12186 10362
rect 12186 10310 12198 10362
rect 12198 10310 12212 10362
rect 12236 10310 12250 10362
rect 12250 10310 12262 10362
rect 12262 10310 12292 10362
rect 12316 10310 12326 10362
rect 12326 10310 12372 10362
rect 12076 10308 12132 10310
rect 12156 10308 12212 10310
rect 12236 10308 12292 10310
rect 12316 10308 12372 10310
rect 12076 9274 12132 9276
rect 12156 9274 12212 9276
rect 12236 9274 12292 9276
rect 12316 9274 12372 9276
rect 12076 9222 12122 9274
rect 12122 9222 12132 9274
rect 12156 9222 12186 9274
rect 12186 9222 12198 9274
rect 12198 9222 12212 9274
rect 12236 9222 12250 9274
rect 12250 9222 12262 9274
rect 12262 9222 12292 9274
rect 12316 9222 12326 9274
rect 12326 9222 12372 9274
rect 12076 9220 12132 9222
rect 12156 9220 12212 9222
rect 12236 9220 12292 9222
rect 12316 9220 12372 9222
rect 12076 8186 12132 8188
rect 12156 8186 12212 8188
rect 12236 8186 12292 8188
rect 12316 8186 12372 8188
rect 12076 8134 12122 8186
rect 12122 8134 12132 8186
rect 12156 8134 12186 8186
rect 12186 8134 12198 8186
rect 12198 8134 12212 8186
rect 12236 8134 12250 8186
rect 12250 8134 12262 8186
rect 12262 8134 12292 8186
rect 12316 8134 12326 8186
rect 12326 8134 12372 8186
rect 12076 8132 12132 8134
rect 12156 8132 12212 8134
rect 12236 8132 12292 8134
rect 12316 8132 12372 8134
rect 12076 7098 12132 7100
rect 12156 7098 12212 7100
rect 12236 7098 12292 7100
rect 12316 7098 12372 7100
rect 12076 7046 12122 7098
rect 12122 7046 12132 7098
rect 12156 7046 12186 7098
rect 12186 7046 12198 7098
rect 12198 7046 12212 7098
rect 12236 7046 12250 7098
rect 12250 7046 12262 7098
rect 12262 7046 12292 7098
rect 12316 7046 12326 7098
rect 12326 7046 12372 7098
rect 12076 7044 12132 7046
rect 12156 7044 12212 7046
rect 12236 7044 12292 7046
rect 12316 7044 12372 7046
rect 12076 6010 12132 6012
rect 12156 6010 12212 6012
rect 12236 6010 12292 6012
rect 12316 6010 12372 6012
rect 12076 5958 12122 6010
rect 12122 5958 12132 6010
rect 12156 5958 12186 6010
rect 12186 5958 12198 6010
rect 12198 5958 12212 6010
rect 12236 5958 12250 6010
rect 12250 5958 12262 6010
rect 12262 5958 12292 6010
rect 12316 5958 12326 6010
rect 12326 5958 12372 6010
rect 12076 5956 12132 5958
rect 12156 5956 12212 5958
rect 12236 5956 12292 5958
rect 12316 5956 12372 5958
rect 12076 4922 12132 4924
rect 12156 4922 12212 4924
rect 12236 4922 12292 4924
rect 12316 4922 12372 4924
rect 12076 4870 12122 4922
rect 12122 4870 12132 4922
rect 12156 4870 12186 4922
rect 12186 4870 12198 4922
rect 12198 4870 12212 4922
rect 12236 4870 12250 4922
rect 12250 4870 12262 4922
rect 12262 4870 12292 4922
rect 12316 4870 12326 4922
rect 12326 4870 12372 4922
rect 12076 4868 12132 4870
rect 12156 4868 12212 4870
rect 12236 4868 12292 4870
rect 12316 4868 12372 4870
rect 12622 14320 12678 14376
rect 12806 11600 12862 11656
rect 15474 16496 15530 16552
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14540 14170 14596 14172
rect 14300 14118 14346 14170
rect 14346 14118 14356 14170
rect 14380 14118 14410 14170
rect 14410 14118 14422 14170
rect 14422 14118 14436 14170
rect 14460 14118 14474 14170
rect 14474 14118 14486 14170
rect 14486 14118 14516 14170
rect 14540 14118 14550 14170
rect 14550 14118 14596 14170
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 14540 14116 14596 14118
rect 13818 13640 13874 13696
rect 13174 12144 13230 12200
rect 12530 3984 12586 4040
rect 12076 3834 12132 3836
rect 12156 3834 12212 3836
rect 12236 3834 12292 3836
rect 12316 3834 12372 3836
rect 12076 3782 12122 3834
rect 12122 3782 12132 3834
rect 12156 3782 12186 3834
rect 12186 3782 12198 3834
rect 12198 3782 12212 3834
rect 12236 3782 12250 3834
rect 12250 3782 12262 3834
rect 12262 3782 12292 3834
rect 12316 3782 12326 3834
rect 12326 3782 12372 3834
rect 12076 3780 12132 3782
rect 12156 3780 12212 3782
rect 12236 3780 12292 3782
rect 12316 3780 12372 3782
rect 11150 2896 11206 2952
rect 11794 2760 11850 2816
rect 12622 3576 12678 3632
rect 12070 2896 12126 2952
rect 12076 2746 12132 2748
rect 12156 2746 12212 2748
rect 12236 2746 12292 2748
rect 12316 2746 12372 2748
rect 12076 2694 12122 2746
rect 12122 2694 12132 2746
rect 12156 2694 12186 2746
rect 12186 2694 12198 2746
rect 12198 2694 12212 2746
rect 12236 2694 12250 2746
rect 12250 2694 12262 2746
rect 12262 2694 12292 2746
rect 12316 2694 12326 2746
rect 12326 2694 12372 2746
rect 12076 2692 12132 2694
rect 12156 2692 12212 2694
rect 12236 2692 12292 2694
rect 12316 2692 12372 2694
rect 13542 5208 13598 5264
rect 13542 4820 13598 4856
rect 13818 10648 13874 10704
rect 13726 5208 13782 5264
rect 13542 4800 13544 4820
rect 13544 4800 13596 4820
rect 13596 4800 13598 4820
rect 13818 3032 13874 3088
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14540 13082 14596 13084
rect 14300 13030 14346 13082
rect 14346 13030 14356 13082
rect 14380 13030 14410 13082
rect 14410 13030 14422 13082
rect 14422 13030 14436 13082
rect 14460 13030 14474 13082
rect 14474 13030 14486 13082
rect 14486 13030 14516 13082
rect 14540 13030 14550 13082
rect 14550 13030 14596 13082
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 14540 13028 14596 13030
rect 14278 12688 14334 12744
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14540 11994 14596 11996
rect 14300 11942 14346 11994
rect 14346 11942 14356 11994
rect 14380 11942 14410 11994
rect 14410 11942 14422 11994
rect 14422 11942 14436 11994
rect 14460 11942 14474 11994
rect 14474 11942 14486 11994
rect 14486 11942 14516 11994
rect 14540 11942 14550 11994
rect 14550 11942 14596 11994
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14540 11940 14596 11942
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14540 10906 14596 10908
rect 14300 10854 14346 10906
rect 14346 10854 14356 10906
rect 14380 10854 14410 10906
rect 14410 10854 14422 10906
rect 14422 10854 14436 10906
rect 14460 10854 14474 10906
rect 14474 10854 14486 10906
rect 14486 10854 14516 10906
rect 14540 10854 14550 10906
rect 14550 10854 14596 10906
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14540 10852 14596 10854
rect 14462 10548 14464 10568
rect 14464 10548 14516 10568
rect 14516 10548 14518 10568
rect 14462 10512 14518 10548
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14540 9818 14596 9820
rect 14300 9766 14346 9818
rect 14346 9766 14356 9818
rect 14380 9766 14410 9818
rect 14410 9766 14422 9818
rect 14422 9766 14436 9818
rect 14460 9766 14474 9818
rect 14474 9766 14486 9818
rect 14486 9766 14516 9818
rect 14540 9766 14550 9818
rect 14550 9766 14596 9818
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14540 9764 14596 9766
rect 15290 15680 15346 15736
rect 15014 13368 15070 13424
rect 16210 16088 16266 16144
rect 16026 14864 16082 14920
rect 15842 14048 15898 14104
rect 15198 13268 15200 13288
rect 15200 13268 15252 13288
rect 15252 13268 15254 13288
rect 15198 13232 15254 13268
rect 15290 11192 15346 11248
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14540 8730 14596 8732
rect 14300 8678 14346 8730
rect 14346 8678 14356 8730
rect 14380 8678 14410 8730
rect 14410 8678 14422 8730
rect 14422 8678 14436 8730
rect 14460 8678 14474 8730
rect 14474 8678 14486 8730
rect 14486 8678 14516 8730
rect 14540 8678 14550 8730
rect 14550 8678 14596 8730
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14540 8676 14596 8678
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14540 7642 14596 7644
rect 14300 7590 14346 7642
rect 14346 7590 14356 7642
rect 14380 7590 14410 7642
rect 14410 7590 14422 7642
rect 14422 7590 14436 7642
rect 14460 7590 14474 7642
rect 14474 7590 14486 7642
rect 14486 7590 14516 7642
rect 14540 7590 14550 7642
rect 14550 7590 14596 7642
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14540 7588 14596 7590
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14540 6554 14596 6556
rect 14300 6502 14346 6554
rect 14346 6502 14356 6554
rect 14380 6502 14410 6554
rect 14410 6502 14422 6554
rect 14422 6502 14436 6554
rect 14460 6502 14474 6554
rect 14474 6502 14486 6554
rect 14486 6502 14516 6554
rect 14540 6502 14550 6554
rect 14550 6502 14596 6554
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 14540 6500 14596 6502
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14540 5466 14596 5468
rect 14300 5414 14346 5466
rect 14346 5414 14356 5466
rect 14380 5414 14410 5466
rect 14410 5414 14422 5466
rect 14422 5414 14436 5466
rect 14460 5414 14474 5466
rect 14474 5414 14486 5466
rect 14486 5414 14516 5466
rect 14540 5414 14550 5466
rect 14550 5414 14596 5466
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 14540 5412 14596 5414
rect 14094 5072 14150 5128
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14540 4378 14596 4380
rect 14300 4326 14346 4378
rect 14346 4326 14356 4378
rect 14380 4326 14410 4378
rect 14410 4326 14422 4378
rect 14422 4326 14436 4378
rect 14460 4326 14474 4378
rect 14474 4326 14486 4378
rect 14486 4326 14516 4378
rect 14540 4326 14550 4378
rect 14550 4326 14596 4378
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 14540 4324 14596 4326
rect 14738 5652 14740 5672
rect 14740 5652 14792 5672
rect 14792 5652 14794 5672
rect 14738 5616 14794 5652
rect 14738 4120 14794 4176
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14540 3290 14596 3292
rect 14300 3238 14346 3290
rect 14346 3238 14356 3290
rect 14380 3238 14410 3290
rect 14410 3238 14422 3290
rect 14422 3238 14436 3290
rect 14460 3238 14474 3290
rect 14474 3238 14486 3290
rect 14486 3238 14516 3290
rect 14540 3238 14550 3290
rect 14550 3238 14596 3290
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 14540 3236 14596 3238
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14540 2202 14596 2204
rect 14300 2150 14346 2202
rect 14346 2150 14356 2202
rect 14380 2150 14410 2202
rect 14410 2150 14422 2202
rect 14422 2150 14436 2202
rect 14460 2150 14474 2202
rect 14474 2150 14486 2202
rect 14486 2150 14516 2202
rect 14540 2150 14550 2202
rect 14550 2150 14596 2202
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 14540 2148 14596 2150
rect 15934 13368 15990 13424
rect 15382 6840 15438 6896
rect 15382 6160 15438 6216
rect 15382 4800 15438 4856
rect 15842 12824 15898 12880
rect 16118 14456 16174 14512
rect 15934 10104 15990 10160
rect 17130 15272 17186 15328
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16764 14714 16820 14716
rect 16524 14662 16570 14714
rect 16570 14662 16580 14714
rect 16604 14662 16634 14714
rect 16634 14662 16646 14714
rect 16646 14662 16660 14714
rect 16684 14662 16698 14714
rect 16698 14662 16710 14714
rect 16710 14662 16740 14714
rect 16764 14662 16774 14714
rect 16774 14662 16820 14714
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16764 14660 16820 14662
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16764 13626 16820 13628
rect 16524 13574 16570 13626
rect 16570 13574 16580 13626
rect 16604 13574 16634 13626
rect 16634 13574 16646 13626
rect 16646 13574 16660 13626
rect 16684 13574 16698 13626
rect 16698 13574 16710 13626
rect 16710 13574 16740 13626
rect 16764 13574 16774 13626
rect 16774 13574 16820 13626
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16764 13572 16820 13574
rect 16302 12008 16358 12064
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16764 12538 16820 12540
rect 16524 12486 16570 12538
rect 16570 12486 16580 12538
rect 16604 12486 16634 12538
rect 16634 12486 16646 12538
rect 16646 12486 16660 12538
rect 16684 12486 16698 12538
rect 16698 12486 16710 12538
rect 16710 12486 16740 12538
rect 16764 12486 16774 12538
rect 16774 12486 16820 12538
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 16764 12484 16820 12486
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16764 11450 16820 11452
rect 16524 11398 16570 11450
rect 16570 11398 16580 11450
rect 16604 11398 16634 11450
rect 16634 11398 16646 11450
rect 16646 11398 16660 11450
rect 16684 11398 16698 11450
rect 16698 11398 16710 11450
rect 16710 11398 16740 11450
rect 16764 11398 16774 11450
rect 16774 11398 16820 11450
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16764 11396 16820 11398
rect 16486 11056 16542 11112
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16764 10362 16820 10364
rect 16524 10310 16570 10362
rect 16570 10310 16580 10362
rect 16604 10310 16634 10362
rect 16634 10310 16646 10362
rect 16646 10310 16660 10362
rect 16684 10310 16698 10362
rect 16698 10310 16710 10362
rect 16710 10310 16740 10362
rect 16764 10310 16774 10362
rect 16774 10310 16820 10362
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16764 10308 16820 10310
rect 16394 9424 16450 9480
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16764 9274 16820 9276
rect 16524 9222 16570 9274
rect 16570 9222 16580 9274
rect 16604 9222 16634 9274
rect 16634 9222 16646 9274
rect 16646 9222 16660 9274
rect 16684 9222 16698 9274
rect 16698 9222 16710 9274
rect 16710 9222 16740 9274
rect 16764 9222 16774 9274
rect 16774 9222 16820 9274
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16764 9220 16820 9222
rect 16302 8744 16358 8800
rect 16026 6840 16082 6896
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16764 8186 16820 8188
rect 16524 8134 16570 8186
rect 16570 8134 16580 8186
rect 16604 8134 16634 8186
rect 16634 8134 16646 8186
rect 16646 8134 16660 8186
rect 16684 8134 16698 8186
rect 16698 8134 16710 8186
rect 16710 8134 16740 8186
rect 16764 8134 16774 8186
rect 16774 8134 16820 8186
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16764 8132 16820 8134
rect 16394 7284 16396 7304
rect 16396 7284 16448 7304
rect 16448 7284 16450 7304
rect 16394 7248 16450 7284
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16764 7098 16820 7100
rect 16524 7046 16570 7098
rect 16570 7046 16580 7098
rect 16604 7046 16634 7098
rect 16634 7046 16646 7098
rect 16646 7046 16660 7098
rect 16684 7046 16698 7098
rect 16698 7046 16710 7098
rect 16710 7046 16740 7098
rect 16764 7046 16774 7098
rect 16774 7046 16820 7098
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16764 7044 16820 7046
rect 18418 12144 18474 12200
rect 17498 10784 17554 10840
rect 17038 6740 17040 6760
rect 17040 6740 17092 6760
rect 17092 6740 17094 6760
rect 17038 6704 17094 6740
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16764 6010 16820 6012
rect 16524 5958 16570 6010
rect 16570 5958 16580 6010
rect 16604 5958 16634 6010
rect 16634 5958 16646 6010
rect 16646 5958 16660 6010
rect 16684 5958 16698 6010
rect 16698 5958 16710 6010
rect 16710 5958 16740 6010
rect 16764 5958 16774 6010
rect 16774 5958 16820 6010
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 16764 5956 16820 5958
rect 15842 4664 15898 4720
rect 15934 4564 15936 4584
rect 15936 4564 15988 4584
rect 15988 4564 15990 4584
rect 15934 4528 15990 4564
rect 15750 3732 15806 3768
rect 15750 3712 15752 3732
rect 15752 3712 15804 3732
rect 15804 3712 15806 3732
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16764 4922 16820 4924
rect 16524 4870 16570 4922
rect 16570 4870 16580 4922
rect 16604 4870 16634 4922
rect 16634 4870 16646 4922
rect 16646 4870 16660 4922
rect 16684 4870 16698 4922
rect 16698 4870 16710 4922
rect 16710 4870 16740 4922
rect 16764 4870 16774 4922
rect 16774 4870 16820 4922
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16764 4868 16820 4870
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16764 3834 16820 3836
rect 16524 3782 16570 3834
rect 16570 3782 16580 3834
rect 16604 3782 16634 3834
rect 16634 3782 16646 3834
rect 16646 3782 16660 3834
rect 16684 3782 16698 3834
rect 16698 3782 16710 3834
rect 16710 3782 16740 3834
rect 16764 3782 16774 3834
rect 16774 3782 16820 3834
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 16764 3780 16820 3782
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16764 2746 16820 2748
rect 16524 2694 16570 2746
rect 16570 2694 16580 2746
rect 16604 2694 16634 2746
rect 16634 2694 16646 2746
rect 16646 2694 16660 2746
rect 16684 2694 16698 2746
rect 16698 2694 16710 2746
rect 16710 2694 16740 2746
rect 16764 2694 16774 2746
rect 16774 2694 16820 2746
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16764 2692 16820 2694
rect 17682 9580 17738 9616
rect 17682 9560 17684 9580
rect 17684 9560 17736 9580
rect 17736 9560 17738 9580
rect 17498 9152 17554 9208
rect 17498 6840 17554 6896
rect 17222 4256 17278 4312
rect 17590 5616 17646 5672
rect 17498 5208 17554 5264
rect 17314 3576 17370 3632
rect 16854 1400 16910 1456
rect 18050 8336 18106 8392
rect 18142 7520 18198 7576
rect 18050 7148 18052 7168
rect 18052 7148 18104 7168
rect 18104 7148 18106 7168
rect 18050 7112 18106 7148
rect 18050 6296 18106 6352
rect 17774 5888 17830 5944
rect 18234 5072 18290 5128
rect 17958 4664 18014 4720
rect 17958 3884 17960 3904
rect 17960 3884 18012 3904
rect 18012 3884 18014 3904
rect 17958 3848 18014 3884
rect 17774 3032 17830 3088
rect 17682 992 17738 1048
rect 18510 9968 18566 10024
rect 18418 7928 18474 7984
rect 18418 6704 18474 6760
rect 18418 5516 18420 5536
rect 18420 5516 18472 5536
rect 18472 5516 18474 5536
rect 18418 5480 18474 5516
rect 18326 2624 18382 2680
rect 18050 2252 18052 2272
rect 18052 2252 18104 2272
rect 18104 2252 18106 2272
rect 18050 2216 18106 2252
rect 18602 3440 18658 3496
rect 18510 1808 18566 1864
rect 16394 584 16450 640
<< metal3 >>
rect 0 16690 800 16720
rect 0 16630 2790 16690
rect 0 16600 800 16630
rect 2730 16418 2790 16630
rect 15469 16554 15535 16557
rect 19200 16554 20000 16584
rect 15469 16552 20000 16554
rect 15469 16496 15474 16552
rect 15530 16496 20000 16552
rect 15469 16494 20000 16496
rect 15469 16491 15535 16494
rect 19200 16464 20000 16494
rect 3049 16418 3115 16421
rect 2730 16416 3115 16418
rect 2730 16360 3054 16416
rect 3110 16360 3115 16416
rect 2730 16358 3115 16360
rect 3049 16355 3115 16358
rect 0 16282 800 16312
rect 2773 16282 2839 16285
rect 0 16280 2839 16282
rect 0 16224 2778 16280
rect 2834 16224 2839 16280
rect 0 16222 2839 16224
rect 0 16192 800 16222
rect 2773 16219 2839 16222
rect 16205 16146 16271 16149
rect 19200 16146 20000 16176
rect 16205 16144 20000 16146
rect 16205 16088 16210 16144
rect 16266 16088 20000 16144
rect 16205 16086 20000 16088
rect 16205 16083 16271 16086
rect 19200 16056 20000 16086
rect 0 15874 800 15904
rect 3969 15874 4035 15877
rect 0 15872 4035 15874
rect 0 15816 3974 15872
rect 4030 15816 4035 15872
rect 0 15814 4035 15816
rect 0 15784 800 15814
rect 3969 15811 4035 15814
rect 15285 15738 15351 15741
rect 19200 15738 20000 15768
rect 15285 15736 20000 15738
rect 15285 15680 15290 15736
rect 15346 15680 20000 15736
rect 15285 15678 20000 15680
rect 15285 15675 15351 15678
rect 19200 15648 20000 15678
rect 0 15466 800 15496
rect 3785 15466 3851 15469
rect 0 15464 3851 15466
rect 0 15408 3790 15464
rect 3846 15408 3851 15464
rect 0 15406 3851 15408
rect 0 15376 800 15406
rect 3785 15403 3851 15406
rect 17125 15330 17191 15333
rect 19200 15330 20000 15360
rect 17125 15328 20000 15330
rect 17125 15272 17130 15328
rect 17186 15272 20000 15328
rect 17125 15270 20000 15272
rect 17125 15267 17191 15270
rect 19200 15240 20000 15270
rect 0 15058 800 15088
rect 3601 15058 3667 15061
rect 0 15056 3667 15058
rect 0 15000 3606 15056
rect 3662 15000 3667 15056
rect 0 14998 3667 15000
rect 0 14968 800 14998
rect 3601 14995 3667 14998
rect 16021 14922 16087 14925
rect 19200 14922 20000 14952
rect 16021 14920 20000 14922
rect 16021 14864 16026 14920
rect 16082 14864 20000 14920
rect 16021 14862 20000 14864
rect 16021 14859 16087 14862
rect 19200 14832 20000 14862
rect 3170 14720 3486 14721
rect 0 14650 800 14680
rect 3170 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3486 14720
rect 3170 14655 3486 14656
rect 7618 14720 7934 14721
rect 7618 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7934 14720
rect 7618 14655 7934 14656
rect 12066 14720 12382 14721
rect 12066 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12382 14720
rect 12066 14655 12382 14656
rect 16514 14720 16830 14721
rect 16514 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16830 14720
rect 16514 14655 16830 14656
rect 2957 14650 3023 14653
rect 0 14648 3023 14650
rect 0 14592 2962 14648
rect 3018 14592 3023 14648
rect 0 14590 3023 14592
rect 0 14560 800 14590
rect 2957 14587 3023 14590
rect 16113 14514 16179 14517
rect 19200 14514 20000 14544
rect 16113 14512 20000 14514
rect 16113 14456 16118 14512
rect 16174 14456 20000 14512
rect 16113 14454 20000 14456
rect 16113 14451 16179 14454
rect 19200 14424 20000 14454
rect 4153 14378 4219 14381
rect 12617 14378 12683 14381
rect 4153 14376 12683 14378
rect 4153 14320 4158 14376
rect 4214 14320 12622 14376
rect 12678 14320 12683 14376
rect 4153 14318 12683 14320
rect 4153 14315 4219 14318
rect 12617 14315 12683 14318
rect 0 14242 800 14272
rect 4061 14242 4127 14245
rect 0 14240 4127 14242
rect 0 14184 4066 14240
rect 4122 14184 4127 14240
rect 0 14182 4127 14184
rect 0 14152 800 14182
rect 4061 14179 4127 14182
rect 5394 14176 5710 14177
rect 5394 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5710 14176
rect 5394 14111 5710 14112
rect 9842 14176 10158 14177
rect 9842 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10158 14176
rect 9842 14111 10158 14112
rect 14290 14176 14606 14177
rect 14290 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14606 14176
rect 14290 14111 14606 14112
rect 15837 14106 15903 14109
rect 19200 14106 20000 14136
rect 15837 14104 20000 14106
rect 15837 14048 15842 14104
rect 15898 14048 20000 14104
rect 15837 14046 20000 14048
rect 15837 14043 15903 14046
rect 19200 14016 20000 14046
rect 8845 13970 8911 13973
rect 9438 13970 9444 13972
rect 8845 13968 9444 13970
rect 8845 13912 8850 13968
rect 8906 13912 9444 13968
rect 8845 13910 9444 13912
rect 8845 13907 8911 13910
rect 9438 13908 9444 13910
rect 9508 13908 9514 13972
rect 0 13834 800 13864
rect 2129 13834 2195 13837
rect 0 13832 2195 13834
rect 0 13776 2134 13832
rect 2190 13776 2195 13832
rect 0 13774 2195 13776
rect 0 13744 800 13774
rect 2129 13771 2195 13774
rect 8886 13772 8892 13836
rect 8956 13834 8962 13836
rect 9121 13834 9187 13837
rect 8956 13832 9187 13834
rect 8956 13776 9126 13832
rect 9182 13776 9187 13832
rect 8956 13774 9187 13776
rect 8956 13772 8962 13774
rect 9121 13771 9187 13774
rect 13813 13698 13879 13701
rect 14958 13698 14964 13700
rect 13813 13696 14964 13698
rect 13813 13640 13818 13696
rect 13874 13640 14964 13696
rect 13813 13638 14964 13640
rect 13813 13635 13879 13638
rect 14958 13636 14964 13638
rect 15028 13636 15034 13700
rect 19200 13698 20000 13728
rect 16990 13638 20000 13698
rect 3170 13632 3486 13633
rect 3170 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3486 13632
rect 3170 13567 3486 13568
rect 7618 13632 7934 13633
rect 7618 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7934 13632
rect 7618 13567 7934 13568
rect 12066 13632 12382 13633
rect 12066 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12382 13632
rect 12066 13567 12382 13568
rect 16514 13632 16830 13633
rect 16514 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16830 13632
rect 16514 13567 16830 13568
rect 0 13426 800 13456
rect 4061 13426 4127 13429
rect 0 13424 4127 13426
rect 0 13368 4066 13424
rect 4122 13368 4127 13424
rect 0 13366 4127 13368
rect 0 13336 800 13366
rect 4061 13363 4127 13366
rect 5257 13426 5323 13429
rect 15009 13426 15075 13429
rect 5257 13424 15075 13426
rect 5257 13368 5262 13424
rect 5318 13368 15014 13424
rect 15070 13368 15075 13424
rect 5257 13366 15075 13368
rect 5257 13363 5323 13366
rect 15009 13363 15075 13366
rect 15929 13426 15995 13429
rect 16990 13426 17050 13638
rect 19200 13608 20000 13638
rect 15929 13424 17050 13426
rect 15929 13368 15934 13424
rect 15990 13368 17050 13424
rect 15929 13366 17050 13368
rect 15929 13363 15995 13366
rect 15193 13290 15259 13293
rect 19200 13290 20000 13320
rect 15193 13288 20000 13290
rect 15193 13232 15198 13288
rect 15254 13232 20000 13288
rect 15193 13230 20000 13232
rect 15193 13227 15259 13230
rect 19200 13200 20000 13230
rect 5394 13088 5710 13089
rect 0 13018 800 13048
rect 5394 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5710 13088
rect 5394 13023 5710 13024
rect 9842 13088 10158 13089
rect 9842 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10158 13088
rect 9842 13023 10158 13024
rect 14290 13088 14606 13089
rect 14290 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14606 13088
rect 14290 13023 14606 13024
rect 1342 13018 1348 13020
rect 0 12958 1348 13018
rect 0 12928 800 12958
rect 1342 12956 1348 12958
rect 1412 12956 1418 13020
rect 3877 12884 3943 12885
rect 3877 12880 3924 12884
rect 3988 12882 3994 12884
rect 15837 12882 15903 12885
rect 19200 12882 20000 12912
rect 3877 12824 3882 12880
rect 3877 12820 3924 12824
rect 3988 12822 4034 12882
rect 15837 12880 20000 12882
rect 15837 12824 15842 12880
rect 15898 12824 20000 12880
rect 15837 12822 20000 12824
rect 3988 12820 3994 12822
rect 3877 12819 3943 12820
rect 15837 12819 15903 12822
rect 19200 12792 20000 12822
rect 3693 12746 3759 12749
rect 2730 12744 3759 12746
rect 2730 12688 3698 12744
rect 3754 12688 3759 12744
rect 2730 12686 3759 12688
rect 0 12610 800 12640
rect 2730 12610 2790 12686
rect 3693 12683 3759 12686
rect 10501 12746 10567 12749
rect 14273 12746 14339 12749
rect 10501 12744 14339 12746
rect 10501 12688 10506 12744
rect 10562 12688 14278 12744
rect 14334 12688 14339 12744
rect 10501 12686 14339 12688
rect 10501 12683 10567 12686
rect 14273 12683 14339 12686
rect 15150 12686 17050 12746
rect 0 12550 2790 12610
rect 0 12520 800 12550
rect 3170 12544 3486 12545
rect 3170 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3486 12544
rect 3170 12479 3486 12480
rect 7618 12544 7934 12545
rect 7618 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7934 12544
rect 7618 12479 7934 12480
rect 12066 12544 12382 12545
rect 12066 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12382 12544
rect 12066 12479 12382 12480
rect 9765 12338 9831 12341
rect 15150 12338 15210 12686
rect 16514 12544 16830 12545
rect 16514 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16830 12544
rect 16514 12479 16830 12480
rect 16990 12474 17050 12686
rect 19200 12474 20000 12504
rect 16990 12414 20000 12474
rect 19200 12384 20000 12414
rect 9765 12336 15210 12338
rect 9765 12280 9770 12336
rect 9826 12280 15210 12336
rect 9765 12278 15210 12280
rect 9765 12275 9831 12278
rect 0 12202 800 12232
rect 4102 12202 4108 12204
rect 0 12142 4108 12202
rect 0 12112 800 12142
rect 4102 12140 4108 12142
rect 4172 12140 4178 12204
rect 13169 12202 13235 12205
rect 18413 12202 18479 12205
rect 13169 12200 18479 12202
rect 13169 12144 13174 12200
rect 13230 12144 18418 12200
rect 18474 12144 18479 12200
rect 13169 12142 18479 12144
rect 13169 12139 13235 12142
rect 18413 12139 18479 12142
rect 16297 12066 16363 12069
rect 19200 12066 20000 12096
rect 16297 12064 20000 12066
rect 16297 12008 16302 12064
rect 16358 12008 20000 12064
rect 16297 12006 20000 12008
rect 16297 12003 16363 12006
rect 5394 12000 5710 12001
rect 5394 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5710 12000
rect 5394 11935 5710 11936
rect 9842 12000 10158 12001
rect 9842 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10158 12000
rect 9842 11935 10158 11936
rect 14290 12000 14606 12001
rect 14290 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14606 12000
rect 19200 11976 20000 12006
rect 14290 11935 14606 11936
rect 0 11794 800 11824
rect 4061 11794 4127 11797
rect 0 11792 4127 11794
rect 0 11736 4066 11792
rect 4122 11736 4127 11792
rect 0 11734 4127 11736
rect 0 11704 800 11734
rect 4061 11731 4127 11734
rect 6453 11658 6519 11661
rect 12801 11658 12867 11661
rect 19200 11658 20000 11688
rect 6453 11656 20000 11658
rect 6453 11600 6458 11656
rect 6514 11600 12806 11656
rect 12862 11600 20000 11656
rect 6453 11598 20000 11600
rect 6453 11595 6519 11598
rect 12801 11595 12867 11598
rect 19200 11568 20000 11598
rect 3170 11456 3486 11457
rect 0 11386 800 11416
rect 3170 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3486 11456
rect 3170 11391 3486 11392
rect 7618 11456 7934 11457
rect 7618 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7934 11456
rect 7618 11391 7934 11392
rect 12066 11456 12382 11457
rect 12066 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12382 11456
rect 12066 11391 12382 11392
rect 16514 11456 16830 11457
rect 16514 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16830 11456
rect 16514 11391 16830 11392
rect 0 11326 2100 11386
rect 0 11296 800 11326
rect 2040 11250 2100 11326
rect 3601 11250 3667 11253
rect 8569 11250 8635 11253
rect 2040 11190 2790 11250
rect 2730 11114 2790 11190
rect 3601 11248 8635 11250
rect 3601 11192 3606 11248
rect 3662 11192 8574 11248
rect 8630 11192 8635 11248
rect 3601 11190 8635 11192
rect 3601 11187 3667 11190
rect 8569 11187 8635 11190
rect 15285 11250 15351 11253
rect 19200 11250 20000 11280
rect 15285 11248 20000 11250
rect 15285 11192 15290 11248
rect 15346 11192 20000 11248
rect 15285 11190 20000 11192
rect 15285 11187 15351 11190
rect 19200 11160 20000 11190
rect 3601 11114 3667 11117
rect 2730 11112 3667 11114
rect 2730 11056 3606 11112
rect 3662 11056 3667 11112
rect 2730 11054 3667 11056
rect 3601 11051 3667 11054
rect 10501 11114 10567 11117
rect 16481 11114 16547 11117
rect 10501 11112 16547 11114
rect 10501 11056 10506 11112
rect 10562 11056 16486 11112
rect 16542 11056 16547 11112
rect 10501 11054 16547 11056
rect 10501 11051 10567 11054
rect 16481 11051 16547 11054
rect 0 10978 800 11008
rect 4061 10978 4127 10981
rect 0 10976 4127 10978
rect 0 10920 4066 10976
rect 4122 10920 4127 10976
rect 0 10918 4127 10920
rect 0 10888 800 10918
rect 4061 10915 4127 10918
rect 5394 10912 5710 10913
rect 5394 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5710 10912
rect 5394 10847 5710 10848
rect 9842 10912 10158 10913
rect 9842 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10158 10912
rect 9842 10847 10158 10848
rect 14290 10912 14606 10913
rect 14290 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14606 10912
rect 14290 10847 14606 10848
rect 17493 10842 17559 10845
rect 19200 10842 20000 10872
rect 17493 10840 20000 10842
rect 17493 10784 17498 10840
rect 17554 10784 20000 10840
rect 17493 10782 20000 10784
rect 17493 10779 17559 10782
rect 19200 10752 20000 10782
rect 2681 10706 2747 10709
rect 13813 10706 13879 10709
rect 2681 10704 13879 10706
rect 2681 10648 2686 10704
rect 2742 10648 13818 10704
rect 13874 10648 13879 10704
rect 2681 10646 13879 10648
rect 2681 10643 2747 10646
rect 13813 10643 13879 10646
rect 0 10570 800 10600
rect 1577 10570 1643 10573
rect 0 10568 1643 10570
rect 0 10512 1582 10568
rect 1638 10512 1643 10568
rect 0 10510 1643 10512
rect 0 10480 800 10510
rect 1577 10507 1643 10510
rect 3877 10570 3943 10573
rect 14457 10570 14523 10573
rect 3877 10568 14523 10570
rect 3877 10512 3882 10568
rect 3938 10512 14462 10568
rect 14518 10512 14523 10568
rect 3877 10510 14523 10512
rect 3877 10507 3943 10510
rect 14457 10507 14523 10510
rect 19200 10434 20000 10464
rect 16990 10374 20000 10434
rect 3170 10368 3486 10369
rect 3170 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3486 10368
rect 3170 10303 3486 10304
rect 7618 10368 7934 10369
rect 7618 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7934 10368
rect 7618 10303 7934 10304
rect 12066 10368 12382 10369
rect 12066 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12382 10368
rect 12066 10303 12382 10304
rect 16514 10368 16830 10369
rect 16514 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16830 10368
rect 16514 10303 16830 10304
rect 0 10162 800 10192
rect 4061 10162 4127 10165
rect 0 10160 4127 10162
rect 0 10104 4066 10160
rect 4122 10104 4127 10160
rect 0 10102 4127 10104
rect 0 10072 800 10102
rect 4061 10099 4127 10102
rect 15929 10162 15995 10165
rect 16990 10162 17050 10374
rect 19200 10344 20000 10374
rect 15929 10160 17050 10162
rect 15929 10104 15934 10160
rect 15990 10104 17050 10160
rect 15929 10102 17050 10104
rect 15929 10099 15995 10102
rect 18505 10026 18571 10029
rect 19200 10026 20000 10056
rect 18505 10024 20000 10026
rect 18505 9968 18510 10024
rect 18566 9968 20000 10024
rect 18505 9966 20000 9968
rect 18505 9963 18571 9966
rect 19200 9936 20000 9966
rect 5394 9824 5710 9825
rect 0 9754 800 9784
rect 5394 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5710 9824
rect 5394 9759 5710 9760
rect 9842 9824 10158 9825
rect 9842 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10158 9824
rect 9842 9759 10158 9760
rect 14290 9824 14606 9825
rect 14290 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14606 9824
rect 14290 9759 14606 9760
rect 4337 9754 4403 9757
rect 0 9752 4403 9754
rect 0 9696 4342 9752
rect 4398 9696 4403 9752
rect 0 9694 4403 9696
rect 0 9664 800 9694
rect 4337 9691 4403 9694
rect 3918 9556 3924 9620
rect 3988 9618 3994 9620
rect 17677 9618 17743 9621
rect 19200 9618 20000 9648
rect 3988 9616 17743 9618
rect 3988 9560 17682 9616
rect 17738 9560 17743 9616
rect 3988 9558 17743 9560
rect 3988 9556 3994 9558
rect 17677 9555 17743 9558
rect 17910 9558 20000 9618
rect 4061 9482 4127 9485
rect 2730 9480 4127 9482
rect 2730 9424 4066 9480
rect 4122 9424 4127 9480
rect 2730 9422 4127 9424
rect 0 9346 800 9376
rect 2730 9346 2790 9422
rect 4061 9419 4127 9422
rect 16389 9482 16455 9485
rect 17910 9482 17970 9558
rect 19200 9528 20000 9558
rect 16389 9480 17970 9482
rect 16389 9424 16394 9480
rect 16450 9424 17970 9480
rect 16389 9422 17970 9424
rect 16389 9419 16455 9422
rect 0 9286 2790 9346
rect 0 9256 800 9286
rect 3170 9280 3486 9281
rect 3170 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3486 9280
rect 3170 9215 3486 9216
rect 7618 9280 7934 9281
rect 7618 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7934 9280
rect 7618 9215 7934 9216
rect 12066 9280 12382 9281
rect 12066 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12382 9280
rect 12066 9215 12382 9216
rect 16514 9280 16830 9281
rect 16514 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16830 9280
rect 16514 9215 16830 9216
rect 17493 9210 17559 9213
rect 19200 9210 20000 9240
rect 17493 9208 20000 9210
rect 17493 9152 17498 9208
rect 17554 9152 20000 9208
rect 17493 9150 20000 9152
rect 17493 9147 17559 9150
rect 19200 9120 20000 9150
rect 4102 9012 4108 9076
rect 4172 9074 4178 9076
rect 7557 9074 7623 9077
rect 4172 9072 7623 9074
rect 4172 9016 7562 9072
rect 7618 9016 7623 9072
rect 4172 9014 7623 9016
rect 4172 9012 4178 9014
rect 7557 9011 7623 9014
rect 0 8938 800 8968
rect 1669 8938 1735 8941
rect 0 8936 1735 8938
rect 0 8880 1674 8936
rect 1730 8880 1735 8936
rect 0 8878 1735 8880
rect 0 8848 800 8878
rect 1669 8875 1735 8878
rect 2630 8740 2636 8804
rect 2700 8802 2706 8804
rect 2957 8802 3023 8805
rect 2700 8800 3023 8802
rect 2700 8744 2962 8800
rect 3018 8744 3023 8800
rect 2700 8742 3023 8744
rect 2700 8740 2706 8742
rect 2957 8739 3023 8742
rect 16297 8802 16363 8805
rect 19200 8802 20000 8832
rect 16297 8800 20000 8802
rect 16297 8744 16302 8800
rect 16358 8744 20000 8800
rect 16297 8742 20000 8744
rect 16297 8739 16363 8742
rect 5394 8736 5710 8737
rect 5394 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5710 8736
rect 5394 8671 5710 8672
rect 9842 8736 10158 8737
rect 9842 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10158 8736
rect 9842 8671 10158 8672
rect 14290 8736 14606 8737
rect 14290 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14606 8736
rect 19200 8712 20000 8742
rect 14290 8671 14606 8672
rect 0 8530 800 8560
rect 2773 8530 2839 8533
rect 0 8528 2839 8530
rect 0 8472 2778 8528
rect 2834 8472 2839 8528
rect 0 8470 2839 8472
rect 0 8440 800 8470
rect 2773 8467 2839 8470
rect 18045 8394 18111 8397
rect 19200 8394 20000 8424
rect 18045 8392 20000 8394
rect 18045 8336 18050 8392
rect 18106 8336 20000 8392
rect 18045 8334 20000 8336
rect 18045 8331 18111 8334
rect 19200 8304 20000 8334
rect 1342 8196 1348 8260
rect 1412 8258 1418 8260
rect 1485 8258 1551 8261
rect 1412 8256 1551 8258
rect 1412 8200 1490 8256
rect 1546 8200 1551 8256
rect 1412 8198 1551 8200
rect 1412 8196 1418 8198
rect 1485 8195 1551 8198
rect 3170 8192 3486 8193
rect 0 8122 800 8152
rect 3170 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3486 8192
rect 3170 8127 3486 8128
rect 7618 8192 7934 8193
rect 7618 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7934 8192
rect 7618 8127 7934 8128
rect 12066 8192 12382 8193
rect 12066 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12382 8192
rect 12066 8127 12382 8128
rect 16514 8192 16830 8193
rect 16514 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16830 8192
rect 16514 8127 16830 8128
rect 1393 8122 1459 8125
rect 0 8120 1459 8122
rect 0 8064 1398 8120
rect 1454 8064 1459 8120
rect 0 8062 1459 8064
rect 0 8032 800 8062
rect 1393 8059 1459 8062
rect 18413 7986 18479 7989
rect 19200 7986 20000 8016
rect 18413 7984 20000 7986
rect 18413 7928 18418 7984
rect 18474 7928 20000 7984
rect 18413 7926 20000 7928
rect 18413 7923 18479 7926
rect 19200 7896 20000 7926
rect 2773 7850 2839 7853
rect 2773 7848 12450 7850
rect 2773 7792 2778 7848
rect 2834 7792 12450 7848
rect 2773 7790 12450 7792
rect 2773 7787 2839 7790
rect 0 7714 800 7744
rect 3785 7714 3851 7717
rect 0 7712 3851 7714
rect 0 7656 3790 7712
rect 3846 7656 3851 7712
rect 0 7654 3851 7656
rect 0 7624 800 7654
rect 3785 7651 3851 7654
rect 5394 7648 5710 7649
rect 5394 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5710 7648
rect 5394 7583 5710 7584
rect 9842 7648 10158 7649
rect 9842 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10158 7648
rect 9842 7583 10158 7584
rect 0 7306 800 7336
rect 1577 7306 1643 7309
rect 0 7304 1643 7306
rect 0 7248 1582 7304
rect 1638 7248 1643 7304
rect 0 7246 1643 7248
rect 12390 7306 12450 7790
rect 14290 7648 14606 7649
rect 14290 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14606 7648
rect 14290 7583 14606 7584
rect 18137 7578 18203 7581
rect 19200 7578 20000 7608
rect 18137 7576 20000 7578
rect 18137 7520 18142 7576
rect 18198 7520 20000 7576
rect 18137 7518 20000 7520
rect 18137 7515 18203 7518
rect 19200 7488 20000 7518
rect 16389 7306 16455 7309
rect 12390 7304 16455 7306
rect 12390 7248 16394 7304
rect 16450 7248 16455 7304
rect 12390 7246 16455 7248
rect 0 7216 800 7246
rect 1577 7243 1643 7246
rect 16389 7243 16455 7246
rect 18045 7170 18111 7173
rect 19200 7170 20000 7200
rect 18045 7168 20000 7170
rect 18045 7112 18050 7168
rect 18106 7112 20000 7168
rect 18045 7110 20000 7112
rect 18045 7107 18111 7110
rect 3170 7104 3486 7105
rect 3170 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3486 7104
rect 3170 7039 3486 7040
rect 7618 7104 7934 7105
rect 7618 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7934 7104
rect 7618 7039 7934 7040
rect 12066 7104 12382 7105
rect 12066 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12382 7104
rect 12066 7039 12382 7040
rect 16514 7104 16830 7105
rect 16514 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16830 7104
rect 19200 7080 20000 7110
rect 16514 7039 16830 7040
rect 0 6898 800 6928
rect 2037 6898 2103 6901
rect 0 6896 2103 6898
rect 0 6840 2042 6896
rect 2098 6840 2103 6896
rect 0 6838 2103 6840
rect 0 6808 800 6838
rect 2037 6835 2103 6838
rect 15377 6898 15443 6901
rect 16021 6898 16087 6901
rect 17493 6898 17559 6901
rect 15377 6896 17559 6898
rect 15377 6840 15382 6896
rect 15438 6840 16026 6896
rect 16082 6840 17498 6896
rect 17554 6840 17559 6896
rect 15377 6838 17559 6840
rect 15377 6835 15443 6838
rect 16021 6835 16087 6838
rect 17493 6835 17559 6838
rect 1945 6762 2011 6765
rect 2630 6762 2636 6764
rect 1945 6760 2636 6762
rect 1945 6704 1950 6760
rect 2006 6704 2636 6760
rect 1945 6702 2636 6704
rect 1945 6699 2011 6702
rect 2630 6700 2636 6702
rect 2700 6762 2706 6764
rect 17033 6762 17099 6765
rect 2700 6760 17099 6762
rect 2700 6704 17038 6760
rect 17094 6704 17099 6760
rect 2700 6702 17099 6704
rect 2700 6700 2706 6702
rect 17033 6699 17099 6702
rect 18413 6762 18479 6765
rect 19200 6762 20000 6792
rect 18413 6760 20000 6762
rect 18413 6704 18418 6760
rect 18474 6704 20000 6760
rect 18413 6702 20000 6704
rect 18413 6699 18479 6702
rect 19200 6672 20000 6702
rect 5394 6560 5710 6561
rect 0 6490 800 6520
rect 5394 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5710 6560
rect 5394 6495 5710 6496
rect 9842 6560 10158 6561
rect 9842 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10158 6560
rect 9842 6495 10158 6496
rect 14290 6560 14606 6561
rect 14290 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14606 6560
rect 14290 6495 14606 6496
rect 1577 6490 1643 6493
rect 0 6488 1643 6490
rect 0 6432 1582 6488
rect 1638 6432 1643 6488
rect 0 6430 1643 6432
rect 0 6400 800 6430
rect 1577 6427 1643 6430
rect 3785 6490 3851 6493
rect 3785 6488 3986 6490
rect 3785 6432 3790 6488
rect 3846 6432 3986 6488
rect 3785 6430 3986 6432
rect 3785 6427 3851 6430
rect 3693 6218 3759 6221
rect 1902 6216 3759 6218
rect 1902 6160 3698 6216
rect 3754 6160 3759 6216
rect 1902 6158 3759 6160
rect 0 6082 800 6112
rect 1902 6082 1962 6158
rect 3693 6155 3759 6158
rect 0 6022 1962 6082
rect 0 5992 800 6022
rect 3170 6016 3486 6017
rect 3170 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3486 6016
rect 3170 5951 3486 5952
rect 3926 5813 3986 6430
rect 18045 6354 18111 6357
rect 19200 6354 20000 6384
rect 18045 6352 20000 6354
rect 18045 6296 18050 6352
rect 18106 6296 20000 6352
rect 18045 6294 20000 6296
rect 18045 6291 18111 6294
rect 19200 6264 20000 6294
rect 6545 6218 6611 6221
rect 15377 6218 15443 6221
rect 6545 6216 15443 6218
rect 6545 6160 6550 6216
rect 6606 6160 15382 6216
rect 15438 6160 15443 6216
rect 6545 6158 15443 6160
rect 6545 6155 6611 6158
rect 15377 6155 15443 6158
rect 7618 6016 7934 6017
rect 7618 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7934 6016
rect 7618 5951 7934 5952
rect 12066 6016 12382 6017
rect 12066 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12382 6016
rect 12066 5951 12382 5952
rect 16514 6016 16830 6017
rect 16514 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16830 6016
rect 16514 5951 16830 5952
rect 17769 5946 17835 5949
rect 19200 5946 20000 5976
rect 17769 5944 20000 5946
rect 17769 5888 17774 5944
rect 17830 5888 20000 5944
rect 17769 5886 20000 5888
rect 17769 5883 17835 5886
rect 19200 5856 20000 5886
rect 3877 5808 3986 5813
rect 3877 5752 3882 5808
rect 3938 5752 3986 5808
rect 3877 5750 3986 5752
rect 3877 5747 3943 5750
rect 0 5674 800 5704
rect 2865 5674 2931 5677
rect 0 5672 2931 5674
rect 0 5616 2870 5672
rect 2926 5616 2931 5672
rect 0 5614 2931 5616
rect 0 5584 800 5614
rect 2865 5611 2931 5614
rect 14733 5674 14799 5677
rect 17585 5674 17651 5677
rect 14733 5672 17651 5674
rect 14733 5616 14738 5672
rect 14794 5616 17590 5672
rect 17646 5616 17651 5672
rect 14733 5614 17651 5616
rect 14733 5611 14799 5614
rect 17585 5611 17651 5614
rect 18413 5538 18479 5541
rect 19200 5538 20000 5568
rect 18413 5536 20000 5538
rect 18413 5480 18418 5536
rect 18474 5480 20000 5536
rect 18413 5478 20000 5480
rect 18413 5475 18479 5478
rect 5394 5472 5710 5473
rect 5394 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5710 5472
rect 5394 5407 5710 5408
rect 9842 5472 10158 5473
rect 9842 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10158 5472
rect 9842 5407 10158 5408
rect 14290 5472 14606 5473
rect 14290 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14606 5472
rect 19200 5448 20000 5478
rect 14290 5407 14606 5408
rect 3049 5402 3115 5405
rect 1902 5400 3115 5402
rect 1902 5344 3054 5400
rect 3110 5344 3115 5400
rect 1902 5342 3115 5344
rect 0 5266 800 5296
rect 1902 5266 1962 5342
rect 3049 5339 3115 5342
rect 0 5206 1962 5266
rect 2405 5266 2471 5269
rect 13537 5266 13603 5269
rect 2405 5264 13603 5266
rect 2405 5208 2410 5264
rect 2466 5208 13542 5264
rect 13598 5208 13603 5264
rect 2405 5206 13603 5208
rect 0 5176 800 5206
rect 2405 5203 2471 5206
rect 13537 5203 13603 5206
rect 13721 5266 13787 5269
rect 17493 5266 17559 5269
rect 13721 5264 17559 5266
rect 13721 5208 13726 5264
rect 13782 5208 17498 5264
rect 17554 5208 17559 5264
rect 13721 5206 17559 5208
rect 13721 5203 13787 5206
rect 17493 5203 17559 5206
rect 3785 5130 3851 5133
rect 14089 5130 14155 5133
rect 3785 5128 14155 5130
rect 3785 5072 3790 5128
rect 3846 5072 14094 5128
rect 14150 5072 14155 5128
rect 3785 5070 14155 5072
rect 3785 5067 3851 5070
rect 14089 5067 14155 5070
rect 18229 5130 18295 5133
rect 19200 5130 20000 5160
rect 18229 5128 20000 5130
rect 18229 5072 18234 5128
rect 18290 5072 20000 5128
rect 18229 5070 20000 5072
rect 18229 5067 18295 5070
rect 19200 5040 20000 5070
rect 3170 4928 3486 4929
rect 0 4858 800 4888
rect 3170 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3486 4928
rect 3170 4863 3486 4864
rect 7618 4928 7934 4929
rect 7618 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7934 4928
rect 7618 4863 7934 4864
rect 12066 4928 12382 4929
rect 12066 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12382 4928
rect 12066 4863 12382 4864
rect 16514 4928 16830 4929
rect 16514 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16830 4928
rect 16514 4863 16830 4864
rect 2773 4858 2839 4861
rect 0 4856 2839 4858
rect 0 4800 2778 4856
rect 2834 4800 2839 4856
rect 0 4798 2839 4800
rect 0 4768 800 4798
rect 2773 4795 2839 4798
rect 4102 4796 4108 4860
rect 4172 4858 4178 4860
rect 5901 4858 5967 4861
rect 4172 4856 5967 4858
rect 4172 4800 5906 4856
rect 5962 4800 5967 4856
rect 4172 4798 5967 4800
rect 4172 4796 4178 4798
rect 5901 4795 5967 4798
rect 13537 4858 13603 4861
rect 15377 4858 15443 4861
rect 13537 4856 15443 4858
rect 13537 4800 13542 4856
rect 13598 4800 15382 4856
rect 15438 4800 15443 4856
rect 13537 4798 15443 4800
rect 13537 4795 13603 4798
rect 15377 4795 15443 4798
rect 3049 4722 3115 4725
rect 3969 4722 4035 4725
rect 7465 4722 7531 4725
rect 15837 4722 15903 4725
rect 3049 4720 15903 4722
rect 3049 4664 3054 4720
rect 3110 4664 3974 4720
rect 4030 4664 7470 4720
rect 7526 4664 15842 4720
rect 15898 4664 15903 4720
rect 3049 4662 15903 4664
rect 3049 4659 3115 4662
rect 3969 4659 4035 4662
rect 7465 4659 7531 4662
rect 15837 4659 15903 4662
rect 17953 4722 18019 4725
rect 19200 4722 20000 4752
rect 17953 4720 20000 4722
rect 17953 4664 17958 4720
rect 18014 4664 20000 4720
rect 17953 4662 20000 4664
rect 17953 4659 18019 4662
rect 19200 4632 20000 4662
rect 3877 4586 3943 4589
rect 15929 4586 15995 4589
rect 3877 4584 15995 4586
rect 3877 4528 3882 4584
rect 3938 4528 15934 4584
rect 15990 4528 15995 4584
rect 3877 4526 15995 4528
rect 3877 4523 3943 4526
rect 15929 4523 15995 4526
rect 0 4450 800 4480
rect 1485 4450 1551 4453
rect 0 4448 1551 4450
rect 0 4392 1490 4448
rect 1546 4392 1551 4448
rect 0 4390 1551 4392
rect 0 4360 800 4390
rect 1485 4387 1551 4390
rect 5394 4384 5710 4385
rect 5394 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5710 4384
rect 5394 4319 5710 4320
rect 9842 4384 10158 4385
rect 9842 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10158 4384
rect 9842 4319 10158 4320
rect 14290 4384 14606 4385
rect 14290 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14606 4384
rect 14290 4319 14606 4320
rect 17217 4314 17283 4317
rect 19200 4314 20000 4344
rect 17217 4312 20000 4314
rect 17217 4256 17222 4312
rect 17278 4256 20000 4312
rect 17217 4254 20000 4256
rect 17217 4251 17283 4254
rect 19200 4224 20000 4254
rect 3233 4178 3299 4181
rect 14733 4178 14799 4181
rect 3233 4176 14799 4178
rect 3233 4120 3238 4176
rect 3294 4120 14738 4176
rect 14794 4120 14799 4176
rect 3233 4118 14799 4120
rect 3233 4115 3299 4118
rect 14733 4115 14799 4118
rect 0 4042 800 4072
rect 2313 4042 2379 4045
rect 0 4040 2379 4042
rect 0 3984 2318 4040
rect 2374 3984 2379 4040
rect 0 3982 2379 3984
rect 0 3952 800 3982
rect 2313 3979 2379 3982
rect 8753 4042 8819 4045
rect 8886 4042 8892 4044
rect 8753 4040 8892 4042
rect 8753 3984 8758 4040
rect 8814 3984 8892 4040
rect 8753 3982 8892 3984
rect 8753 3979 8819 3982
rect 8886 3980 8892 3982
rect 8956 3980 8962 4044
rect 9305 4042 9371 4045
rect 9438 4042 9444 4044
rect 9305 4040 9444 4042
rect 9305 3984 9310 4040
rect 9366 3984 9444 4040
rect 9305 3982 9444 3984
rect 9305 3979 9371 3982
rect 9438 3980 9444 3982
rect 9508 3980 9514 4044
rect 9673 4042 9739 4045
rect 12525 4042 12591 4045
rect 9673 4040 12591 4042
rect 9673 3984 9678 4040
rect 9734 3984 12530 4040
rect 12586 3984 12591 4040
rect 9673 3982 12591 3984
rect 9673 3979 9739 3982
rect 12525 3979 12591 3982
rect 17953 3906 18019 3909
rect 19200 3906 20000 3936
rect 17953 3904 20000 3906
rect 17953 3848 17958 3904
rect 18014 3848 20000 3904
rect 17953 3846 20000 3848
rect 17953 3843 18019 3846
rect 3170 3840 3486 3841
rect 3170 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3486 3840
rect 3170 3775 3486 3776
rect 7618 3840 7934 3841
rect 7618 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7934 3840
rect 7618 3775 7934 3776
rect 12066 3840 12382 3841
rect 12066 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12382 3840
rect 12066 3775 12382 3776
rect 16514 3840 16830 3841
rect 16514 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16830 3840
rect 19200 3816 20000 3846
rect 16514 3775 16830 3776
rect 14958 3708 14964 3772
rect 15028 3770 15034 3772
rect 15745 3770 15811 3773
rect 15028 3768 15811 3770
rect 15028 3712 15750 3768
rect 15806 3712 15811 3768
rect 15028 3710 15811 3712
rect 15028 3708 15034 3710
rect 15745 3707 15811 3710
rect 0 3634 800 3664
rect 1577 3634 1643 3637
rect 0 3632 1643 3634
rect 0 3576 1582 3632
rect 1638 3576 1643 3632
rect 0 3574 1643 3576
rect 0 3544 800 3574
rect 1577 3571 1643 3574
rect 12617 3634 12683 3637
rect 17309 3634 17375 3637
rect 12617 3632 17375 3634
rect 12617 3576 12622 3632
rect 12678 3576 17314 3632
rect 17370 3576 17375 3632
rect 12617 3574 17375 3576
rect 12617 3571 12683 3574
rect 17309 3571 17375 3574
rect 2681 3498 2747 3501
rect 10501 3498 10567 3501
rect 2681 3496 10567 3498
rect 2681 3440 2686 3496
rect 2742 3440 10506 3496
rect 10562 3440 10567 3496
rect 2681 3438 10567 3440
rect 2681 3435 2747 3438
rect 10501 3435 10567 3438
rect 18597 3498 18663 3501
rect 19200 3498 20000 3528
rect 18597 3496 20000 3498
rect 18597 3440 18602 3496
rect 18658 3440 20000 3496
rect 18597 3438 20000 3440
rect 18597 3435 18663 3438
rect 19200 3408 20000 3438
rect 5394 3296 5710 3297
rect 0 3226 800 3256
rect 5394 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5710 3296
rect 5394 3231 5710 3232
rect 9842 3296 10158 3297
rect 9842 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10158 3296
rect 9842 3231 10158 3232
rect 14290 3296 14606 3297
rect 14290 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14606 3296
rect 14290 3231 14606 3232
rect 2221 3226 2287 3229
rect 0 3224 2287 3226
rect 0 3168 2226 3224
rect 2282 3168 2287 3224
rect 0 3166 2287 3168
rect 0 3136 800 3166
rect 2221 3163 2287 3166
rect 5073 3090 5139 3093
rect 13813 3090 13879 3093
rect 5073 3088 13879 3090
rect 5073 3032 5078 3088
rect 5134 3032 13818 3088
rect 13874 3032 13879 3088
rect 5073 3030 13879 3032
rect 5073 3027 5139 3030
rect 13813 3027 13879 3030
rect 17769 3090 17835 3093
rect 19200 3090 20000 3120
rect 17769 3088 20000 3090
rect 17769 3032 17774 3088
rect 17830 3032 20000 3088
rect 17769 3030 20000 3032
rect 17769 3027 17835 3030
rect 19200 3000 20000 3030
rect 7373 2954 7439 2957
rect 11145 2954 11211 2957
rect 12065 2954 12131 2957
rect 7373 2952 11211 2954
rect 7373 2896 7378 2952
rect 7434 2896 11150 2952
rect 11206 2896 11211 2952
rect 7373 2894 11211 2896
rect 7373 2891 7439 2894
rect 11145 2891 11211 2894
rect 11838 2952 12131 2954
rect 11838 2896 12070 2952
rect 12126 2896 12131 2952
rect 11838 2894 12131 2896
rect 0 2818 800 2848
rect 11838 2821 11898 2894
rect 12065 2891 12131 2894
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 11789 2816 11898 2821
rect 11789 2760 11794 2816
rect 11850 2760 11898 2816
rect 11789 2758 11898 2760
rect 11789 2755 11855 2758
rect 3170 2752 3486 2753
rect 3170 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3486 2752
rect 3170 2687 3486 2688
rect 7618 2752 7934 2753
rect 7618 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7934 2752
rect 7618 2687 7934 2688
rect 12066 2752 12382 2753
rect 12066 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12382 2752
rect 12066 2687 12382 2688
rect 16514 2752 16830 2753
rect 16514 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16830 2752
rect 16514 2687 16830 2688
rect 18321 2682 18387 2685
rect 19200 2682 20000 2712
rect 18321 2680 20000 2682
rect 18321 2624 18326 2680
rect 18382 2624 20000 2680
rect 18321 2622 20000 2624
rect 18321 2619 18387 2622
rect 19200 2592 20000 2622
rect 0 2410 800 2440
rect 2957 2410 3023 2413
rect 0 2408 3023 2410
rect 0 2352 2962 2408
rect 3018 2352 3023 2408
rect 0 2350 3023 2352
rect 0 2320 800 2350
rect 2957 2347 3023 2350
rect 18045 2274 18111 2277
rect 19200 2274 20000 2304
rect 18045 2272 20000 2274
rect 18045 2216 18050 2272
rect 18106 2216 20000 2272
rect 18045 2214 20000 2216
rect 18045 2211 18111 2214
rect 5394 2208 5710 2209
rect 5394 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5710 2208
rect 5394 2143 5710 2144
rect 9842 2208 10158 2209
rect 9842 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10158 2208
rect 9842 2143 10158 2144
rect 14290 2208 14606 2209
rect 14290 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14606 2208
rect 19200 2184 20000 2214
rect 14290 2143 14606 2144
rect 0 2002 800 2032
rect 2773 2002 2839 2005
rect 0 2000 2839 2002
rect 0 1944 2778 2000
rect 2834 1944 2839 2000
rect 0 1942 2839 1944
rect 0 1912 800 1942
rect 2773 1939 2839 1942
rect 18505 1866 18571 1869
rect 19200 1866 20000 1896
rect 18505 1864 20000 1866
rect 18505 1808 18510 1864
rect 18566 1808 20000 1864
rect 18505 1806 20000 1808
rect 18505 1803 18571 1806
rect 19200 1776 20000 1806
rect 0 1594 800 1624
rect 1945 1594 2011 1597
rect 0 1592 2011 1594
rect 0 1536 1950 1592
rect 2006 1536 2011 1592
rect 0 1534 2011 1536
rect 0 1504 800 1534
rect 1945 1531 2011 1534
rect 16849 1458 16915 1461
rect 19200 1458 20000 1488
rect 16849 1456 20000 1458
rect 16849 1400 16854 1456
rect 16910 1400 20000 1456
rect 16849 1398 20000 1400
rect 16849 1395 16915 1398
rect 19200 1368 20000 1398
rect 0 1186 800 1216
rect 3509 1186 3575 1189
rect 0 1184 3575 1186
rect 0 1128 3514 1184
rect 3570 1128 3575 1184
rect 0 1126 3575 1128
rect 0 1096 800 1126
rect 3509 1123 3575 1126
rect 17677 1050 17743 1053
rect 19200 1050 20000 1080
rect 17677 1048 20000 1050
rect 17677 992 17682 1048
rect 17738 992 20000 1048
rect 17677 990 20000 992
rect 17677 987 17743 990
rect 19200 960 20000 990
rect 3785 914 3851 917
rect 1350 912 3851 914
rect 1350 856 3790 912
rect 3846 856 3851 912
rect 1350 854 3851 856
rect 0 778 800 808
rect 1350 778 1410 854
rect 3785 851 3851 854
rect 0 718 1410 778
rect 0 688 800 718
rect 16389 642 16455 645
rect 19200 642 20000 672
rect 16389 640 20000 642
rect 16389 584 16394 640
rect 16450 584 20000 640
rect 16389 582 20000 584
rect 16389 579 16455 582
rect 19200 552 20000 582
rect 0 370 800 400
rect 2865 370 2931 373
rect 0 368 2931 370
rect 0 312 2870 368
rect 2926 312 2931 368
rect 0 310 2931 312
rect 0 280 800 310
rect 2865 307 2931 310
<< via3 >>
rect 3176 14716 3240 14720
rect 3176 14660 3180 14716
rect 3180 14660 3236 14716
rect 3236 14660 3240 14716
rect 3176 14656 3240 14660
rect 3256 14716 3320 14720
rect 3256 14660 3260 14716
rect 3260 14660 3316 14716
rect 3316 14660 3320 14716
rect 3256 14656 3320 14660
rect 3336 14716 3400 14720
rect 3336 14660 3340 14716
rect 3340 14660 3396 14716
rect 3396 14660 3400 14716
rect 3336 14656 3400 14660
rect 3416 14716 3480 14720
rect 3416 14660 3420 14716
rect 3420 14660 3476 14716
rect 3476 14660 3480 14716
rect 3416 14656 3480 14660
rect 7624 14716 7688 14720
rect 7624 14660 7628 14716
rect 7628 14660 7684 14716
rect 7684 14660 7688 14716
rect 7624 14656 7688 14660
rect 7704 14716 7768 14720
rect 7704 14660 7708 14716
rect 7708 14660 7764 14716
rect 7764 14660 7768 14716
rect 7704 14656 7768 14660
rect 7784 14716 7848 14720
rect 7784 14660 7788 14716
rect 7788 14660 7844 14716
rect 7844 14660 7848 14716
rect 7784 14656 7848 14660
rect 7864 14716 7928 14720
rect 7864 14660 7868 14716
rect 7868 14660 7924 14716
rect 7924 14660 7928 14716
rect 7864 14656 7928 14660
rect 12072 14716 12136 14720
rect 12072 14660 12076 14716
rect 12076 14660 12132 14716
rect 12132 14660 12136 14716
rect 12072 14656 12136 14660
rect 12152 14716 12216 14720
rect 12152 14660 12156 14716
rect 12156 14660 12212 14716
rect 12212 14660 12216 14716
rect 12152 14656 12216 14660
rect 12232 14716 12296 14720
rect 12232 14660 12236 14716
rect 12236 14660 12292 14716
rect 12292 14660 12296 14716
rect 12232 14656 12296 14660
rect 12312 14716 12376 14720
rect 12312 14660 12316 14716
rect 12316 14660 12372 14716
rect 12372 14660 12376 14716
rect 12312 14656 12376 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 16760 14716 16824 14720
rect 16760 14660 16764 14716
rect 16764 14660 16820 14716
rect 16820 14660 16824 14716
rect 16760 14656 16824 14660
rect 5400 14172 5464 14176
rect 5400 14116 5404 14172
rect 5404 14116 5460 14172
rect 5460 14116 5464 14172
rect 5400 14112 5464 14116
rect 5480 14172 5544 14176
rect 5480 14116 5484 14172
rect 5484 14116 5540 14172
rect 5540 14116 5544 14172
rect 5480 14112 5544 14116
rect 5560 14172 5624 14176
rect 5560 14116 5564 14172
rect 5564 14116 5620 14172
rect 5620 14116 5624 14172
rect 5560 14112 5624 14116
rect 5640 14172 5704 14176
rect 5640 14116 5644 14172
rect 5644 14116 5700 14172
rect 5700 14116 5704 14172
rect 5640 14112 5704 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 14536 14172 14600 14176
rect 14536 14116 14540 14172
rect 14540 14116 14596 14172
rect 14596 14116 14600 14172
rect 14536 14112 14600 14116
rect 9444 13908 9508 13972
rect 8892 13772 8956 13836
rect 14964 13636 15028 13700
rect 3176 13628 3240 13632
rect 3176 13572 3180 13628
rect 3180 13572 3236 13628
rect 3236 13572 3240 13628
rect 3176 13568 3240 13572
rect 3256 13628 3320 13632
rect 3256 13572 3260 13628
rect 3260 13572 3316 13628
rect 3316 13572 3320 13628
rect 3256 13568 3320 13572
rect 3336 13628 3400 13632
rect 3336 13572 3340 13628
rect 3340 13572 3396 13628
rect 3396 13572 3400 13628
rect 3336 13568 3400 13572
rect 3416 13628 3480 13632
rect 3416 13572 3420 13628
rect 3420 13572 3476 13628
rect 3476 13572 3480 13628
rect 3416 13568 3480 13572
rect 7624 13628 7688 13632
rect 7624 13572 7628 13628
rect 7628 13572 7684 13628
rect 7684 13572 7688 13628
rect 7624 13568 7688 13572
rect 7704 13628 7768 13632
rect 7704 13572 7708 13628
rect 7708 13572 7764 13628
rect 7764 13572 7768 13628
rect 7704 13568 7768 13572
rect 7784 13628 7848 13632
rect 7784 13572 7788 13628
rect 7788 13572 7844 13628
rect 7844 13572 7848 13628
rect 7784 13568 7848 13572
rect 7864 13628 7928 13632
rect 7864 13572 7868 13628
rect 7868 13572 7924 13628
rect 7924 13572 7928 13628
rect 7864 13568 7928 13572
rect 12072 13628 12136 13632
rect 12072 13572 12076 13628
rect 12076 13572 12132 13628
rect 12132 13572 12136 13628
rect 12072 13568 12136 13572
rect 12152 13628 12216 13632
rect 12152 13572 12156 13628
rect 12156 13572 12212 13628
rect 12212 13572 12216 13628
rect 12152 13568 12216 13572
rect 12232 13628 12296 13632
rect 12232 13572 12236 13628
rect 12236 13572 12292 13628
rect 12292 13572 12296 13628
rect 12232 13568 12296 13572
rect 12312 13628 12376 13632
rect 12312 13572 12316 13628
rect 12316 13572 12372 13628
rect 12372 13572 12376 13628
rect 12312 13568 12376 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 16760 13628 16824 13632
rect 16760 13572 16764 13628
rect 16764 13572 16820 13628
rect 16820 13572 16824 13628
rect 16760 13568 16824 13572
rect 5400 13084 5464 13088
rect 5400 13028 5404 13084
rect 5404 13028 5460 13084
rect 5460 13028 5464 13084
rect 5400 13024 5464 13028
rect 5480 13084 5544 13088
rect 5480 13028 5484 13084
rect 5484 13028 5540 13084
rect 5540 13028 5544 13084
rect 5480 13024 5544 13028
rect 5560 13084 5624 13088
rect 5560 13028 5564 13084
rect 5564 13028 5620 13084
rect 5620 13028 5624 13084
rect 5560 13024 5624 13028
rect 5640 13084 5704 13088
rect 5640 13028 5644 13084
rect 5644 13028 5700 13084
rect 5700 13028 5704 13084
rect 5640 13024 5704 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 14536 13084 14600 13088
rect 14536 13028 14540 13084
rect 14540 13028 14596 13084
rect 14596 13028 14600 13084
rect 14536 13024 14600 13028
rect 1348 12956 1412 13020
rect 3924 12880 3988 12884
rect 3924 12824 3938 12880
rect 3938 12824 3988 12880
rect 3924 12820 3988 12824
rect 3176 12540 3240 12544
rect 3176 12484 3180 12540
rect 3180 12484 3236 12540
rect 3236 12484 3240 12540
rect 3176 12480 3240 12484
rect 3256 12540 3320 12544
rect 3256 12484 3260 12540
rect 3260 12484 3316 12540
rect 3316 12484 3320 12540
rect 3256 12480 3320 12484
rect 3336 12540 3400 12544
rect 3336 12484 3340 12540
rect 3340 12484 3396 12540
rect 3396 12484 3400 12540
rect 3336 12480 3400 12484
rect 3416 12540 3480 12544
rect 3416 12484 3420 12540
rect 3420 12484 3476 12540
rect 3476 12484 3480 12540
rect 3416 12480 3480 12484
rect 7624 12540 7688 12544
rect 7624 12484 7628 12540
rect 7628 12484 7684 12540
rect 7684 12484 7688 12540
rect 7624 12480 7688 12484
rect 7704 12540 7768 12544
rect 7704 12484 7708 12540
rect 7708 12484 7764 12540
rect 7764 12484 7768 12540
rect 7704 12480 7768 12484
rect 7784 12540 7848 12544
rect 7784 12484 7788 12540
rect 7788 12484 7844 12540
rect 7844 12484 7848 12540
rect 7784 12480 7848 12484
rect 7864 12540 7928 12544
rect 7864 12484 7868 12540
rect 7868 12484 7924 12540
rect 7924 12484 7928 12540
rect 7864 12480 7928 12484
rect 12072 12540 12136 12544
rect 12072 12484 12076 12540
rect 12076 12484 12132 12540
rect 12132 12484 12136 12540
rect 12072 12480 12136 12484
rect 12152 12540 12216 12544
rect 12152 12484 12156 12540
rect 12156 12484 12212 12540
rect 12212 12484 12216 12540
rect 12152 12480 12216 12484
rect 12232 12540 12296 12544
rect 12232 12484 12236 12540
rect 12236 12484 12292 12540
rect 12292 12484 12296 12540
rect 12232 12480 12296 12484
rect 12312 12540 12376 12544
rect 12312 12484 12316 12540
rect 12316 12484 12372 12540
rect 12372 12484 12376 12540
rect 12312 12480 12376 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 16760 12540 16824 12544
rect 16760 12484 16764 12540
rect 16764 12484 16820 12540
rect 16820 12484 16824 12540
rect 16760 12480 16824 12484
rect 4108 12140 4172 12204
rect 5400 11996 5464 12000
rect 5400 11940 5404 11996
rect 5404 11940 5460 11996
rect 5460 11940 5464 11996
rect 5400 11936 5464 11940
rect 5480 11996 5544 12000
rect 5480 11940 5484 11996
rect 5484 11940 5540 11996
rect 5540 11940 5544 11996
rect 5480 11936 5544 11940
rect 5560 11996 5624 12000
rect 5560 11940 5564 11996
rect 5564 11940 5620 11996
rect 5620 11940 5624 11996
rect 5560 11936 5624 11940
rect 5640 11996 5704 12000
rect 5640 11940 5644 11996
rect 5644 11940 5700 11996
rect 5700 11940 5704 11996
rect 5640 11936 5704 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 14536 11996 14600 12000
rect 14536 11940 14540 11996
rect 14540 11940 14596 11996
rect 14596 11940 14600 11996
rect 14536 11936 14600 11940
rect 3176 11452 3240 11456
rect 3176 11396 3180 11452
rect 3180 11396 3236 11452
rect 3236 11396 3240 11452
rect 3176 11392 3240 11396
rect 3256 11452 3320 11456
rect 3256 11396 3260 11452
rect 3260 11396 3316 11452
rect 3316 11396 3320 11452
rect 3256 11392 3320 11396
rect 3336 11452 3400 11456
rect 3336 11396 3340 11452
rect 3340 11396 3396 11452
rect 3396 11396 3400 11452
rect 3336 11392 3400 11396
rect 3416 11452 3480 11456
rect 3416 11396 3420 11452
rect 3420 11396 3476 11452
rect 3476 11396 3480 11452
rect 3416 11392 3480 11396
rect 7624 11452 7688 11456
rect 7624 11396 7628 11452
rect 7628 11396 7684 11452
rect 7684 11396 7688 11452
rect 7624 11392 7688 11396
rect 7704 11452 7768 11456
rect 7704 11396 7708 11452
rect 7708 11396 7764 11452
rect 7764 11396 7768 11452
rect 7704 11392 7768 11396
rect 7784 11452 7848 11456
rect 7784 11396 7788 11452
rect 7788 11396 7844 11452
rect 7844 11396 7848 11452
rect 7784 11392 7848 11396
rect 7864 11452 7928 11456
rect 7864 11396 7868 11452
rect 7868 11396 7924 11452
rect 7924 11396 7928 11452
rect 7864 11392 7928 11396
rect 12072 11452 12136 11456
rect 12072 11396 12076 11452
rect 12076 11396 12132 11452
rect 12132 11396 12136 11452
rect 12072 11392 12136 11396
rect 12152 11452 12216 11456
rect 12152 11396 12156 11452
rect 12156 11396 12212 11452
rect 12212 11396 12216 11452
rect 12152 11392 12216 11396
rect 12232 11452 12296 11456
rect 12232 11396 12236 11452
rect 12236 11396 12292 11452
rect 12292 11396 12296 11452
rect 12232 11392 12296 11396
rect 12312 11452 12376 11456
rect 12312 11396 12316 11452
rect 12316 11396 12372 11452
rect 12372 11396 12376 11452
rect 12312 11392 12376 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 16760 11452 16824 11456
rect 16760 11396 16764 11452
rect 16764 11396 16820 11452
rect 16820 11396 16824 11452
rect 16760 11392 16824 11396
rect 5400 10908 5464 10912
rect 5400 10852 5404 10908
rect 5404 10852 5460 10908
rect 5460 10852 5464 10908
rect 5400 10848 5464 10852
rect 5480 10908 5544 10912
rect 5480 10852 5484 10908
rect 5484 10852 5540 10908
rect 5540 10852 5544 10908
rect 5480 10848 5544 10852
rect 5560 10908 5624 10912
rect 5560 10852 5564 10908
rect 5564 10852 5620 10908
rect 5620 10852 5624 10908
rect 5560 10848 5624 10852
rect 5640 10908 5704 10912
rect 5640 10852 5644 10908
rect 5644 10852 5700 10908
rect 5700 10852 5704 10908
rect 5640 10848 5704 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 14536 10908 14600 10912
rect 14536 10852 14540 10908
rect 14540 10852 14596 10908
rect 14596 10852 14600 10908
rect 14536 10848 14600 10852
rect 3176 10364 3240 10368
rect 3176 10308 3180 10364
rect 3180 10308 3236 10364
rect 3236 10308 3240 10364
rect 3176 10304 3240 10308
rect 3256 10364 3320 10368
rect 3256 10308 3260 10364
rect 3260 10308 3316 10364
rect 3316 10308 3320 10364
rect 3256 10304 3320 10308
rect 3336 10364 3400 10368
rect 3336 10308 3340 10364
rect 3340 10308 3396 10364
rect 3396 10308 3400 10364
rect 3336 10304 3400 10308
rect 3416 10364 3480 10368
rect 3416 10308 3420 10364
rect 3420 10308 3476 10364
rect 3476 10308 3480 10364
rect 3416 10304 3480 10308
rect 7624 10364 7688 10368
rect 7624 10308 7628 10364
rect 7628 10308 7684 10364
rect 7684 10308 7688 10364
rect 7624 10304 7688 10308
rect 7704 10364 7768 10368
rect 7704 10308 7708 10364
rect 7708 10308 7764 10364
rect 7764 10308 7768 10364
rect 7704 10304 7768 10308
rect 7784 10364 7848 10368
rect 7784 10308 7788 10364
rect 7788 10308 7844 10364
rect 7844 10308 7848 10364
rect 7784 10304 7848 10308
rect 7864 10364 7928 10368
rect 7864 10308 7868 10364
rect 7868 10308 7924 10364
rect 7924 10308 7928 10364
rect 7864 10304 7928 10308
rect 12072 10364 12136 10368
rect 12072 10308 12076 10364
rect 12076 10308 12132 10364
rect 12132 10308 12136 10364
rect 12072 10304 12136 10308
rect 12152 10364 12216 10368
rect 12152 10308 12156 10364
rect 12156 10308 12212 10364
rect 12212 10308 12216 10364
rect 12152 10304 12216 10308
rect 12232 10364 12296 10368
rect 12232 10308 12236 10364
rect 12236 10308 12292 10364
rect 12292 10308 12296 10364
rect 12232 10304 12296 10308
rect 12312 10364 12376 10368
rect 12312 10308 12316 10364
rect 12316 10308 12372 10364
rect 12372 10308 12376 10364
rect 12312 10304 12376 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 16760 10364 16824 10368
rect 16760 10308 16764 10364
rect 16764 10308 16820 10364
rect 16820 10308 16824 10364
rect 16760 10304 16824 10308
rect 5400 9820 5464 9824
rect 5400 9764 5404 9820
rect 5404 9764 5460 9820
rect 5460 9764 5464 9820
rect 5400 9760 5464 9764
rect 5480 9820 5544 9824
rect 5480 9764 5484 9820
rect 5484 9764 5540 9820
rect 5540 9764 5544 9820
rect 5480 9760 5544 9764
rect 5560 9820 5624 9824
rect 5560 9764 5564 9820
rect 5564 9764 5620 9820
rect 5620 9764 5624 9820
rect 5560 9760 5624 9764
rect 5640 9820 5704 9824
rect 5640 9764 5644 9820
rect 5644 9764 5700 9820
rect 5700 9764 5704 9820
rect 5640 9760 5704 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 14536 9820 14600 9824
rect 14536 9764 14540 9820
rect 14540 9764 14596 9820
rect 14596 9764 14600 9820
rect 14536 9760 14600 9764
rect 3924 9556 3988 9620
rect 3176 9276 3240 9280
rect 3176 9220 3180 9276
rect 3180 9220 3236 9276
rect 3236 9220 3240 9276
rect 3176 9216 3240 9220
rect 3256 9276 3320 9280
rect 3256 9220 3260 9276
rect 3260 9220 3316 9276
rect 3316 9220 3320 9276
rect 3256 9216 3320 9220
rect 3336 9276 3400 9280
rect 3336 9220 3340 9276
rect 3340 9220 3396 9276
rect 3396 9220 3400 9276
rect 3336 9216 3400 9220
rect 3416 9276 3480 9280
rect 3416 9220 3420 9276
rect 3420 9220 3476 9276
rect 3476 9220 3480 9276
rect 3416 9216 3480 9220
rect 7624 9276 7688 9280
rect 7624 9220 7628 9276
rect 7628 9220 7684 9276
rect 7684 9220 7688 9276
rect 7624 9216 7688 9220
rect 7704 9276 7768 9280
rect 7704 9220 7708 9276
rect 7708 9220 7764 9276
rect 7764 9220 7768 9276
rect 7704 9216 7768 9220
rect 7784 9276 7848 9280
rect 7784 9220 7788 9276
rect 7788 9220 7844 9276
rect 7844 9220 7848 9276
rect 7784 9216 7848 9220
rect 7864 9276 7928 9280
rect 7864 9220 7868 9276
rect 7868 9220 7924 9276
rect 7924 9220 7928 9276
rect 7864 9216 7928 9220
rect 12072 9276 12136 9280
rect 12072 9220 12076 9276
rect 12076 9220 12132 9276
rect 12132 9220 12136 9276
rect 12072 9216 12136 9220
rect 12152 9276 12216 9280
rect 12152 9220 12156 9276
rect 12156 9220 12212 9276
rect 12212 9220 12216 9276
rect 12152 9216 12216 9220
rect 12232 9276 12296 9280
rect 12232 9220 12236 9276
rect 12236 9220 12292 9276
rect 12292 9220 12296 9276
rect 12232 9216 12296 9220
rect 12312 9276 12376 9280
rect 12312 9220 12316 9276
rect 12316 9220 12372 9276
rect 12372 9220 12376 9276
rect 12312 9216 12376 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 16760 9276 16824 9280
rect 16760 9220 16764 9276
rect 16764 9220 16820 9276
rect 16820 9220 16824 9276
rect 16760 9216 16824 9220
rect 4108 9012 4172 9076
rect 2636 8740 2700 8804
rect 5400 8732 5464 8736
rect 5400 8676 5404 8732
rect 5404 8676 5460 8732
rect 5460 8676 5464 8732
rect 5400 8672 5464 8676
rect 5480 8732 5544 8736
rect 5480 8676 5484 8732
rect 5484 8676 5540 8732
rect 5540 8676 5544 8732
rect 5480 8672 5544 8676
rect 5560 8732 5624 8736
rect 5560 8676 5564 8732
rect 5564 8676 5620 8732
rect 5620 8676 5624 8732
rect 5560 8672 5624 8676
rect 5640 8732 5704 8736
rect 5640 8676 5644 8732
rect 5644 8676 5700 8732
rect 5700 8676 5704 8732
rect 5640 8672 5704 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 14536 8732 14600 8736
rect 14536 8676 14540 8732
rect 14540 8676 14596 8732
rect 14596 8676 14600 8732
rect 14536 8672 14600 8676
rect 1348 8196 1412 8260
rect 3176 8188 3240 8192
rect 3176 8132 3180 8188
rect 3180 8132 3236 8188
rect 3236 8132 3240 8188
rect 3176 8128 3240 8132
rect 3256 8188 3320 8192
rect 3256 8132 3260 8188
rect 3260 8132 3316 8188
rect 3316 8132 3320 8188
rect 3256 8128 3320 8132
rect 3336 8188 3400 8192
rect 3336 8132 3340 8188
rect 3340 8132 3396 8188
rect 3396 8132 3400 8188
rect 3336 8128 3400 8132
rect 3416 8188 3480 8192
rect 3416 8132 3420 8188
rect 3420 8132 3476 8188
rect 3476 8132 3480 8188
rect 3416 8128 3480 8132
rect 7624 8188 7688 8192
rect 7624 8132 7628 8188
rect 7628 8132 7684 8188
rect 7684 8132 7688 8188
rect 7624 8128 7688 8132
rect 7704 8188 7768 8192
rect 7704 8132 7708 8188
rect 7708 8132 7764 8188
rect 7764 8132 7768 8188
rect 7704 8128 7768 8132
rect 7784 8188 7848 8192
rect 7784 8132 7788 8188
rect 7788 8132 7844 8188
rect 7844 8132 7848 8188
rect 7784 8128 7848 8132
rect 7864 8188 7928 8192
rect 7864 8132 7868 8188
rect 7868 8132 7924 8188
rect 7924 8132 7928 8188
rect 7864 8128 7928 8132
rect 12072 8188 12136 8192
rect 12072 8132 12076 8188
rect 12076 8132 12132 8188
rect 12132 8132 12136 8188
rect 12072 8128 12136 8132
rect 12152 8188 12216 8192
rect 12152 8132 12156 8188
rect 12156 8132 12212 8188
rect 12212 8132 12216 8188
rect 12152 8128 12216 8132
rect 12232 8188 12296 8192
rect 12232 8132 12236 8188
rect 12236 8132 12292 8188
rect 12292 8132 12296 8188
rect 12232 8128 12296 8132
rect 12312 8188 12376 8192
rect 12312 8132 12316 8188
rect 12316 8132 12372 8188
rect 12372 8132 12376 8188
rect 12312 8128 12376 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 16760 8188 16824 8192
rect 16760 8132 16764 8188
rect 16764 8132 16820 8188
rect 16820 8132 16824 8188
rect 16760 8128 16824 8132
rect 5400 7644 5464 7648
rect 5400 7588 5404 7644
rect 5404 7588 5460 7644
rect 5460 7588 5464 7644
rect 5400 7584 5464 7588
rect 5480 7644 5544 7648
rect 5480 7588 5484 7644
rect 5484 7588 5540 7644
rect 5540 7588 5544 7644
rect 5480 7584 5544 7588
rect 5560 7644 5624 7648
rect 5560 7588 5564 7644
rect 5564 7588 5620 7644
rect 5620 7588 5624 7644
rect 5560 7584 5624 7588
rect 5640 7644 5704 7648
rect 5640 7588 5644 7644
rect 5644 7588 5700 7644
rect 5700 7588 5704 7644
rect 5640 7584 5704 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 14536 7644 14600 7648
rect 14536 7588 14540 7644
rect 14540 7588 14596 7644
rect 14596 7588 14600 7644
rect 14536 7584 14600 7588
rect 3176 7100 3240 7104
rect 3176 7044 3180 7100
rect 3180 7044 3236 7100
rect 3236 7044 3240 7100
rect 3176 7040 3240 7044
rect 3256 7100 3320 7104
rect 3256 7044 3260 7100
rect 3260 7044 3316 7100
rect 3316 7044 3320 7100
rect 3256 7040 3320 7044
rect 3336 7100 3400 7104
rect 3336 7044 3340 7100
rect 3340 7044 3396 7100
rect 3396 7044 3400 7100
rect 3336 7040 3400 7044
rect 3416 7100 3480 7104
rect 3416 7044 3420 7100
rect 3420 7044 3476 7100
rect 3476 7044 3480 7100
rect 3416 7040 3480 7044
rect 7624 7100 7688 7104
rect 7624 7044 7628 7100
rect 7628 7044 7684 7100
rect 7684 7044 7688 7100
rect 7624 7040 7688 7044
rect 7704 7100 7768 7104
rect 7704 7044 7708 7100
rect 7708 7044 7764 7100
rect 7764 7044 7768 7100
rect 7704 7040 7768 7044
rect 7784 7100 7848 7104
rect 7784 7044 7788 7100
rect 7788 7044 7844 7100
rect 7844 7044 7848 7100
rect 7784 7040 7848 7044
rect 7864 7100 7928 7104
rect 7864 7044 7868 7100
rect 7868 7044 7924 7100
rect 7924 7044 7928 7100
rect 7864 7040 7928 7044
rect 12072 7100 12136 7104
rect 12072 7044 12076 7100
rect 12076 7044 12132 7100
rect 12132 7044 12136 7100
rect 12072 7040 12136 7044
rect 12152 7100 12216 7104
rect 12152 7044 12156 7100
rect 12156 7044 12212 7100
rect 12212 7044 12216 7100
rect 12152 7040 12216 7044
rect 12232 7100 12296 7104
rect 12232 7044 12236 7100
rect 12236 7044 12292 7100
rect 12292 7044 12296 7100
rect 12232 7040 12296 7044
rect 12312 7100 12376 7104
rect 12312 7044 12316 7100
rect 12316 7044 12372 7100
rect 12372 7044 12376 7100
rect 12312 7040 12376 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 16760 7100 16824 7104
rect 16760 7044 16764 7100
rect 16764 7044 16820 7100
rect 16820 7044 16824 7100
rect 16760 7040 16824 7044
rect 2636 6700 2700 6764
rect 5400 6556 5464 6560
rect 5400 6500 5404 6556
rect 5404 6500 5460 6556
rect 5460 6500 5464 6556
rect 5400 6496 5464 6500
rect 5480 6556 5544 6560
rect 5480 6500 5484 6556
rect 5484 6500 5540 6556
rect 5540 6500 5544 6556
rect 5480 6496 5544 6500
rect 5560 6556 5624 6560
rect 5560 6500 5564 6556
rect 5564 6500 5620 6556
rect 5620 6500 5624 6556
rect 5560 6496 5624 6500
rect 5640 6556 5704 6560
rect 5640 6500 5644 6556
rect 5644 6500 5700 6556
rect 5700 6500 5704 6556
rect 5640 6496 5704 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 14536 6556 14600 6560
rect 14536 6500 14540 6556
rect 14540 6500 14596 6556
rect 14596 6500 14600 6556
rect 14536 6496 14600 6500
rect 3176 6012 3240 6016
rect 3176 5956 3180 6012
rect 3180 5956 3236 6012
rect 3236 5956 3240 6012
rect 3176 5952 3240 5956
rect 3256 6012 3320 6016
rect 3256 5956 3260 6012
rect 3260 5956 3316 6012
rect 3316 5956 3320 6012
rect 3256 5952 3320 5956
rect 3336 6012 3400 6016
rect 3336 5956 3340 6012
rect 3340 5956 3396 6012
rect 3396 5956 3400 6012
rect 3336 5952 3400 5956
rect 3416 6012 3480 6016
rect 3416 5956 3420 6012
rect 3420 5956 3476 6012
rect 3476 5956 3480 6012
rect 3416 5952 3480 5956
rect 7624 6012 7688 6016
rect 7624 5956 7628 6012
rect 7628 5956 7684 6012
rect 7684 5956 7688 6012
rect 7624 5952 7688 5956
rect 7704 6012 7768 6016
rect 7704 5956 7708 6012
rect 7708 5956 7764 6012
rect 7764 5956 7768 6012
rect 7704 5952 7768 5956
rect 7784 6012 7848 6016
rect 7784 5956 7788 6012
rect 7788 5956 7844 6012
rect 7844 5956 7848 6012
rect 7784 5952 7848 5956
rect 7864 6012 7928 6016
rect 7864 5956 7868 6012
rect 7868 5956 7924 6012
rect 7924 5956 7928 6012
rect 7864 5952 7928 5956
rect 12072 6012 12136 6016
rect 12072 5956 12076 6012
rect 12076 5956 12132 6012
rect 12132 5956 12136 6012
rect 12072 5952 12136 5956
rect 12152 6012 12216 6016
rect 12152 5956 12156 6012
rect 12156 5956 12212 6012
rect 12212 5956 12216 6012
rect 12152 5952 12216 5956
rect 12232 6012 12296 6016
rect 12232 5956 12236 6012
rect 12236 5956 12292 6012
rect 12292 5956 12296 6012
rect 12232 5952 12296 5956
rect 12312 6012 12376 6016
rect 12312 5956 12316 6012
rect 12316 5956 12372 6012
rect 12372 5956 12376 6012
rect 12312 5952 12376 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 16760 6012 16824 6016
rect 16760 5956 16764 6012
rect 16764 5956 16820 6012
rect 16820 5956 16824 6012
rect 16760 5952 16824 5956
rect 5400 5468 5464 5472
rect 5400 5412 5404 5468
rect 5404 5412 5460 5468
rect 5460 5412 5464 5468
rect 5400 5408 5464 5412
rect 5480 5468 5544 5472
rect 5480 5412 5484 5468
rect 5484 5412 5540 5468
rect 5540 5412 5544 5468
rect 5480 5408 5544 5412
rect 5560 5468 5624 5472
rect 5560 5412 5564 5468
rect 5564 5412 5620 5468
rect 5620 5412 5624 5468
rect 5560 5408 5624 5412
rect 5640 5468 5704 5472
rect 5640 5412 5644 5468
rect 5644 5412 5700 5468
rect 5700 5412 5704 5468
rect 5640 5408 5704 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 14536 5468 14600 5472
rect 14536 5412 14540 5468
rect 14540 5412 14596 5468
rect 14596 5412 14600 5468
rect 14536 5408 14600 5412
rect 3176 4924 3240 4928
rect 3176 4868 3180 4924
rect 3180 4868 3236 4924
rect 3236 4868 3240 4924
rect 3176 4864 3240 4868
rect 3256 4924 3320 4928
rect 3256 4868 3260 4924
rect 3260 4868 3316 4924
rect 3316 4868 3320 4924
rect 3256 4864 3320 4868
rect 3336 4924 3400 4928
rect 3336 4868 3340 4924
rect 3340 4868 3396 4924
rect 3396 4868 3400 4924
rect 3336 4864 3400 4868
rect 3416 4924 3480 4928
rect 3416 4868 3420 4924
rect 3420 4868 3476 4924
rect 3476 4868 3480 4924
rect 3416 4864 3480 4868
rect 7624 4924 7688 4928
rect 7624 4868 7628 4924
rect 7628 4868 7684 4924
rect 7684 4868 7688 4924
rect 7624 4864 7688 4868
rect 7704 4924 7768 4928
rect 7704 4868 7708 4924
rect 7708 4868 7764 4924
rect 7764 4868 7768 4924
rect 7704 4864 7768 4868
rect 7784 4924 7848 4928
rect 7784 4868 7788 4924
rect 7788 4868 7844 4924
rect 7844 4868 7848 4924
rect 7784 4864 7848 4868
rect 7864 4924 7928 4928
rect 7864 4868 7868 4924
rect 7868 4868 7924 4924
rect 7924 4868 7928 4924
rect 7864 4864 7928 4868
rect 12072 4924 12136 4928
rect 12072 4868 12076 4924
rect 12076 4868 12132 4924
rect 12132 4868 12136 4924
rect 12072 4864 12136 4868
rect 12152 4924 12216 4928
rect 12152 4868 12156 4924
rect 12156 4868 12212 4924
rect 12212 4868 12216 4924
rect 12152 4864 12216 4868
rect 12232 4924 12296 4928
rect 12232 4868 12236 4924
rect 12236 4868 12292 4924
rect 12292 4868 12296 4924
rect 12232 4864 12296 4868
rect 12312 4924 12376 4928
rect 12312 4868 12316 4924
rect 12316 4868 12372 4924
rect 12372 4868 12376 4924
rect 12312 4864 12376 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 16760 4924 16824 4928
rect 16760 4868 16764 4924
rect 16764 4868 16820 4924
rect 16820 4868 16824 4924
rect 16760 4864 16824 4868
rect 4108 4796 4172 4860
rect 5400 4380 5464 4384
rect 5400 4324 5404 4380
rect 5404 4324 5460 4380
rect 5460 4324 5464 4380
rect 5400 4320 5464 4324
rect 5480 4380 5544 4384
rect 5480 4324 5484 4380
rect 5484 4324 5540 4380
rect 5540 4324 5544 4380
rect 5480 4320 5544 4324
rect 5560 4380 5624 4384
rect 5560 4324 5564 4380
rect 5564 4324 5620 4380
rect 5620 4324 5624 4380
rect 5560 4320 5624 4324
rect 5640 4380 5704 4384
rect 5640 4324 5644 4380
rect 5644 4324 5700 4380
rect 5700 4324 5704 4380
rect 5640 4320 5704 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 14536 4380 14600 4384
rect 14536 4324 14540 4380
rect 14540 4324 14596 4380
rect 14596 4324 14600 4380
rect 14536 4320 14600 4324
rect 8892 3980 8956 4044
rect 9444 3980 9508 4044
rect 3176 3836 3240 3840
rect 3176 3780 3180 3836
rect 3180 3780 3236 3836
rect 3236 3780 3240 3836
rect 3176 3776 3240 3780
rect 3256 3836 3320 3840
rect 3256 3780 3260 3836
rect 3260 3780 3316 3836
rect 3316 3780 3320 3836
rect 3256 3776 3320 3780
rect 3336 3836 3400 3840
rect 3336 3780 3340 3836
rect 3340 3780 3396 3836
rect 3396 3780 3400 3836
rect 3336 3776 3400 3780
rect 3416 3836 3480 3840
rect 3416 3780 3420 3836
rect 3420 3780 3476 3836
rect 3476 3780 3480 3836
rect 3416 3776 3480 3780
rect 7624 3836 7688 3840
rect 7624 3780 7628 3836
rect 7628 3780 7684 3836
rect 7684 3780 7688 3836
rect 7624 3776 7688 3780
rect 7704 3836 7768 3840
rect 7704 3780 7708 3836
rect 7708 3780 7764 3836
rect 7764 3780 7768 3836
rect 7704 3776 7768 3780
rect 7784 3836 7848 3840
rect 7784 3780 7788 3836
rect 7788 3780 7844 3836
rect 7844 3780 7848 3836
rect 7784 3776 7848 3780
rect 7864 3836 7928 3840
rect 7864 3780 7868 3836
rect 7868 3780 7924 3836
rect 7924 3780 7928 3836
rect 7864 3776 7928 3780
rect 12072 3836 12136 3840
rect 12072 3780 12076 3836
rect 12076 3780 12132 3836
rect 12132 3780 12136 3836
rect 12072 3776 12136 3780
rect 12152 3836 12216 3840
rect 12152 3780 12156 3836
rect 12156 3780 12212 3836
rect 12212 3780 12216 3836
rect 12152 3776 12216 3780
rect 12232 3836 12296 3840
rect 12232 3780 12236 3836
rect 12236 3780 12292 3836
rect 12292 3780 12296 3836
rect 12232 3776 12296 3780
rect 12312 3836 12376 3840
rect 12312 3780 12316 3836
rect 12316 3780 12372 3836
rect 12372 3780 12376 3836
rect 12312 3776 12376 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 16760 3836 16824 3840
rect 16760 3780 16764 3836
rect 16764 3780 16820 3836
rect 16820 3780 16824 3836
rect 16760 3776 16824 3780
rect 14964 3708 15028 3772
rect 5400 3292 5464 3296
rect 5400 3236 5404 3292
rect 5404 3236 5460 3292
rect 5460 3236 5464 3292
rect 5400 3232 5464 3236
rect 5480 3292 5544 3296
rect 5480 3236 5484 3292
rect 5484 3236 5540 3292
rect 5540 3236 5544 3292
rect 5480 3232 5544 3236
rect 5560 3292 5624 3296
rect 5560 3236 5564 3292
rect 5564 3236 5620 3292
rect 5620 3236 5624 3292
rect 5560 3232 5624 3236
rect 5640 3292 5704 3296
rect 5640 3236 5644 3292
rect 5644 3236 5700 3292
rect 5700 3236 5704 3292
rect 5640 3232 5704 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 14536 3292 14600 3296
rect 14536 3236 14540 3292
rect 14540 3236 14596 3292
rect 14596 3236 14600 3292
rect 14536 3232 14600 3236
rect 3176 2748 3240 2752
rect 3176 2692 3180 2748
rect 3180 2692 3236 2748
rect 3236 2692 3240 2748
rect 3176 2688 3240 2692
rect 3256 2748 3320 2752
rect 3256 2692 3260 2748
rect 3260 2692 3316 2748
rect 3316 2692 3320 2748
rect 3256 2688 3320 2692
rect 3336 2748 3400 2752
rect 3336 2692 3340 2748
rect 3340 2692 3396 2748
rect 3396 2692 3400 2748
rect 3336 2688 3400 2692
rect 3416 2748 3480 2752
rect 3416 2692 3420 2748
rect 3420 2692 3476 2748
rect 3476 2692 3480 2748
rect 3416 2688 3480 2692
rect 7624 2748 7688 2752
rect 7624 2692 7628 2748
rect 7628 2692 7684 2748
rect 7684 2692 7688 2748
rect 7624 2688 7688 2692
rect 7704 2748 7768 2752
rect 7704 2692 7708 2748
rect 7708 2692 7764 2748
rect 7764 2692 7768 2748
rect 7704 2688 7768 2692
rect 7784 2748 7848 2752
rect 7784 2692 7788 2748
rect 7788 2692 7844 2748
rect 7844 2692 7848 2748
rect 7784 2688 7848 2692
rect 7864 2748 7928 2752
rect 7864 2692 7868 2748
rect 7868 2692 7924 2748
rect 7924 2692 7928 2748
rect 7864 2688 7928 2692
rect 12072 2748 12136 2752
rect 12072 2692 12076 2748
rect 12076 2692 12132 2748
rect 12132 2692 12136 2748
rect 12072 2688 12136 2692
rect 12152 2748 12216 2752
rect 12152 2692 12156 2748
rect 12156 2692 12212 2748
rect 12212 2692 12216 2748
rect 12152 2688 12216 2692
rect 12232 2748 12296 2752
rect 12232 2692 12236 2748
rect 12236 2692 12292 2748
rect 12292 2692 12296 2748
rect 12232 2688 12296 2692
rect 12312 2748 12376 2752
rect 12312 2692 12316 2748
rect 12316 2692 12372 2748
rect 12372 2692 12376 2748
rect 12312 2688 12376 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 16760 2748 16824 2752
rect 16760 2692 16764 2748
rect 16764 2692 16820 2748
rect 16820 2692 16824 2748
rect 16760 2688 16824 2692
rect 5400 2204 5464 2208
rect 5400 2148 5404 2204
rect 5404 2148 5460 2204
rect 5460 2148 5464 2204
rect 5400 2144 5464 2148
rect 5480 2204 5544 2208
rect 5480 2148 5484 2204
rect 5484 2148 5540 2204
rect 5540 2148 5544 2204
rect 5480 2144 5544 2148
rect 5560 2204 5624 2208
rect 5560 2148 5564 2204
rect 5564 2148 5620 2204
rect 5620 2148 5624 2204
rect 5560 2144 5624 2148
rect 5640 2204 5704 2208
rect 5640 2148 5644 2204
rect 5644 2148 5700 2204
rect 5700 2148 5704 2204
rect 5640 2144 5704 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 14536 2204 14600 2208
rect 14536 2148 14540 2204
rect 14540 2148 14596 2204
rect 14596 2148 14600 2204
rect 14536 2144 14600 2148
<< metal4 >>
rect 3168 14720 3488 14736
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3168 13632 3488 14656
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 1347 13020 1413 13021
rect 1347 12956 1348 13020
rect 1412 12956 1413 13020
rect 1347 12955 1413 12956
rect 1350 8261 1410 12955
rect 3168 12544 3488 13568
rect 5392 14176 5712 14736
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 5392 13088 5712 14112
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 3923 12884 3989 12885
rect 3923 12820 3924 12884
rect 3988 12820 3989 12884
rect 3923 12819 3989 12820
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 3168 11456 3488 12480
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 3168 10368 3488 11392
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3168 9280 3488 10304
rect 3926 9621 3986 12819
rect 4107 12204 4173 12205
rect 4107 12140 4108 12204
rect 4172 12140 4173 12204
rect 4107 12139 4173 12140
rect 3923 9620 3989 9621
rect 3923 9556 3924 9620
rect 3988 9556 3989 9620
rect 3923 9555 3989 9556
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 2635 8804 2701 8805
rect 2635 8740 2636 8804
rect 2700 8740 2701 8804
rect 2635 8739 2701 8740
rect 1347 8260 1413 8261
rect 1347 8196 1348 8260
rect 1412 8196 1413 8260
rect 1347 8195 1413 8196
rect 2638 6765 2698 8739
rect 3168 8192 3488 9216
rect 4110 9077 4170 12139
rect 5392 12000 5712 13024
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5392 10912 5712 11936
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 9824 5712 10848
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 4107 9076 4173 9077
rect 4107 9012 4108 9076
rect 4172 9012 4173 9076
rect 4107 9011 4173 9012
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 3168 7104 3488 8128
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 2635 6764 2701 6765
rect 2635 6700 2636 6764
rect 2700 6700 2701 6764
rect 2635 6699 2701 6700
rect 3168 6016 3488 7040
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 3168 4928 3488 5952
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 3168 3840 3488 4864
rect 4110 4861 4170 9011
rect 5392 8736 5712 9760
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 7648 5712 8672
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5392 6560 5712 7584
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5392 5472 5712 6496
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 4107 4860 4173 4861
rect 4107 4796 4108 4860
rect 4172 4796 4173 4860
rect 4107 4795 4173 4796
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 3168 2752 3488 3776
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2128 3488 2688
rect 5392 4384 5712 5408
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 5392 3296 5712 4320
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 5392 2208 5712 3232
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2128 5712 2144
rect 7616 14720 7936 14736
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 7616 13632 7936 14656
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9443 13972 9509 13973
rect 9443 13908 9444 13972
rect 9508 13908 9509 13972
rect 9443 13907 9509 13908
rect 8891 13836 8957 13837
rect 8891 13772 8892 13836
rect 8956 13772 8957 13836
rect 8891 13771 8957 13772
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 7616 12544 7936 13568
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 7616 11456 7936 12480
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7616 10368 7936 11392
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7616 9280 7936 10304
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7616 8192 7936 9216
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7616 7104 7936 8128
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 6016 7936 7040
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 4928 7936 5952
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 3840 7936 4864
rect 8894 4045 8954 13771
rect 9446 4045 9506 13907
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 8891 4044 8957 4045
rect 8891 3980 8892 4044
rect 8956 3980 8957 4044
rect 8891 3979 8957 3980
rect 9443 4044 9509 4045
rect 9443 3980 9444 4044
rect 9508 3980 9509 4044
rect 9443 3979 9509 3980
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 7616 2752 7936 3776
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 7616 2128 7936 2688
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12064 14720 12384 14736
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 13632 12384 14656
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 12064 12544 12384 13568
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 12064 11456 12384 12480
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 10368 12384 11392
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 9280 12384 10304
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 8192 12384 9216
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 7104 12384 8128
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 6016 12384 7040
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 4928 12384 5952
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 3840 12384 4864
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 2752 12384 3776
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 12064 2128 12384 2688
rect 14288 14176 14608 14736
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 14288 13088 14608 14112
rect 16512 14720 16832 14736
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 14963 13700 15029 13701
rect 14963 13636 14964 13700
rect 15028 13636 15029 13700
rect 14963 13635 15029 13636
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 14288 12000 14608 13024
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 14288 10912 14608 11936
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 9824 14608 10848
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 14288 8736 14608 9760
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 14288 7648 14608 8672
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 6560 14608 7584
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 14288 5472 14608 6496
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 14288 4384 14608 5408
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 14288 3296 14608 4320
rect 14966 3773 15026 13635
rect 16512 13632 16832 14656
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 12544 16832 13568
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 16512 11456 16832 12480
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 10368 16832 11392
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 16512 9280 16832 10304
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 8192 16832 9216
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 16512 7104 16832 8128
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16512 6016 16832 7040
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16512 4928 16832 5952
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 16512 3840 16832 4864
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 14963 3772 15029 3773
rect 14963 3708 14964 3772
rect 15028 3708 15029 3772
rect 14963 3707 15029 3708
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 14288 2208 14608 3232
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 14288 2128 14608 2144
rect 16512 2752 16832 3776
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 16512 2128 16832 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1649977179
transform -1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1649977179
transform 1 0 2576 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1649977179
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1649977179
transform -1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1649977179
transform 1 0 1656 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1649977179
transform -1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1649977179
transform -1 0 2668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1649977179
transform -1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1649977179
transform 1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1649977179
transform -1 0 2668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1649977179
transform -1 0 1564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1649977179
transform -1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1649977179
transform 1 0 2024 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1649977179
transform -1 0 2852 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1649977179
transform -1 0 16468 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1649977179
transform -1 0 17664 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform -1 0 17204 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform 1 0 17664 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform 1 0 17664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform -1 0 17848 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 17480 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform -1 0 17756 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform -1 0 17756 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform -1 0 17756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform 1 0 17664 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1649977179
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform 1 0 17296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform 1 0 17664 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform -1 0 18216 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform -1 0 17848 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform -1 0 18400 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform -1 0 18216 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1649977179
transform -1 0 17848 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform 1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1649977179
transform 1 0 9016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1649977179
transform 1 0 7636 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1649977179
transform 1 0 11776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1649977179
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1649977179
transform -1 0 7268 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1649977179
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1649977179
transform -1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1649977179
transform 1 0 2208 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 9108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 10304 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 12880 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 7912 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 11132 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 13156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 7912 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 12236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 13984 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 12052 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 9844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 15640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 10120 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform 1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 14628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform 1 0 15732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 6164 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3036 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 1932 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 1748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 9384 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 9936 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6900 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 7636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 2576 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 2208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 8740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7544 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 5428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3312 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4048 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 6532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 5336 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 6256 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14444 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 16284 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 18400 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16744 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 16560 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17204 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16008 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16192 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 16468 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 15916 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14168 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 16560 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 13892 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 15456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 13984 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 13064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15272 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14168 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14536 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16928 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1649977179
transform 1 0 2760 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2208 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1649977179
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91
timestamp 1649977179
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95
timestamp 1649977179
transform 1 0 9844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_105
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_158
timestamp 1649977179
transform 1 0 15640 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1649977179
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_177
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_186
timestamp 1649977179
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_12
timestamp 1649977179
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_45
timestamp 1649977179
transform 1 0 5244 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_84
timestamp 1649977179
transform 1 0 8832 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_126
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1649977179
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1649977179
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_45
timestamp 1649977179
transform 1 0 5244 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_52
timestamp 1649977179
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 1649977179
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_90
timestamp 1649977179
transform 1 0 9384 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_100 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10304 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_125
timestamp 1649977179
transform 1 0 12604 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_128
timestamp 1649977179
transform 1 0 12880 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_137
timestamp 1649977179
transform 1 0 13708 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154
timestamp 1649977179
transform 1 0 15272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_158
timestamp 1649977179
transform 1 0 15640 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_174
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_186
timestamp 1649977179
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_24
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_36
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_48
timestamp 1649977179
transform 1 0 5520 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_59
timestamp 1649977179
transform 1 0 6532 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_71
timestamp 1649977179
transform 1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_115
timestamp 1649977179
transform 1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1649977179
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_135
timestamp 1649977179
transform 1 0 13524 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1649977179
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_177
timestamp 1649977179
transform 1 0 17388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_185
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_23
timestamp 1649977179
transform 1 0 3220 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_46
timestamp 1649977179
transform 1 0 5336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_69
timestamp 1649977179
transform 1 0 7452 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_73
timestamp 1649977179
transform 1 0 7820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_76
timestamp 1649977179
transform 1 0 8096 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_119
timestamp 1649977179
transform 1 0 12052 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_147
timestamp 1649977179
transform 1 0 14628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_169
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_184
timestamp 1649977179
transform 1 0 18032 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_25
timestamp 1649977179
transform 1 0 3404 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_85
timestamp 1649977179
transform 1 0 8924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_106
timestamp 1649977179
transform 1 0 10856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_126
timestamp 1649977179
transform 1 0 12696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_175
timestamp 1649977179
transform 1 0 17204 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_185
timestamp 1649977179
transform 1 0 18124 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1649977179
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_33
timestamp 1649977179
transform 1 0 4140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_64
timestamp 1649977179
transform 1 0 6992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_78
timestamp 1649977179
transform 1 0 8280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_94
timestamp 1649977179
transform 1 0 9752 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_156
timestamp 1649977179
transform 1 0 15456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_179
timestamp 1649977179
transform 1 0 17572 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_75
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_83
timestamp 1649977179
transform 1 0 8740 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_100
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_133
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_173
timestamp 1649977179
transform 1 0 17020 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 1649977179
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1649977179
transform 1 0 4324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_52
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1649977179
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_156
timestamp 1649977179
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_179
timestamp 1649977179
transform 1 0 17572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_183
timestamp 1649977179
transform 1 0 17940 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_77
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_85
timestamp 1649977179
transform 1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 1649977179
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_135
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_159
timestamp 1649977179
transform 1 0 15732 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_165
timestamp 1649977179
transform 1 0 16284 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_5
timestamp 1649977179
transform 1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_20
timestamp 1649977179
transform 1 0 2944 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1649977179
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_61
timestamp 1649977179
transform 1 0 6716 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1649977179
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_101
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_118
timestamp 1649977179
transform 1 0 11960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1649977179
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_158
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_170
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_33
timestamp 1649977179
transform 1 0 4140 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_73
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_85
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_102
timestamp 1649977179
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_145
timestamp 1649977179
transform 1 0 14444 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_177
timestamp 1649977179
transform 1 0 17388 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_184
timestamp 1649977179
transform 1 0 18032 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_63
timestamp 1649977179
transform 1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_67
timestamp 1649977179
transform 1 0 7268 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_114
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_155
timestamp 1649977179
transform 1 0 15364 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_167
timestamp 1649977179
transform 1 0 16468 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_175
timestamp 1649977179
transform 1 0 17204 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1649977179
transform 1 0 17848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1649977179
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_11
timestamp 1649977179
transform 1 0 2116 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_21
timestamp 1649977179
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_33
timestamp 1649977179
transform 1 0 4140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_65
timestamp 1649977179
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_97
timestamp 1649977179
transform 1 0 10028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_133
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_145
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_153
timestamp 1649977179
transform 1 0 15180 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_156
timestamp 1649977179
transform 1 0 15456 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_177
timestamp 1649977179
transform 1 0 17388 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_22
timestamp 1649977179
transform 1 0 3128 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1649977179
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1649977179
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_102
timestamp 1649977179
transform 1 0 10488 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_110
timestamp 1649977179
transform 1 0 11224 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_128
timestamp 1649977179
transform 1 0 12880 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_179
timestamp 1649977179
transform 1 0 17572 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_186
timestamp 1649977179
transform 1 0 18216 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1649977179
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_34
timestamp 1649977179
transform 1 0 4232 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_61
timestamp 1649977179
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_94
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_156
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_186
timestamp 1649977179
transform 1 0 18216 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1649977179
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_69
timestamp 1649977179
transform 1 0 7452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_98
timestamp 1649977179
transform 1 0 10120 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_110
timestamp 1649977179
transform 1 0 11224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_114
timestamp 1649977179
transform 1 0 11592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_159
timestamp 1649977179
transform 1 0 15732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_181
timestamp 1649977179
transform 1 0 17756 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_19
timestamp 1649977179
transform 1 0 2852 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1649977179
transform 1 0 3772 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_40
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_44
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_59
timestamp 1649977179
transform 1 0 6532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_103
timestamp 1649977179
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_119
timestamp 1649977179
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_133
timestamp 1649977179
transform 1 0 13340 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_174
timestamp 1649977179
transform 1 0 17112 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_186
timestamp 1649977179
transform 1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_13
timestamp 1649977179
transform 1 0 2300 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_104
timestamp 1649977179
transform 1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_115
timestamp 1649977179
transform 1 0 11684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_150
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_156
timestamp 1649977179
transform 1 0 15456 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_168
timestamp 1649977179
transform 1 0 16560 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_176
timestamp 1649977179
transform 1 0 17296 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_185
timestamp 1649977179
transform 1 0 18124 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_19
timestamp 1649977179
transform 1 0 2852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_23
timestamp 1649977179
transform 1 0 3220 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_37
timestamp 1649977179
transform 1 0 4508 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_49
timestamp 1649977179
transform 1 0 5612 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1649977179
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1649977179
transform 1 0 6624 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_65
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_77
timestamp 1649977179
transform 1 0 8188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1649977179
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_127
timestamp 1649977179
transform 1 0 12788 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_150
timestamp 1649977179
transform 1 0 14904 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_73
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1649977179
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_99
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_130
timestamp 1649977179
transform 1 0 13064 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_136
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_73
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_88
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_94
timestamp 1649977179
transform 1 0 9752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_101
timestamp 1649977179
transform 1 0 10396 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_107
timestamp 1649977179
transform 1 0 10948 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_118
timestamp 1649977179
transform 1 0 11960 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_128
timestamp 1649977179
transform 1 0 12880 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_142
timestamp 1649977179
transform 1 0 14168 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_154
timestamp 1649977179
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_57
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_69
timestamp 1649977179
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_113
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_125
timestamp 1649977179
transform 1 0 12604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1649977179
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_169
timestamp 1649977179
transform 1 0 16652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_181
timestamp 1649977179
transform 1 0 17756 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _09_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _10_
timestamp 1649977179
transform -1 0 6624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _11_
timestamp 1649977179
transform -1 0 3128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _12_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _13_
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _14_
timestamp 1649977179
transform -1 0 9660 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _15_
timestamp 1649977179
transform -1 0 17020 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1649977179
transform 1 0 12604 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1649977179
transform -1 0 15272 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _18_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1649977179
transform -1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1649977179
transform -1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1649977179
transform -1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1649977179
transform -1 0 2116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1649977179
transform -1 0 2576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1649977179
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1649977179
transform -1 0 3036 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1649977179
transform -1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1649977179
transform -1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1649977179
transform -1 0 2116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1649977179
transform -1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1649977179
transform -1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1649977179
transform -1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1649977179
transform -1 0 2116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1649977179
transform -1 0 2024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1649977179
transform -1 0 2116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1649977179
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1649977179
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1649977179
transform 1 0 17848 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1649977179
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1649977179
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1649977179
transform 1 0 17664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1649977179
transform 1 0 17756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1649977179
transform 1 0 17020 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1649977179
transform 1 0 17848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1649977179
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1649977179
transform 1 0 17480 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1649977179
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1649977179
transform 1 0 17848 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1649977179
transform 1 0 17848 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1649977179
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1649977179
transform 1 0 17848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1649977179
transform -1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1649977179
transform -1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1649977179
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1649977179
transform -1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1649977179
transform -1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1649977179
transform -1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1649977179
transform -1 0 10764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1649977179
transform -1 0 10856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1649977179
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1649977179
transform 1 0 16008 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1649977179
transform 1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1649977179
transform -1 0 13616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1649977179
transform -1 0 12880 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1649977179
transform -1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1649977179
transform -1 0 15272 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1649977179
transform -1 0 8464 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1649977179
transform -1 0 8832 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1649977179
transform -1 0 7636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1649977179
transform -1 0 11408 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1649977179
transform -1 0 10212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1649977179
transform -1 0 7084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1649977179
transform -1 0 3036 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1649977179
transform -1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1649977179
transform -1 0 2208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7636 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8924 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 7636 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10304 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform -1 0 10488 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 8924 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8004 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform -1 0 7912 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8188 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 11776 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 8096 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 10120 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6900 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 12420 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform -1 0 9752 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 10856 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 9016 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10672 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 12788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 13064 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 10028 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 12144 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9292 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 14168 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 10304 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 14720 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13892 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 14904 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 15916 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12420 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 4508 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4416 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11592 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10488 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9752 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7820 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5980 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5428 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4508 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5428 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8004 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5888 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 5980 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4508 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6256 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 8556 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11684 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12880 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6808 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10488 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13432 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13340 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12052 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3036 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 3588 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 1932 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3128 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2208 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2300 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2116 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2208 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1472 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9568 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8740 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7728 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6808 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6624 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5152 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3864 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1649977179
transform 1 0 3496 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3036 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2576 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2392 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3220 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1840 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2024 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1472 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6900 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7728 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6072 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4416 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3496 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3680 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2576 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6164 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5336 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6440 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5336 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13616 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12788 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16560 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16928 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16100 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8740 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9200 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8740 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7268 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15548 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16376 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15180 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15180 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16560 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14352 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15732 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 13524 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13892 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13156 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13064 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11776 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11592 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11960 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10948 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10856 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15364 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15456 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15180 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15640 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15456 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14904 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14076 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1649977179
transform -1 0 2208 0 1 3264
box -38 -48 590 592
<< labels >>
flabel metal2 s 7378 16400 7434 17200 0 FreeSans 224 90 0 0 IO_ISOL_N
port 0 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 SC_IN_BOT
port 1 nsew signal input
flabel metal2 s 6090 16400 6146 17200 0 FreeSans 224 90 0 0 SC_IN_TOP
port 2 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 3 nsew signal tristate
flabel metal2 s 6734 16400 6790 17200 0 FreeSans 224 90 0 0 SC_OUT_TOP
port 4 nsew signal tristate
flabel metal4 s 5392 2128 5712 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 9840 2128 10160 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 14288 2128 14608 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 3168 2128 3488 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 7616 2128 7936 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 12064 2128 12384 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 16512 2128 16832 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 bottom_grid_pin_0_
port 7 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 bottom_grid_pin_10_
port 8 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_grid_pin_12_
port 9 nsew signal tristate
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 bottom_grid_pin_14_
port 10 nsew signal tristate
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 bottom_grid_pin_16_
port 11 nsew signal tristate
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 bottom_grid_pin_2_
port 12 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 bottom_grid_pin_4_
port 13 nsew signal tristate
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 bottom_grid_pin_6_
port 14 nsew signal tristate
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 bottom_grid_pin_8_
port 15 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 ccff_head
port 16 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 ccff_tail
port 17 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 18 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 19 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 20 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 21 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 22 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 23 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 24 nsew signal input
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 25 nsew signal input
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 26 nsew signal input
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 27 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 28 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 29 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 30 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 31 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 32 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 33 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 34 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 35 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 36 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 37 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 38 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 39 nsew signal tristate
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 40 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 41 nsew signal tristate
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 42 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 43 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 44 nsew signal tristate
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 45 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 46 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 47 nsew signal tristate
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 48 nsew signal tristate
flabel metal3 s 0 1096 800 1216 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 49 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 50 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 51 nsew signal tristate
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 52 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 53 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 54 nsew signal tristate
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 55 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 56 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 57 nsew signal tristate
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 58 nsew signal input
flabel metal3 s 19200 12792 20000 12912 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 59 nsew signal input
flabel metal3 s 19200 13200 20000 13320 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 60 nsew signal input
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 61 nsew signal input
flabel metal3 s 19200 14016 20000 14136 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 62 nsew signal input
flabel metal3 s 19200 14424 20000 14544 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 63 nsew signal input
flabel metal3 s 19200 14832 20000 14952 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 64 nsew signal input
flabel metal3 s 19200 15240 20000 15360 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 65 nsew signal input
flabel metal3 s 19200 15648 20000 15768 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 66 nsew signal input
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 67 nsew signal input
flabel metal3 s 19200 16464 20000 16584 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 68 nsew signal input
flabel metal3 s 19200 9120 20000 9240 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 69 nsew signal input
flabel metal3 s 19200 9528 20000 9648 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 70 nsew signal input
flabel metal3 s 19200 9936 20000 10056 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 71 nsew signal input
flabel metal3 s 19200 10344 20000 10464 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 72 nsew signal input
flabel metal3 s 19200 10752 20000 10872 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 73 nsew signal input
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 74 nsew signal input
flabel metal3 s 19200 11568 20000 11688 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 75 nsew signal input
flabel metal3 s 19200 11976 20000 12096 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 76 nsew signal input
flabel metal3 s 19200 12384 20000 12504 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 77 nsew signal input
flabel metal3 s 19200 552 20000 672 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 78 nsew signal tristate
flabel metal3 s 19200 4632 20000 4752 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 79 nsew signal tristate
flabel metal3 s 19200 5040 20000 5160 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 80 nsew signal tristate
flabel metal3 s 19200 5448 20000 5568 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 81 nsew signal tristate
flabel metal3 s 19200 5856 20000 5976 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 82 nsew signal tristate
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 83 nsew signal tristate
flabel metal3 s 19200 6672 20000 6792 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 84 nsew signal tristate
flabel metal3 s 19200 7080 20000 7200 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 85 nsew signal tristate
flabel metal3 s 19200 7488 20000 7608 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 86 nsew signal tristate
flabel metal3 s 19200 7896 20000 8016 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 87 nsew signal tristate
flabel metal3 s 19200 8304 20000 8424 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 88 nsew signal tristate
flabel metal3 s 19200 960 20000 1080 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 89 nsew signal tristate
flabel metal3 s 19200 1368 20000 1488 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 90 nsew signal tristate
flabel metal3 s 19200 1776 20000 1896 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 91 nsew signal tristate
flabel metal3 s 19200 2184 20000 2304 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 92 nsew signal tristate
flabel metal3 s 19200 2592 20000 2712 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 93 nsew signal tristate
flabel metal3 s 19200 3000 20000 3120 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 94 nsew signal tristate
flabel metal3 s 19200 3408 20000 3528 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 95 nsew signal tristate
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 96 nsew signal tristate
flabel metal3 s 19200 4224 20000 4344 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 97 nsew signal tristate
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
port 98 nsew signal tristate
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
port 99 nsew signal tristate
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
port 100 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
port 101 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
port 102 nsew signal tristate
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
port 103 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
port 104 nsew signal tristate
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
port 105 nsew signal tristate
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
port 106 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
port 107 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
port 108 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
port 109 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
port 110 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
port 111 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
port 112 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
port 113 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
port 114 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
port 115 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
port 116 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
port 117 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
port 118 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
port 119 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
port 120 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
port 121 nsew signal tristate
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
port 122 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
port 123 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
port 124 nsew signal tristate
flabel metal2 s 8022 16400 8078 17200 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 125 nsew signal input
flabel metal3 s 0 280 800 400 0 FreeSans 480 0 0 0 prog_clk_0_W_out
port 126 nsew signal tristate
flabel metal2 s 8666 16400 8722 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_0_
port 127 nsew signal input
flabel metal2 s 11886 16400 11942 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_10_
port 128 nsew signal input
flabel metal2 s 19614 16400 19670 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_11_lower
port 129 nsew signal tristate
flabel metal2 s 3514 16400 3570 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_11_upper
port 130 nsew signal tristate
flabel metal2 s 12530 16400 12586 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_12_
port 131 nsew signal input
flabel metal2 s 14462 16400 14518 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_13_lower
port 132 nsew signal tristate
flabel metal2 s 4158 16400 4214 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_13_upper
port 133 nsew signal tristate
flabel metal2 s 13174 16400 13230 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_14_
port 134 nsew signal input
flabel metal2 s 15106 16400 15162 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_15_lower
port 135 nsew signal tristate
flabel metal2 s 4802 16400 4858 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_15_upper
port 136 nsew signal tristate
flabel metal2 s 13818 16400 13874 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_16_
port 137 nsew signal input
flabel metal2 s 15750 16400 15806 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_17_lower
port 138 nsew signal tristate
flabel metal2 s 5446 16400 5502 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_17_upper
port 139 nsew signal tristate
flabel metal2 s 16394 16400 16450 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_1_lower
port 140 nsew signal tristate
flabel metal2 s 294 16400 350 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_1_upper
port 141 nsew signal tristate
flabel metal2 s 9310 16400 9366 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_2_
port 142 nsew signal input
flabel metal2 s 17038 16400 17094 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_3_lower
port 143 nsew signal tristate
flabel metal2 s 938 16400 994 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_3_upper
port 144 nsew signal tristate
flabel metal2 s 9954 16400 10010 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_4_
port 145 nsew signal input
flabel metal2 s 17682 16400 17738 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_5_lower
port 146 nsew signal tristate
flabel metal2 s 1582 16400 1638 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_5_upper
port 147 nsew signal tristate
flabel metal2 s 10598 16400 10654 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_6_
port 148 nsew signal input
flabel metal2 s 18326 16400 18382 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_7_lower
port 149 nsew signal tristate
flabel metal2 s 2226 16400 2282 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_7_upper
port 150 nsew signal tristate
flabel metal2 s 11242 16400 11298 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_8_
port 151 nsew signal input
flabel metal2 s 18970 16400 19026 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_9_lower
port 152 nsew signal tristate
flabel metal2 s 2870 16400 2926 17200 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_9_upper
port 153 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
