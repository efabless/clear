magic
tech sky130A
magscale 1 2
timestamp 1656242629
<< viali >>
rect 1869 20553 1903 20587
rect 2237 20553 2271 20587
rect 10333 20553 10367 20587
rect 11897 20553 11931 20587
rect 12265 20553 12299 20587
rect 12633 20553 12667 20587
rect 12909 20553 12943 20587
rect 13369 20553 13403 20587
rect 13645 20553 13679 20587
rect 14289 20553 14323 20587
rect 15025 20553 15059 20587
rect 15393 20553 15427 20587
rect 16129 20553 16163 20587
rect 16865 20553 16899 20587
rect 17233 20553 17267 20587
rect 17969 20553 18003 20587
rect 19533 20553 19567 20587
rect 19993 20553 20027 20587
rect 20361 20553 20395 20587
rect 21465 20553 21499 20587
rect 2697 20485 2731 20519
rect 3065 20485 3099 20519
rect 9045 20485 9079 20519
rect 1685 20417 1719 20451
rect 2053 20417 2087 20451
rect 2421 20417 2455 20451
rect 3525 20417 3559 20451
rect 4629 20417 4663 20451
rect 4721 20417 4755 20451
rect 5089 20417 5123 20451
rect 6561 20417 6595 20451
rect 6929 20417 6963 20451
rect 7021 20417 7055 20451
rect 7573 20417 7607 20451
rect 7757 20417 7791 20451
rect 8493 20417 8527 20451
rect 9965 20417 9999 20451
rect 10149 20417 10183 20451
rect 10517 20417 10551 20451
rect 11713 20417 11747 20451
rect 12081 20417 12115 20451
rect 12449 20417 12483 20451
rect 13093 20417 13127 20451
rect 13185 20417 13219 20451
rect 13829 20417 13863 20451
rect 14105 20417 14139 20451
rect 14473 20417 14507 20451
rect 14841 20417 14875 20451
rect 15209 20417 15243 20451
rect 15577 20417 15611 20451
rect 15945 20417 15979 20451
rect 16313 20417 16347 20451
rect 16681 20417 16715 20451
rect 17049 20417 17083 20451
rect 17417 20417 17451 20451
rect 17785 20417 17819 20451
rect 18153 20417 18187 20451
rect 18521 20417 18555 20451
rect 18889 20417 18923 20451
rect 19717 20417 19751 20451
rect 19809 20417 19843 20451
rect 20177 20417 20211 20451
rect 20545 20417 20579 20451
rect 20913 20417 20947 20451
rect 21281 20417 21315 20451
rect 4353 20349 4387 20383
rect 5917 20349 5951 20383
rect 6193 20349 6227 20383
rect 6745 20349 6779 20383
rect 8769 20349 8803 20383
rect 9689 20349 9723 20383
rect 10793 20349 10827 20383
rect 4905 20281 4939 20315
rect 5273 20281 5307 20315
rect 7389 20281 7423 20315
rect 14657 20281 14691 20315
rect 15761 20281 15795 20315
rect 17601 20281 17635 20315
rect 18705 20281 18739 20315
rect 19073 20281 19107 20315
rect 19349 20281 19383 20315
rect 20729 20281 20763 20315
rect 1501 20213 1535 20247
rect 2789 20213 2823 20247
rect 3157 20213 3191 20247
rect 3433 20213 3467 20247
rect 6377 20213 6411 20247
rect 11621 20213 11655 20247
rect 16497 20213 16531 20247
rect 18337 20213 18371 20247
rect 21097 20213 21131 20247
rect 2237 20009 2271 20043
rect 2605 20009 2639 20043
rect 4077 20009 4111 20043
rect 7113 20009 7147 20043
rect 9137 20009 9171 20043
rect 11437 20009 11471 20043
rect 12081 20009 12115 20043
rect 12541 20009 12575 20043
rect 13093 20009 13127 20043
rect 13369 20009 13403 20043
rect 13645 20009 13679 20043
rect 14289 20009 14323 20043
rect 14657 20009 14691 20043
rect 14933 20009 14967 20043
rect 15209 20009 15243 20043
rect 15761 20009 15795 20043
rect 16037 20009 16071 20043
rect 16773 20009 16807 20043
rect 17417 20009 17451 20043
rect 18245 20009 18279 20043
rect 18429 20009 18463 20043
rect 18705 20009 18739 20043
rect 19533 20009 19567 20043
rect 20545 20009 20579 20043
rect 2881 19941 2915 19975
rect 3249 19941 3283 19975
rect 3617 19941 3651 19975
rect 9597 19941 9631 19975
rect 12817 19941 12851 19975
rect 13737 19941 13771 19975
rect 15485 19941 15519 19975
rect 17049 19941 17083 19975
rect 17785 19941 17819 19975
rect 7849 19873 7883 19907
rect 8217 19873 8251 19907
rect 10977 19873 11011 19907
rect 12173 19873 12207 19907
rect 18981 19873 19015 19907
rect 1685 19805 1719 19839
rect 2053 19805 2087 19839
rect 2421 19805 2455 19839
rect 2697 19805 2731 19839
rect 3065 19805 3099 19839
rect 4261 19805 4295 19839
rect 5733 19805 5767 19839
rect 8953 19805 8987 19839
rect 11069 19805 11103 19839
rect 11621 19805 11655 19839
rect 11897 19805 11931 19839
rect 12357 19781 12391 19815
rect 12625 19805 12659 19839
rect 12909 19805 12943 19839
rect 13185 19805 13219 19839
rect 13461 19805 13495 19839
rect 13921 19805 13955 19839
rect 14105 19805 14139 19839
rect 14473 19805 14507 19839
rect 14749 19805 14783 19839
rect 15025 19805 15059 19839
rect 15301 19805 15335 19839
rect 15577 19805 15611 19839
rect 15853 19805 15887 19839
rect 16129 19805 16163 19839
rect 16497 19805 16531 19839
rect 16957 19805 16991 19839
rect 17233 19805 17267 19839
rect 17693 19805 17727 19839
rect 17969 19805 18003 19839
rect 18061 19805 18095 19839
rect 18613 19805 18647 19839
rect 18889 19805 18923 19839
rect 19441 19805 19475 19839
rect 20177 19805 20211 19839
rect 20361 19805 20395 19839
rect 20729 19805 20763 19839
rect 21281 19805 21315 19839
rect 3433 19737 3467 19771
rect 3985 19737 4019 19771
rect 4528 19737 4562 19771
rect 5978 19737 6012 19771
rect 8401 19737 8435 19771
rect 9229 19737 9263 19771
rect 9413 19737 9447 19771
rect 10710 19737 10744 19771
rect 19901 19737 19935 19771
rect 21005 19737 21039 19771
rect 1501 19669 1535 19703
rect 1869 19669 1903 19703
rect 5641 19669 5675 19703
rect 7205 19669 7239 19703
rect 7573 19669 7607 19703
rect 7665 19669 7699 19703
rect 8309 19669 8343 19703
rect 8769 19669 8803 19703
rect 11253 19669 11287 19703
rect 11805 19669 11839 19703
rect 16313 19669 16347 19703
rect 16681 19669 16715 19703
rect 17509 19669 17543 19703
rect 19257 19669 19291 19703
rect 21465 19669 21499 19703
rect 1869 19465 1903 19499
rect 2329 19465 2363 19499
rect 3709 19465 3743 19499
rect 4905 19465 4939 19499
rect 5365 19465 5399 19499
rect 5733 19465 5767 19499
rect 5825 19465 5859 19499
rect 6193 19465 6227 19499
rect 6745 19465 6779 19499
rect 6837 19465 6871 19499
rect 8677 19465 8711 19499
rect 10517 19465 10551 19499
rect 10977 19465 11011 19499
rect 13001 19465 13035 19499
rect 14013 19465 14047 19499
rect 14381 19465 14415 19499
rect 16497 19465 16531 19499
rect 17233 19465 17267 19499
rect 18153 19465 18187 19499
rect 18429 19465 18463 19499
rect 18797 19465 18831 19499
rect 19073 19465 19107 19499
rect 19809 19465 19843 19499
rect 20177 19465 20211 19499
rect 9014 19397 9048 19431
rect 11161 19397 11195 19431
rect 14933 19397 14967 19431
rect 1685 19329 1719 19363
rect 2053 19329 2087 19363
rect 2145 19329 2179 19363
rect 2789 19329 2823 19363
rect 3617 19329 3651 19363
rect 4353 19329 4387 19363
rect 4997 19329 5031 19363
rect 7564 19329 7598 19363
rect 8769 19329 8803 19363
rect 10609 19329 10643 19363
rect 11529 19329 11563 19363
rect 11796 19329 11830 19363
rect 13185 19329 13219 19363
rect 14197 19329 14231 19363
rect 14473 19329 14507 19363
rect 16313 19329 16347 19363
rect 17049 19329 17083 19363
rect 17969 19329 18003 19363
rect 18245 19329 18279 19363
rect 18521 19329 18555 19363
rect 18981 19329 19015 19363
rect 19257 19329 19291 19363
rect 19349 19329 19383 19363
rect 19625 19329 19659 19363
rect 19993 19329 20027 19363
rect 20361 19329 20395 19363
rect 20729 19329 20763 19363
rect 21281 19329 21315 19363
rect 2605 19261 2639 19295
rect 2697 19261 2731 19295
rect 3893 19261 3927 19295
rect 4813 19261 4847 19295
rect 5549 19261 5583 19295
rect 6653 19261 6687 19295
rect 7297 19261 7331 19295
rect 10425 19261 10459 19295
rect 17877 19261 17911 19295
rect 20913 19261 20947 19295
rect 4169 19193 4203 19227
rect 7205 19193 7239 19227
rect 10149 19193 10183 19227
rect 13461 19193 13495 19227
rect 14657 19193 14691 19227
rect 15301 19193 15335 19227
rect 18705 19193 18739 19227
rect 19533 19193 19567 19227
rect 20545 19193 20579 19227
rect 1501 19125 1535 19159
rect 3157 19125 3191 19159
rect 3249 19125 3283 19159
rect 4445 19125 4479 19159
rect 11253 19125 11287 19159
rect 12909 19125 12943 19159
rect 13277 19125 13311 19159
rect 13645 19125 13679 19159
rect 14841 19125 14875 19159
rect 15209 19125 15243 19159
rect 15485 19125 15519 19159
rect 15669 19125 15703 19159
rect 16129 19125 16163 19159
rect 16865 19125 16899 19159
rect 21465 19125 21499 19159
rect 2145 18921 2179 18955
rect 2789 18921 2823 18955
rect 7849 18921 7883 18955
rect 9689 18921 9723 18955
rect 10241 18921 10275 18955
rect 10517 18921 10551 18955
rect 13737 18921 13771 18955
rect 19349 18921 19383 18955
rect 19625 18921 19659 18955
rect 19901 18921 19935 18955
rect 2421 18853 2455 18887
rect 3893 18853 3927 18887
rect 12909 18853 12943 18887
rect 19073 18853 19107 18887
rect 19993 18853 20027 18887
rect 20269 18853 20303 18887
rect 3341 18785 3375 18819
rect 3433 18785 3467 18819
rect 4169 18785 4203 18819
rect 6193 18785 6227 18819
rect 6469 18785 6503 18819
rect 8493 18785 8527 18819
rect 9045 18785 9079 18819
rect 11989 18785 12023 18819
rect 12173 18785 12207 18819
rect 13461 18785 13495 18819
rect 14289 18785 14323 18819
rect 18797 18785 18831 18819
rect 1685 18717 1719 18751
rect 1777 18717 1811 18751
rect 2329 18717 2363 18751
rect 2605 18717 2639 18751
rect 3249 18717 3283 18751
rect 4077 18717 4111 18751
rect 6101 18717 6135 18751
rect 6736 18717 6770 18751
rect 9965 18717 9999 18751
rect 10333 18717 10367 18751
rect 12357 18717 12391 18751
rect 14381 18717 14415 18751
rect 18889 18717 18923 18751
rect 19441 18717 19475 18751
rect 19717 18693 19751 18727
rect 20177 18717 20211 18751
rect 20453 18717 20487 18751
rect 20637 18717 20671 18751
rect 21281 18717 21315 18751
rect 4436 18649 4470 18683
rect 8401 18649 8435 18683
rect 9781 18649 9815 18683
rect 11744 18649 11778 18683
rect 13369 18649 13403 18683
rect 14473 18649 14507 18683
rect 18613 18649 18647 18683
rect 20913 18649 20947 18683
rect 1501 18581 1535 18615
rect 1961 18581 1995 18615
rect 2881 18581 2915 18615
rect 5549 18581 5583 18615
rect 5641 18581 5675 18615
rect 6009 18581 6043 18615
rect 7941 18581 7975 18615
rect 8309 18581 8343 18615
rect 9229 18581 9263 18615
rect 9321 18581 9355 18615
rect 10609 18581 10643 18615
rect 12449 18581 12483 18615
rect 12817 18581 12851 18615
rect 13277 18581 13311 18615
rect 14841 18581 14875 18615
rect 18429 18581 18463 18615
rect 21465 18581 21499 18615
rect 1777 18377 1811 18411
rect 4905 18377 4939 18411
rect 6193 18377 6227 18411
rect 6377 18377 6411 18411
rect 7389 18377 7423 18411
rect 7757 18377 7791 18411
rect 8217 18377 8251 18411
rect 8677 18377 8711 18411
rect 9137 18377 9171 18411
rect 11345 18377 11379 18411
rect 12633 18377 12667 18411
rect 19625 18377 19659 18411
rect 3166 18309 3200 18343
rect 3801 18309 3835 18343
rect 5733 18309 5767 18343
rect 5825 18309 5859 18343
rect 12265 18309 12299 18343
rect 13360 18309 13394 18343
rect 1685 18241 1719 18275
rect 1961 18241 1995 18275
rect 3433 18241 3467 18275
rect 3893 18241 3927 18275
rect 4353 18241 4387 18275
rect 4997 18241 5031 18275
rect 6745 18241 6779 18275
rect 7205 18241 7239 18275
rect 7849 18241 7883 18275
rect 9505 18241 9539 18275
rect 10149 18241 10183 18275
rect 10333 18241 10367 18275
rect 10977 18241 11011 18275
rect 14749 18241 14783 18275
rect 19441 18241 19475 18275
rect 19717 18241 19751 18275
rect 19993 18241 20027 18275
rect 20361 18241 20395 18275
rect 20637 18241 20671 18275
rect 20913 18241 20947 18275
rect 21281 18241 21315 18275
rect 3617 18173 3651 18207
rect 4721 18173 4755 18207
rect 5641 18173 5675 18207
rect 6837 18173 6871 18207
rect 6929 18173 6963 18207
rect 7573 18173 7607 18207
rect 8401 18173 8435 18207
rect 8585 18173 8619 18207
rect 9597 18173 9631 18207
rect 9689 18173 9723 18207
rect 10701 18173 10735 18207
rect 10885 18173 10919 18207
rect 11529 18173 11563 18207
rect 11989 18173 12023 18207
rect 12173 18173 12207 18207
rect 12725 18173 12759 18207
rect 13093 18173 13127 18207
rect 4261 18105 4295 18139
rect 9045 18105 9079 18139
rect 9965 18105 9999 18139
rect 10517 18105 10551 18139
rect 14565 18105 14599 18139
rect 18981 18105 19015 18139
rect 19165 18105 19199 18139
rect 21097 18105 21131 18139
rect 1501 18037 1535 18071
rect 2053 18037 2087 18071
rect 4537 18037 4571 18071
rect 5365 18037 5399 18071
rect 11713 18037 11747 18071
rect 14473 18037 14507 18071
rect 15577 18037 15611 18071
rect 19349 18037 19383 18071
rect 19901 18037 19935 18071
rect 20177 18037 20211 18071
rect 20545 18037 20579 18071
rect 20821 18037 20855 18071
rect 21465 18037 21499 18071
rect 1869 17833 1903 17867
rect 3617 17833 3651 17867
rect 4629 17833 4663 17867
rect 6101 17833 6135 17867
rect 8769 17833 8803 17867
rect 10149 17833 10183 17867
rect 10425 17833 10459 17867
rect 11069 17833 11103 17867
rect 12265 17833 12299 17867
rect 20269 17833 20303 17867
rect 21189 17833 21223 17867
rect 9965 17765 9999 17799
rect 13277 17765 13311 17799
rect 20729 17765 20763 17799
rect 4077 17697 4111 17731
rect 6745 17697 6779 17731
rect 7205 17697 7239 17731
rect 8217 17697 8251 17731
rect 9413 17697 9447 17731
rect 9597 17697 9631 17731
rect 11529 17697 11563 17731
rect 12817 17697 12851 17731
rect 16313 17697 16347 17731
rect 1685 17629 1719 17663
rect 2053 17629 2087 17663
rect 2237 17629 2271 17663
rect 4169 17629 4203 17663
rect 4721 17629 4755 17663
rect 9781 17629 9815 17663
rect 10333 17629 10367 17663
rect 10609 17629 10643 17663
rect 11345 17629 11379 17663
rect 12633 17629 12667 17663
rect 14197 17629 14231 17663
rect 14464 17629 14498 17663
rect 19717 17629 19751 17663
rect 20085 17629 20119 17663
rect 20545 17629 20579 17663
rect 20913 17629 20947 17663
rect 21005 17629 21039 17663
rect 21281 17629 21315 17663
rect 2504 17561 2538 17595
rect 4988 17561 5022 17595
rect 6561 17561 6595 17595
rect 7389 17561 7423 17595
rect 11713 17561 11747 17595
rect 13461 17561 13495 17595
rect 19901 17561 19935 17595
rect 1501 17493 1535 17527
rect 4261 17493 4295 17527
rect 6193 17493 6227 17527
rect 6653 17493 6687 17527
rect 7297 17493 7331 17527
rect 7757 17493 7791 17527
rect 7941 17493 7975 17527
rect 8309 17493 8343 17527
rect 8401 17493 8435 17527
rect 8953 17493 8987 17527
rect 9321 17493 9355 17527
rect 10701 17493 10735 17527
rect 10885 17493 10919 17527
rect 11805 17493 11839 17527
rect 12173 17493 12207 17527
rect 12725 17493 12759 17527
rect 13093 17493 13127 17527
rect 15577 17493 15611 17527
rect 15669 17493 15703 17527
rect 16037 17493 16071 17527
rect 16129 17493 16163 17527
rect 20361 17493 20395 17527
rect 21465 17493 21499 17527
rect 1869 17289 1903 17323
rect 2145 17289 2179 17323
rect 2697 17289 2731 17323
rect 3157 17289 3191 17323
rect 4629 17289 4663 17323
rect 5457 17289 5491 17323
rect 5917 17289 5951 17323
rect 6837 17289 6871 17323
rect 8217 17289 8251 17323
rect 9045 17289 9079 17323
rect 9505 17289 9539 17323
rect 11713 17289 11747 17323
rect 12081 17289 12115 17323
rect 13001 17289 13035 17323
rect 14197 17289 14231 17323
rect 14657 17289 14691 17323
rect 15761 17289 15795 17323
rect 19993 17289 20027 17323
rect 20729 17289 20763 17323
rect 21005 17289 21039 17323
rect 3494 17221 3528 17255
rect 6469 17221 6503 17255
rect 7297 17221 7331 17255
rect 7665 17221 7699 17255
rect 12909 17221 12943 17255
rect 14105 17221 14139 17255
rect 1685 17153 1719 17187
rect 2053 17153 2087 17187
rect 2329 17153 2363 17187
rect 2789 17153 2823 17187
rect 3249 17153 3283 17187
rect 4721 17153 4755 17187
rect 5181 17153 5215 17187
rect 5365 17153 5399 17187
rect 5825 17153 5859 17187
rect 7205 17153 7239 17187
rect 8585 17153 8619 17187
rect 8677 17153 8711 17187
rect 9413 17153 9447 17187
rect 10129 17153 10163 17187
rect 12173 17153 12207 17187
rect 13737 17153 13771 17187
rect 15025 17153 15059 17187
rect 15853 17153 15887 17187
rect 19809 17153 19843 17187
rect 20545 17153 20579 17187
rect 20821 17153 20855 17187
rect 21281 17153 21315 17187
rect 2605 17085 2639 17119
rect 6009 17085 6043 17119
rect 7481 17085 7515 17119
rect 7941 17085 7975 17119
rect 8861 17085 8895 17119
rect 9597 17085 9631 17119
rect 9873 17085 9907 17119
rect 11621 17085 11655 17119
rect 12265 17085 12299 17119
rect 13093 17085 13127 17119
rect 13921 17085 13955 17119
rect 15117 17085 15151 17119
rect 15209 17085 15243 17119
rect 15577 17085 15611 17119
rect 4905 17017 4939 17051
rect 6653 17017 6687 17051
rect 11253 17017 11287 17051
rect 14565 17017 14599 17051
rect 21189 17017 21223 17051
rect 1501 16949 1535 16983
rect 4997 16949 5031 16983
rect 8033 16949 8067 16983
rect 12541 16949 12575 16983
rect 13553 16949 13587 16983
rect 16221 16949 16255 16983
rect 20361 16949 20395 16983
rect 21465 16949 21499 16983
rect 2145 16745 2179 16779
rect 2789 16745 2823 16779
rect 5641 16745 5675 16779
rect 6653 16745 6687 16779
rect 7665 16745 7699 16779
rect 7849 16745 7883 16779
rect 8769 16745 8803 16779
rect 15577 16745 15611 16779
rect 16405 16745 16439 16779
rect 18429 16745 18463 16779
rect 19441 16745 19475 16779
rect 20821 16745 20855 16779
rect 5549 16677 5583 16711
rect 18245 16677 18279 16711
rect 2973 16609 3007 16643
rect 3157 16609 3191 16643
rect 6469 16609 6503 16643
rect 7113 16609 7147 16643
rect 7297 16609 7331 16643
rect 7573 16609 7607 16643
rect 8125 16609 8159 16643
rect 9321 16609 9355 16643
rect 9689 16609 9723 16643
rect 10885 16609 10919 16643
rect 11713 16609 11747 16643
rect 13921 16609 13955 16643
rect 14105 16609 14139 16643
rect 16037 16609 16071 16643
rect 16129 16609 16163 16643
rect 16957 16609 16991 16643
rect 17325 16609 17359 16643
rect 17509 16609 17543 16643
rect 18061 16609 18095 16643
rect 1685 16541 1719 16575
rect 2053 16541 2087 16575
rect 2329 16541 2363 16575
rect 2605 16541 2639 16575
rect 4169 16541 4203 16575
rect 4436 16541 4470 16575
rect 6193 16541 6227 16575
rect 16865 16541 16899 16575
rect 19257 16541 19291 16575
rect 20637 16541 20671 16575
rect 20913 16541 20947 16575
rect 21281 16541 21315 16575
rect 3249 16473 3283 16507
rect 3801 16473 3835 16507
rect 8401 16473 8435 16507
rect 8953 16473 8987 16507
rect 10793 16473 10827 16507
rect 11621 16473 11655 16507
rect 13676 16473 13710 16507
rect 14372 16473 14406 16507
rect 16773 16473 16807 16507
rect 1501 16405 1535 16439
rect 1869 16405 1903 16439
rect 2421 16405 2455 16439
rect 3617 16405 3651 16439
rect 5825 16405 5859 16439
rect 6285 16405 6319 16439
rect 7021 16405 7055 16439
rect 8309 16405 8343 16439
rect 9781 16405 9815 16439
rect 9873 16405 9907 16439
rect 10241 16405 10275 16439
rect 10333 16405 10367 16439
rect 10701 16405 10735 16439
rect 11161 16405 11195 16439
rect 11529 16405 11563 16439
rect 12081 16405 12115 16439
rect 12541 16405 12575 16439
rect 15485 16405 15519 16439
rect 15945 16405 15979 16439
rect 17601 16405 17635 16439
rect 17969 16405 18003 16439
rect 18613 16405 18647 16439
rect 20453 16405 20487 16439
rect 21097 16405 21131 16439
rect 21465 16405 21499 16439
rect 1869 16201 1903 16235
rect 2329 16201 2363 16235
rect 2697 16201 2731 16235
rect 3341 16201 3375 16235
rect 3709 16201 3743 16235
rect 4169 16201 4203 16235
rect 4629 16201 4663 16235
rect 6193 16201 6227 16235
rect 7113 16201 7147 16235
rect 8677 16201 8711 16235
rect 8953 16201 8987 16235
rect 9321 16201 9355 16235
rect 10793 16201 10827 16235
rect 13461 16201 13495 16235
rect 15025 16201 15059 16235
rect 15393 16201 15427 16235
rect 15853 16201 15887 16235
rect 16405 16201 16439 16235
rect 16681 16201 16715 16235
rect 17509 16201 17543 16235
rect 17969 16201 18003 16235
rect 18337 16201 18371 16235
rect 18797 16201 18831 16235
rect 20453 16201 20487 16235
rect 20729 16201 20763 16235
rect 21005 16201 21039 16235
rect 5733 16133 5767 16167
rect 6653 16133 6687 16167
rect 9045 16133 9079 16167
rect 13124 16133 13158 16167
rect 14657 16133 14691 16167
rect 18705 16133 18739 16167
rect 21097 16133 21131 16167
rect 1685 16065 1719 16099
rect 2053 16065 2087 16099
rect 2145 16065 2179 16099
rect 2513 16065 2547 16099
rect 4261 16065 4295 16099
rect 4997 16065 5031 16099
rect 5825 16065 5859 16099
rect 6377 16065 6411 16099
rect 7481 16065 7515 16099
rect 8125 16065 8159 16099
rect 8585 16065 8619 16099
rect 9669 16065 9703 16099
rect 11069 16065 11103 16099
rect 13369 16065 13403 16099
rect 13829 16065 13863 16099
rect 14565 16065 14599 16099
rect 15485 16065 15519 16099
rect 16129 16065 16163 16099
rect 17049 16065 17083 16099
rect 17877 16065 17911 16099
rect 20269 16065 20303 16099
rect 20545 16065 20579 16099
rect 20821 16065 20855 16099
rect 21281 16065 21315 16099
rect 3065 15997 3099 16031
rect 3249 15997 3283 16031
rect 4353 15997 4387 16031
rect 5089 15997 5123 16031
rect 5273 15997 5307 16031
rect 5641 15997 5675 16031
rect 7573 15997 7607 16031
rect 7665 15997 7699 16031
rect 9413 15997 9447 16031
rect 13921 15997 13955 16031
rect 14013 15997 14047 16031
rect 14473 15997 14507 16031
rect 15301 15997 15335 16031
rect 17141 15997 17175 16031
rect 17233 15997 17267 16031
rect 18061 15997 18095 16031
rect 18981 15997 19015 16031
rect 20177 15997 20211 16031
rect 3801 15929 3835 15963
rect 8033 15929 8067 15963
rect 1501 15861 1535 15895
rect 2881 15861 2915 15895
rect 6929 15861 6963 15895
rect 8401 15861 8435 15895
rect 10885 15861 10919 15895
rect 11253 15861 11287 15895
rect 11989 15861 12023 15895
rect 21465 15861 21499 15895
rect 1869 15657 1903 15691
rect 2145 15657 2179 15691
rect 2421 15657 2455 15691
rect 3157 15657 3191 15691
rect 3801 15657 3835 15691
rect 4629 15657 4663 15691
rect 4997 15657 5031 15691
rect 5641 15657 5675 15691
rect 6377 15657 6411 15691
rect 11897 15657 11931 15691
rect 13369 15657 13403 15691
rect 17049 15657 17083 15691
rect 19257 15657 19291 15691
rect 20729 15657 20763 15691
rect 6193 15589 6227 15623
rect 14657 15589 14691 15623
rect 20361 15589 20395 15623
rect 4353 15521 4387 15555
rect 5457 15521 5491 15555
rect 6009 15521 6043 15555
rect 7113 15521 7147 15555
rect 10517 15521 10551 15555
rect 12449 15521 12483 15555
rect 12633 15521 12667 15555
rect 14105 15521 14139 15555
rect 19809 15521 19843 15555
rect 1685 15453 1719 15487
rect 2053 15453 2087 15487
rect 2329 15453 2363 15487
rect 2605 15453 2639 15487
rect 2697 15453 2731 15487
rect 2973 15453 3007 15487
rect 3249 15453 3283 15487
rect 4813 15453 4847 15487
rect 5181 15453 5215 15487
rect 7389 15453 7423 15487
rect 8953 15453 8987 15487
rect 13829 15453 13863 15487
rect 15025 15453 15059 15487
rect 15485 15453 15519 15487
rect 15577 15453 15611 15487
rect 15844 15453 15878 15487
rect 18429 15453 18463 15487
rect 18981 15453 19015 15487
rect 19717 15453 19751 15487
rect 20085 15453 20119 15487
rect 20545 15453 20579 15487
rect 20821 15453 20855 15487
rect 21281 15453 21315 15487
rect 5365 15385 5399 15419
rect 7656 15385 7690 15419
rect 9220 15385 9254 15419
rect 10784 15385 10818 15419
rect 12725 15385 12759 15419
rect 18162 15385 18196 15419
rect 18705 15385 18739 15419
rect 19625 15385 19659 15419
rect 1501 15317 1535 15351
rect 2881 15317 2915 15351
rect 3433 15317 3467 15351
rect 3617 15317 3651 15351
rect 4169 15317 4203 15351
rect 4261 15317 4295 15351
rect 5917 15317 5951 15351
rect 6561 15317 6595 15351
rect 6929 15317 6963 15351
rect 7021 15317 7055 15351
rect 8769 15317 8803 15351
rect 10333 15317 10367 15351
rect 13093 15317 13127 15351
rect 13645 15317 13679 15351
rect 14289 15317 14323 15351
rect 14565 15317 14599 15351
rect 15301 15317 15335 15351
rect 16957 15317 16991 15351
rect 18797 15317 18831 15351
rect 20269 15317 20303 15351
rect 21005 15317 21039 15351
rect 21189 15317 21223 15351
rect 21465 15317 21499 15351
rect 2329 15113 2363 15147
rect 2421 15113 2455 15147
rect 4629 15113 4663 15147
rect 5089 15113 5123 15147
rect 5457 15113 5491 15147
rect 5917 15113 5951 15147
rect 6929 15113 6963 15147
rect 7389 15113 7423 15147
rect 8033 15113 8067 15147
rect 8493 15113 8527 15147
rect 8585 15113 8619 15147
rect 8953 15113 8987 15147
rect 9781 15113 9815 15147
rect 13001 15113 13035 15147
rect 13461 15113 13495 15147
rect 13921 15113 13955 15147
rect 14473 15113 14507 15147
rect 16957 15113 16991 15147
rect 19165 15113 19199 15147
rect 19901 15113 19935 15147
rect 3924 15045 3958 15079
rect 9413 15045 9447 15079
rect 11345 15045 11379 15079
rect 11897 15045 11931 15079
rect 17478 15045 17512 15079
rect 20085 15045 20119 15079
rect 20637 15045 20671 15079
rect 1685 14977 1719 15011
rect 2053 14977 2087 15011
rect 2145 14977 2179 15011
rect 2605 14977 2639 15011
rect 4169 14977 4203 15011
rect 4353 14977 4387 15011
rect 4997 14977 5031 15011
rect 5825 14977 5859 15011
rect 6745 14977 6779 15011
rect 7297 14977 7331 15011
rect 10241 14977 10275 15011
rect 10701 14977 10735 15011
rect 11989 14977 12023 15011
rect 13829 14977 13863 15011
rect 14289 14977 14323 15011
rect 15025 14977 15059 15011
rect 16037 14977 16071 15011
rect 17141 14977 17175 15011
rect 17233 14977 17267 15011
rect 19717 14977 19751 15011
rect 20913 14977 20947 15011
rect 21281 14977 21315 15011
rect 5273 14909 5307 14943
rect 6009 14909 6043 14943
rect 6653 14909 6687 14943
rect 7573 14909 7607 14943
rect 8401 14909 8435 14943
rect 9229 14909 9263 14943
rect 9321 14909 9355 14943
rect 10333 14909 10367 14943
rect 10425 14909 10459 14943
rect 12081 14909 12115 14943
rect 12725 14909 12759 14943
rect 12909 14909 12943 14943
rect 14013 14909 14047 14943
rect 15761 14909 15795 14943
rect 15945 14909 15979 14943
rect 20177 14909 20211 14943
rect 20821 14909 20855 14943
rect 1869 14841 1903 14875
rect 2789 14841 2823 14875
rect 4537 14841 4571 14875
rect 6469 14841 6503 14875
rect 11529 14841 11563 14875
rect 21097 14841 21131 14875
rect 1501 14773 1535 14807
rect 7849 14773 7883 14807
rect 9873 14773 9907 14807
rect 10977 14773 11011 14807
rect 12449 14773 12483 14807
rect 13369 14773 13403 14807
rect 15209 14773 15243 14807
rect 16405 14773 16439 14807
rect 18613 14773 18647 14807
rect 20453 14773 20487 14807
rect 21465 14773 21499 14807
rect 2145 14569 2179 14603
rect 2421 14569 2455 14603
rect 3525 14569 3559 14603
rect 4813 14569 4847 14603
rect 6285 14569 6319 14603
rect 7941 14569 7975 14603
rect 9965 14569 9999 14603
rect 16957 14569 16991 14603
rect 17785 14569 17819 14603
rect 19349 14569 19383 14603
rect 20729 14569 20763 14603
rect 21005 14569 21039 14603
rect 1869 14501 1903 14535
rect 2697 14501 2731 14535
rect 3801 14501 3835 14535
rect 9873 14501 9907 14535
rect 3249 14433 3283 14467
rect 4261 14433 4295 14467
rect 8493 14433 8527 14467
rect 9229 14433 9263 14467
rect 10609 14433 10643 14467
rect 13921 14433 13955 14467
rect 17141 14433 17175 14467
rect 17325 14433 17359 14467
rect 21097 14433 21131 14467
rect 1685 14365 1719 14399
rect 2053 14365 2087 14399
rect 2329 14365 2363 14399
rect 2605 14365 2639 14399
rect 2881 14365 2915 14399
rect 2973 14365 3007 14399
rect 4905 14365 4939 14399
rect 5172 14365 5206 14399
rect 7593 14365 7627 14399
rect 7849 14365 7883 14399
rect 8401 14365 8435 14399
rect 9045 14365 9079 14399
rect 9505 14365 9539 14399
rect 11906 14365 11940 14399
rect 12173 14365 12207 14399
rect 12265 14365 12299 14399
rect 14105 14365 14139 14399
rect 15577 14365 15611 14399
rect 20361 14365 20395 14399
rect 20545 14365 20579 14399
rect 20821 14365 20855 14399
rect 21281 14365 21315 14399
rect 3341 14297 3375 14331
rect 10425 14297 10459 14331
rect 12510 14297 12544 14331
rect 14350 14297 14384 14331
rect 15844 14297 15878 14331
rect 19441 14297 19475 14331
rect 19901 14297 19935 14331
rect 20269 14297 20303 14331
rect 1501 14229 1535 14263
rect 4353 14229 4387 14263
rect 4445 14229 4479 14263
rect 6469 14229 6503 14263
rect 8309 14229 8343 14263
rect 9413 14229 9447 14263
rect 10333 14229 10367 14263
rect 10793 14229 10827 14263
rect 13645 14229 13679 14263
rect 15485 14229 15519 14263
rect 17417 14229 17451 14263
rect 18889 14229 18923 14263
rect 19625 14229 19659 14263
rect 19993 14229 20027 14263
rect 21465 14229 21499 14263
rect 1869 14025 1903 14059
rect 2237 14025 2271 14059
rect 2605 14025 2639 14059
rect 3065 14025 3099 14059
rect 5641 14025 5675 14059
rect 6469 14025 6503 14059
rect 8493 14025 8527 14059
rect 8677 14025 8711 14059
rect 9413 14025 9447 14059
rect 9873 14025 9907 14059
rect 10333 14025 10367 14059
rect 11069 14025 11103 14059
rect 11253 14025 11287 14059
rect 12173 14025 12207 14059
rect 13369 14025 13403 14059
rect 13461 14025 13495 14059
rect 15669 14025 15703 14059
rect 16497 14025 16531 14059
rect 21005 14025 21039 14059
rect 4528 13957 4562 13991
rect 7358 13957 7392 13991
rect 11529 13957 11563 13991
rect 15209 13957 15243 13991
rect 1685 13889 1719 13923
rect 2053 13889 2087 13923
rect 2697 13889 2731 13923
rect 3433 13889 3467 13923
rect 3525 13889 3559 13923
rect 3985 13889 4019 13923
rect 4261 13889 4295 13923
rect 6009 13889 6043 13923
rect 6653 13889 6687 13923
rect 7113 13889 7147 13923
rect 9505 13889 9539 13923
rect 10241 13889 10275 13923
rect 12541 13889 12575 13923
rect 13001 13889 13035 13923
rect 13829 13889 13863 13923
rect 13921 13889 13955 13923
rect 14381 13889 14415 13923
rect 14841 13889 14875 13923
rect 15301 13889 15335 13923
rect 16129 13889 16163 13923
rect 17693 13889 17727 13923
rect 17960 13889 17994 13923
rect 19441 13889 19475 13923
rect 19533 13889 19567 13923
rect 20545 13889 20579 13923
rect 20821 13889 20855 13923
rect 21281 13889 21315 13923
rect 2789 13821 2823 13855
rect 3709 13821 3743 13855
rect 4169 13821 4203 13855
rect 5733 13821 5767 13855
rect 6745 13821 6779 13855
rect 6929 13821 6963 13855
rect 9689 13821 9723 13855
rect 10425 13821 10459 13855
rect 10885 13821 10919 13855
rect 11713 13821 11747 13855
rect 11897 13821 11931 13855
rect 12265 13821 12299 13855
rect 12817 13821 12851 13855
rect 12909 13821 12943 13855
rect 14105 13821 14139 13855
rect 15117 13821 15151 13855
rect 15853 13821 15887 13855
rect 16037 13821 16071 13855
rect 19257 13821 19291 13855
rect 20177 13821 20211 13855
rect 20361 13821 20395 13855
rect 21097 13821 21131 13855
rect 8953 13753 8987 13787
rect 20729 13753 20763 13787
rect 1501 13685 1535 13719
rect 9045 13685 9079 13719
rect 19073 13685 19107 13719
rect 19901 13685 19935 13719
rect 21465 13685 21499 13719
rect 4169 13481 4203 13515
rect 6929 13481 6963 13515
rect 11805 13481 11839 13515
rect 12449 13481 12483 13515
rect 15853 13481 15887 13515
rect 16221 13481 16255 13515
rect 18981 13481 19015 13515
rect 19257 13481 19291 13515
rect 20085 13481 20119 13515
rect 4997 13413 5031 13447
rect 8033 13413 8067 13447
rect 8953 13413 8987 13447
rect 11345 13413 11379 13447
rect 12541 13413 12575 13447
rect 13461 13413 13495 13447
rect 15761 13413 15795 13447
rect 4813 13345 4847 13379
rect 5549 13345 5583 13379
rect 7481 13345 7515 13379
rect 8585 13345 8619 13379
rect 10977 13345 11011 13379
rect 12081 13345 12115 13379
rect 12817 13345 12851 13379
rect 13001 13345 13035 13379
rect 16865 13345 16899 13379
rect 17601 13345 17635 13379
rect 19809 13345 19843 13379
rect 20637 13345 20671 13379
rect 1685 13277 1719 13311
rect 2053 13277 2087 13311
rect 3361 13277 3395 13311
rect 3617 13277 3651 13311
rect 5365 13277 5399 13311
rect 6745 13277 6779 13311
rect 8401 13277 8435 13311
rect 10333 13277 10367 13311
rect 10793 13277 10827 13311
rect 11713 13277 11747 13311
rect 13093 13277 13127 13311
rect 13645 13277 13679 13311
rect 14381 13277 14415 13311
rect 17325 13277 17359 13311
rect 17857 13277 17891 13311
rect 19625 13277 19659 13311
rect 20453 13277 20487 13311
rect 20913 13277 20947 13311
rect 21281 13277 21315 13311
rect 4629 13209 4663 13243
rect 5825 13209 5859 13243
rect 6009 13209 6043 13243
rect 6469 13209 6503 13243
rect 7297 13209 7331 13243
rect 8493 13209 8527 13243
rect 10066 13209 10100 13243
rect 14648 13209 14682 13243
rect 16589 13209 16623 13243
rect 20545 13209 20579 13243
rect 1501 13141 1535 13175
rect 1869 13141 1903 13175
rect 2237 13141 2271 13175
rect 3801 13141 3835 13175
rect 3985 13141 4019 13175
rect 4537 13141 4571 13175
rect 5457 13141 5491 13175
rect 6193 13141 6227 13175
rect 6561 13141 6595 13175
rect 7389 13141 7423 13175
rect 7849 13141 7883 13175
rect 10425 13141 10459 13175
rect 10885 13141 10919 13175
rect 11529 13141 11563 13175
rect 16037 13141 16071 13175
rect 16681 13141 16715 13175
rect 17233 13141 17267 13175
rect 17509 13141 17543 13175
rect 19717 13141 19751 13175
rect 21097 13141 21131 13175
rect 21465 13141 21499 13175
rect 2973 12937 3007 12971
rect 3249 12937 3283 12971
rect 3525 12937 3559 12971
rect 3893 12937 3927 12971
rect 7849 12937 7883 12971
rect 8309 12937 8343 12971
rect 9137 12937 9171 12971
rect 9505 12937 9539 12971
rect 9873 12937 9907 12971
rect 9965 12937 9999 12971
rect 10793 12937 10827 12971
rect 12909 12937 12943 12971
rect 13369 12937 13403 12971
rect 15209 12937 15243 12971
rect 18245 12937 18279 12971
rect 19809 12937 19843 12971
rect 20177 12937 20211 12971
rect 20269 12937 20303 12971
rect 20637 12937 20671 12971
rect 21005 12937 21039 12971
rect 2636 12869 2670 12903
rect 5273 12869 5307 12903
rect 8217 12869 8251 12903
rect 9045 12869 9079 12903
rect 14096 12869 14130 12903
rect 16405 12869 16439 12903
rect 18604 12869 18638 12903
rect 3157 12801 3191 12835
rect 3433 12801 3467 12835
rect 3985 12801 4019 12835
rect 5181 12801 5215 12835
rect 6101 12801 6135 12835
rect 6377 12801 6411 12835
rect 6644 12801 6678 12835
rect 10885 12801 10919 12835
rect 11345 12801 11379 12835
rect 11529 12801 11563 12835
rect 11796 12801 11830 12835
rect 13737 12801 13771 12835
rect 13829 12801 13863 12835
rect 15669 12801 15703 12835
rect 16865 12801 16899 12835
rect 17877 12801 17911 12835
rect 18337 12801 18371 12835
rect 20821 12801 20855 12835
rect 21281 12801 21315 12835
rect 2881 12733 2915 12767
rect 4077 12733 4111 12767
rect 4353 12733 4387 12767
rect 5457 12733 5491 12767
rect 8493 12733 8527 12767
rect 9229 12733 9263 12767
rect 10057 12733 10091 12767
rect 10333 12733 10367 12767
rect 10609 12733 10643 12767
rect 13001 12733 13035 12767
rect 15393 12733 15427 12767
rect 15577 12733 15611 12767
rect 17693 12733 17727 12767
rect 17785 12733 17819 12767
rect 20361 12733 20395 12767
rect 4813 12665 4847 12699
rect 5917 12665 5951 12699
rect 7757 12665 7791 12699
rect 13185 12665 13219 12699
rect 13553 12665 13587 12699
rect 16037 12665 16071 12699
rect 16313 12665 16347 12699
rect 19717 12665 19751 12699
rect 21189 12665 21223 12699
rect 1501 12597 1535 12631
rect 4629 12597 4663 12631
rect 5825 12597 5859 12631
rect 8677 12597 8711 12631
rect 11161 12597 11195 12631
rect 16773 12597 16807 12631
rect 17049 12597 17083 12631
rect 17417 12597 17451 12631
rect 21465 12597 21499 12631
rect 1501 12393 1535 12427
rect 3985 12393 4019 12427
rect 6285 12393 6319 12427
rect 8677 12393 8711 12427
rect 8953 12393 8987 12427
rect 9505 12393 9539 12427
rect 10609 12393 10643 12427
rect 13461 12393 13495 12427
rect 14105 12393 14139 12427
rect 15577 12393 15611 12427
rect 16405 12393 16439 12427
rect 18061 12393 18095 12427
rect 19441 12393 19475 12427
rect 20729 12393 20763 12427
rect 6193 12325 6227 12359
rect 8033 12325 8067 12359
rect 9321 12325 9355 12359
rect 10701 12325 10735 12359
rect 20913 12325 20947 12359
rect 3801 12257 3835 12291
rect 4537 12257 4571 12291
rect 6837 12257 6871 12291
rect 7113 12257 7147 12291
rect 7389 12257 7423 12291
rect 11069 12257 11103 12291
rect 13093 12257 13127 12291
rect 16129 12257 16163 12291
rect 16957 12257 16991 12291
rect 17417 12257 17451 12291
rect 18613 12257 18647 12291
rect 19717 12257 19751 12291
rect 1685 12189 1719 12223
rect 2053 12189 2087 12223
rect 2237 12189 2271 12223
rect 2504 12189 2538 12223
rect 4445 12189 4479 12223
rect 4813 12189 4847 12223
rect 7481 12189 7515 12223
rect 9137 12189 9171 12223
rect 12909 12189 12943 12223
rect 15485 12189 15519 12223
rect 17509 12189 17543 12223
rect 18889 12189 18923 12223
rect 19257 12189 19291 12223
rect 20545 12189 20579 12223
rect 21281 12189 21315 12223
rect 5080 12121 5114 12155
rect 6653 12121 6687 12155
rect 11336 12121 11370 12155
rect 15218 12121 15252 12155
rect 16773 12121 16807 12155
rect 17601 12121 17635 12155
rect 18521 12121 18555 12155
rect 19809 12121 19843 12155
rect 21097 12121 21131 12155
rect 1869 12053 1903 12087
rect 3617 12053 3651 12087
rect 4353 12053 4387 12087
rect 6745 12053 6779 12087
rect 7665 12053 7699 12087
rect 7941 12053 7975 12087
rect 8217 12053 8251 12087
rect 8493 12053 8527 12087
rect 9597 12053 9631 12087
rect 9873 12053 9907 12087
rect 10057 12053 10091 12087
rect 10241 12053 10275 12087
rect 10333 12053 10367 12087
rect 10885 12053 10919 12087
rect 12449 12053 12483 12087
rect 12541 12053 12575 12087
rect 13001 12053 13035 12087
rect 13553 12053 13587 12087
rect 13829 12053 13863 12087
rect 15945 12053 15979 12087
rect 16037 12053 16071 12087
rect 16865 12053 16899 12087
rect 17969 12053 18003 12087
rect 18429 12053 18463 12087
rect 19073 12053 19107 12087
rect 19901 12053 19935 12087
rect 20269 12053 20303 12087
rect 20361 12053 20395 12087
rect 21465 12053 21499 12087
rect 3249 11849 3283 11883
rect 3617 11849 3651 11883
rect 5365 11849 5399 11883
rect 5733 11849 5767 11883
rect 6469 11849 6503 11883
rect 7757 11849 7791 11883
rect 8125 11849 8159 11883
rect 8585 11849 8619 11883
rect 9045 11849 9079 11883
rect 11345 11849 11379 11883
rect 12173 11849 12207 11883
rect 13461 11849 13495 11883
rect 13921 11849 13955 11883
rect 15117 11849 15151 11883
rect 16681 11849 16715 11883
rect 17049 11849 17083 11883
rect 17877 11849 17911 11883
rect 18245 11849 18279 11883
rect 20361 11849 20395 11883
rect 20453 11849 20487 11883
rect 3709 11781 3743 11815
rect 4905 11781 4939 11815
rect 6837 11781 6871 11815
rect 7665 11781 7699 11815
rect 8493 11781 8527 11815
rect 9413 11781 9447 11815
rect 15669 11781 15703 11815
rect 1961 11713 1995 11747
rect 2697 11713 2731 11747
rect 4261 11713 4295 11747
rect 4537 11713 4571 11747
rect 4997 11713 5031 11747
rect 5825 11713 5859 11747
rect 9505 11713 9539 11747
rect 9965 11713 9999 11747
rect 10232 11713 10266 11747
rect 12265 11713 12299 11747
rect 13093 11713 13127 11747
rect 14749 11713 14783 11747
rect 15577 11713 15611 11747
rect 17141 11713 17175 11747
rect 18429 11713 18463 11747
rect 18889 11713 18923 11747
rect 18981 11713 19015 11747
rect 19237 11713 19271 11747
rect 20637 11713 20671 11747
rect 2237 11645 2271 11679
rect 2789 11645 2823 11679
rect 2973 11645 3007 11679
rect 3893 11645 3927 11679
rect 4813 11645 4847 11679
rect 5641 11645 5675 11679
rect 6929 11645 6963 11679
rect 7067 11645 7101 11679
rect 7941 11645 7975 11679
rect 8677 11645 8711 11679
rect 9229 11645 9263 11679
rect 12081 11645 12115 11679
rect 12817 11645 12851 11679
rect 13001 11645 13035 11679
rect 14013 11645 14047 11679
rect 14105 11645 14139 11679
rect 14473 11645 14507 11679
rect 14657 11645 14691 11679
rect 15853 11645 15887 11679
rect 16313 11645 16347 11679
rect 17233 11645 17267 11679
rect 17601 11645 17635 11679
rect 17785 11645 17819 11679
rect 21281 11645 21315 11679
rect 21557 11645 21591 11679
rect 4077 11577 4111 11611
rect 4353 11577 4387 11611
rect 6193 11577 6227 11611
rect 18705 11577 18739 11611
rect 2329 11509 2363 11543
rect 7297 11509 7331 11543
rect 9873 11509 9907 11543
rect 11529 11509 11563 11543
rect 11713 11509 11747 11543
rect 12633 11509 12667 11543
rect 13553 11509 13587 11543
rect 15209 11509 15243 11543
rect 16405 11509 16439 11543
rect 18613 11509 18647 11543
rect 3801 11305 3835 11339
rect 6745 11305 6779 11339
rect 7573 11305 7607 11339
rect 8769 11305 8803 11339
rect 11253 11305 11287 11339
rect 11529 11305 11563 11339
rect 12357 11305 12391 11339
rect 13185 11305 13219 11339
rect 13369 11305 13403 11339
rect 13829 11305 13863 11339
rect 14565 11305 14599 11339
rect 14749 11305 14783 11339
rect 15577 11305 15611 11339
rect 16405 11305 16439 11339
rect 17233 11305 17267 11339
rect 17417 11305 17451 11339
rect 1685 11237 1719 11271
rect 3617 11237 3651 11271
rect 5917 11237 5951 11271
rect 6653 11237 6687 11271
rect 10885 11237 10919 11271
rect 14381 11237 14415 11271
rect 19073 11237 19107 11271
rect 4445 11169 4479 11203
rect 4537 11169 4571 11203
rect 6101 11169 6135 11203
rect 6377 11169 6411 11203
rect 7389 11169 7423 11203
rect 8217 11169 8251 11203
rect 9137 11169 9171 11203
rect 11805 11169 11839 11203
rect 12541 11169 12575 11203
rect 15209 11169 15243 11203
rect 15301 11169 15335 11203
rect 16129 11169 16163 11203
rect 16957 11169 16991 11203
rect 17693 11169 17727 11203
rect 20637 11169 20671 11203
rect 21281 11169 21315 11203
rect 1501 11101 1535 11135
rect 2237 11101 2271 11135
rect 2504 11101 2538 11135
rect 3985 11101 4019 11135
rect 7941 11101 7975 11135
rect 8309 11101 8343 11135
rect 8401 11101 8435 11135
rect 8953 11101 8987 11135
rect 11989 11101 12023 11135
rect 12817 11101 12851 11135
rect 16773 11101 16807 11135
rect 16865 11101 16899 11135
rect 20370 11101 20404 11135
rect 21189 11101 21223 11135
rect 1869 11033 1903 11067
rect 2053 11033 2087 11067
rect 4169 11033 4203 11067
rect 4804 11033 4838 11067
rect 9382 11033 9416 11067
rect 13645 11033 13679 11067
rect 14289 11033 14323 11067
rect 15117 11033 15151 11067
rect 17960 11033 17994 11067
rect 21097 11033 21131 11067
rect 7113 10965 7147 10999
rect 7205 10965 7239 10999
rect 10517 10965 10551 10999
rect 10609 10965 10643 10999
rect 11161 10965 11195 10999
rect 11897 10965 11931 10999
rect 12725 10965 12759 10999
rect 15945 10965 15979 10999
rect 16037 10965 16071 10999
rect 19257 10965 19291 10999
rect 20729 10965 20763 10999
rect 1593 10761 1627 10795
rect 3433 10761 3467 10795
rect 5641 10761 5675 10795
rect 6745 10761 6779 10795
rect 7021 10761 7055 10795
rect 8309 10761 8343 10795
rect 9781 10761 9815 10795
rect 10149 10761 10183 10795
rect 11805 10761 11839 10795
rect 14197 10761 14231 10795
rect 14381 10761 14415 10795
rect 16129 10761 16163 10795
rect 16681 10761 16715 10795
rect 18061 10761 18095 10795
rect 18521 10761 18555 10795
rect 20177 10761 20211 10795
rect 20269 10761 20303 10795
rect 4528 10693 4562 10727
rect 6929 10693 6963 10727
rect 7389 10693 7423 10727
rect 7481 10693 7515 10727
rect 9422 10693 9456 10727
rect 12602 10693 12636 10727
rect 15016 10693 15050 10727
rect 20637 10693 20671 10727
rect 21281 10693 21315 10727
rect 2706 10625 2740 10659
rect 3249 10625 3283 10659
rect 3801 10625 3835 10659
rect 5733 10625 5767 10659
rect 6009 10625 6043 10659
rect 7941 10625 7975 10659
rect 8217 10625 8251 10659
rect 11345 10625 11379 10659
rect 11897 10625 11931 10659
rect 12357 10625 12391 10659
rect 14749 10625 14783 10659
rect 17049 10625 17083 10659
rect 17509 10625 17543 10659
rect 18153 10625 18187 10659
rect 18981 10625 19015 10659
rect 19809 10625 19843 10659
rect 21097 10625 21131 10659
rect 21465 10625 21499 10659
rect 2973 10557 3007 10591
rect 3893 10557 3927 10591
rect 3985 10557 4019 10591
rect 4261 10557 4295 10591
rect 6377 10557 6411 10591
rect 7573 10557 7607 10591
rect 9689 10557 9723 10591
rect 10241 10557 10275 10591
rect 10425 10557 10459 10591
rect 11621 10557 11655 10591
rect 13921 10557 13955 10591
rect 16221 10557 16255 10591
rect 17141 10557 17175 10591
rect 17325 10557 17359 10591
rect 17969 10557 18003 10591
rect 19073 10557 19107 10591
rect 19165 10557 19199 10591
rect 19625 10557 19659 10591
rect 19717 10557 19751 10591
rect 20729 10557 20763 10591
rect 20821 10557 20855 10591
rect 8033 10489 8067 10523
rect 10793 10489 10827 10523
rect 14013 10489 14047 10523
rect 18613 10489 18647 10523
rect 1501 10421 1535 10455
rect 3065 10421 3099 10455
rect 6101 10421 6135 10455
rect 10609 10421 10643 10455
rect 11069 10421 11103 10455
rect 12265 10421 12299 10455
rect 13737 10421 13771 10455
rect 14657 10421 14691 10455
rect 16405 10421 16439 10455
rect 4721 10217 4755 10251
rect 5825 10217 5859 10251
rect 10425 10217 10459 10251
rect 13553 10217 13587 10251
rect 15669 10217 15703 10251
rect 16221 10217 16255 10251
rect 18705 10217 18739 10251
rect 20269 10217 20303 10251
rect 6653 10149 6687 10183
rect 7113 10149 7147 10183
rect 13829 10149 13863 10183
rect 14841 10149 14875 10183
rect 20637 10149 20671 10183
rect 1685 10081 1719 10115
rect 3249 10081 3283 10115
rect 3617 10081 3651 10115
rect 5273 10081 5307 10115
rect 6285 10081 6319 10115
rect 6469 10081 6503 10115
rect 7389 10081 7423 10115
rect 8217 10081 8251 10115
rect 9597 10081 9631 10115
rect 11253 10081 11287 10115
rect 11989 10081 12023 10115
rect 12081 10081 12115 10115
rect 13001 10081 13035 10115
rect 14197 10081 14231 10115
rect 14381 10081 14415 10115
rect 15025 10081 15059 10115
rect 16589 10081 16623 10115
rect 17325 10081 17359 10115
rect 19625 10081 19659 10115
rect 21005 10081 21039 10115
rect 3801 10013 3835 10047
rect 4077 10013 4111 10047
rect 5089 10013 5123 10047
rect 6837 10013 6871 10047
rect 7573 10013 7607 10047
rect 8953 10013 8987 10047
rect 12633 10013 12667 10047
rect 13185 10013 13219 10047
rect 14473 10013 14507 10047
rect 15301 10013 15335 10047
rect 15761 10013 15795 10047
rect 16773 10013 16807 10047
rect 19901 10013 19935 10047
rect 20729 10013 20763 10047
rect 1501 9945 1535 9979
rect 2982 9945 3016 9979
rect 3433 9945 3467 9979
rect 9689 9945 9723 9979
rect 10241 9945 10275 9979
rect 11529 9945 11563 9979
rect 13093 9945 13127 9979
rect 16037 9945 16071 9979
rect 17570 9945 17604 9979
rect 18797 9945 18831 9979
rect 18981 9945 19015 9979
rect 19441 9945 19475 9979
rect 20453 9945 20487 9979
rect 1869 9877 1903 9911
rect 5181 9877 5215 9911
rect 5641 9877 5675 9911
rect 6193 9877 6227 9911
rect 7481 9877 7515 9911
rect 7941 9877 7975 9911
rect 8309 9877 8343 9911
rect 8401 9877 8435 9911
rect 8769 9877 8803 9911
rect 9137 9877 9171 9911
rect 9321 9877 9355 9911
rect 9781 9877 9815 9911
rect 10149 9877 10183 9911
rect 10701 9877 10735 9911
rect 11069 9877 11103 9911
rect 11161 9877 11195 9911
rect 12173 9877 12207 9911
rect 12541 9877 12575 9911
rect 13645 9877 13679 9911
rect 15209 9877 15243 9911
rect 15945 9877 15979 9911
rect 16865 9877 16899 9911
rect 17233 9877 17267 9911
rect 19809 9877 19843 9911
rect 1593 9673 1627 9707
rect 4629 9673 4663 9707
rect 7573 9673 7607 9707
rect 9597 9673 9631 9707
rect 10517 9673 10551 9707
rect 10885 9673 10919 9707
rect 11345 9673 11379 9707
rect 11989 9673 12023 9707
rect 13277 9673 13311 9707
rect 19533 9673 19567 9707
rect 20361 9673 20395 9707
rect 3810 9605 3844 9639
rect 6745 9605 6779 9639
rect 12081 9605 12115 9639
rect 13728 9605 13762 9639
rect 17570 9605 17604 9639
rect 19993 9605 20027 9639
rect 21465 9605 21499 9639
rect 1409 9537 1443 9571
rect 2053 9537 2087 9571
rect 4169 9537 4203 9571
rect 4997 9537 5031 9571
rect 5089 9537 5123 9571
rect 5825 9537 5859 9571
rect 6837 9537 6871 9571
rect 7665 9537 7699 9571
rect 8125 9537 8159 9571
rect 8381 9537 8415 9571
rect 9965 9537 9999 9571
rect 10977 9537 11011 9571
rect 12909 9537 12943 9571
rect 15301 9537 15335 9571
rect 16129 9537 16163 9571
rect 17233 9537 17267 9571
rect 17325 9537 17359 9571
rect 18797 9537 18831 9571
rect 18981 9537 19015 9571
rect 19441 9537 19475 9571
rect 19901 9537 19935 9571
rect 20729 9537 20763 9571
rect 1869 9469 1903 9503
rect 1961 9469 1995 9503
rect 4077 9469 4111 9503
rect 4445 9469 4479 9503
rect 5181 9469 5215 9503
rect 5917 9469 5951 9503
rect 6101 9469 6135 9503
rect 7021 9469 7055 9503
rect 7481 9469 7515 9503
rect 10057 9469 10091 9503
rect 10149 9469 10183 9503
rect 10701 9469 10735 9503
rect 11805 9469 11839 9503
rect 12633 9469 12667 9503
rect 12817 9469 12851 9503
rect 13461 9469 13495 9503
rect 15117 9469 15151 9503
rect 15209 9469 15243 9503
rect 15945 9469 15979 9503
rect 16037 9469 16071 9503
rect 20085 9469 20119 9503
rect 20821 9469 20855 9503
rect 20913 9469 20947 9503
rect 2421 9401 2455 9435
rect 2697 9401 2731 9435
rect 5457 9401 5491 9435
rect 6377 9401 6411 9435
rect 12449 9401 12483 9435
rect 16497 9401 16531 9435
rect 18705 9401 18739 9435
rect 21281 9401 21315 9435
rect 2605 9333 2639 9367
rect 4353 9333 4387 9367
rect 8033 9333 8067 9367
rect 9505 9333 9539 9367
rect 11529 9333 11563 9367
rect 14841 9333 14875 9367
rect 15669 9333 15703 9367
rect 16681 9333 16715 9367
rect 16865 9333 16899 9367
rect 17049 9333 17083 9367
rect 19257 9333 19291 9367
rect 2145 9129 2179 9163
rect 3249 9129 3283 9163
rect 4077 9129 4111 9163
rect 7389 9129 7423 9163
rect 8953 9129 8987 9163
rect 9137 9129 9171 9163
rect 9413 9129 9447 9163
rect 10241 9129 10275 9163
rect 13093 9129 13127 9163
rect 13185 9129 13219 9163
rect 14565 9129 14599 9163
rect 16221 9129 16255 9163
rect 17785 9129 17819 9163
rect 19073 9129 19107 9163
rect 20729 9129 20763 9163
rect 3617 9061 3651 9095
rect 10333 9061 10367 9095
rect 18613 9061 18647 9095
rect 1593 8993 1627 9027
rect 2881 8993 2915 9027
rect 4629 8993 4663 9027
rect 5457 8993 5491 9027
rect 6285 8993 6319 9027
rect 7113 8993 7147 9027
rect 9689 8993 9723 9027
rect 11805 8993 11839 9027
rect 12449 8993 12483 9027
rect 12633 8993 12667 9027
rect 13645 8993 13679 9027
rect 14841 8993 14875 9027
rect 18245 8993 18279 9027
rect 18429 8993 18463 9027
rect 21281 8993 21315 9027
rect 2605 8925 2639 8959
rect 3065 8925 3099 8959
rect 3433 8925 3467 8959
rect 4445 8925 4479 8959
rect 5273 8925 5307 8959
rect 6101 8925 6135 8959
rect 6929 8925 6963 8959
rect 8769 8925 8803 8959
rect 9781 8925 9815 8959
rect 11446 8925 11480 8959
rect 11713 8925 11747 8959
rect 13461 8925 13495 8959
rect 13829 8925 13863 8959
rect 14381 8925 14415 8959
rect 16313 8925 16347 8959
rect 16569 8925 16603 8959
rect 18889 8925 18923 8959
rect 19257 8925 19291 8959
rect 19524 8925 19558 8959
rect 1685 8857 1719 8891
rect 4537 8857 4571 8891
rect 8513 8857 8547 8891
rect 9873 8857 9907 8891
rect 12173 8857 12207 8891
rect 15108 8857 15142 8891
rect 1777 8789 1811 8823
rect 2237 8789 2271 8823
rect 2697 8789 2731 8823
rect 3801 8789 3835 8823
rect 4905 8789 4939 8823
rect 5365 8789 5399 8823
rect 5733 8789 5767 8823
rect 6193 8789 6227 8823
rect 6561 8789 6595 8823
rect 7021 8789 7055 8823
rect 12725 8789 12759 8823
rect 14197 8789 14231 8823
rect 17693 8789 17727 8823
rect 18153 8789 18187 8823
rect 20637 8789 20671 8823
rect 21097 8789 21131 8823
rect 21189 8789 21223 8823
rect 1593 8585 1627 8619
rect 2329 8585 2363 8619
rect 3433 8585 3467 8619
rect 3893 8585 3927 8619
rect 3985 8585 4019 8619
rect 4353 8585 4387 8619
rect 4721 8585 4755 8619
rect 5181 8585 5215 8619
rect 5549 8585 5583 8619
rect 6377 8585 6411 8619
rect 7941 8585 7975 8619
rect 8769 8585 8803 8619
rect 9137 8585 9171 8619
rect 9597 8585 9631 8619
rect 11621 8585 11655 8619
rect 12725 8585 12759 8619
rect 13277 8585 13311 8619
rect 14565 8585 14599 8619
rect 14933 8585 14967 8619
rect 16037 8585 16071 8619
rect 16497 8585 16531 8619
rect 16957 8585 16991 8619
rect 17049 8585 17083 8619
rect 17417 8585 17451 8619
rect 17693 8585 17727 8619
rect 19441 8585 19475 8619
rect 20085 8585 20119 8619
rect 20453 8585 20487 8619
rect 21005 8585 21039 8619
rect 5641 8517 5675 8551
rect 8309 8517 8343 8551
rect 9229 8517 9263 8551
rect 10710 8517 10744 8551
rect 11161 8517 11195 8551
rect 14473 8517 14507 8551
rect 15393 8517 15427 8551
rect 15669 8517 15703 8551
rect 18990 8517 19024 8551
rect 21097 8517 21131 8551
rect 1409 8449 1443 8483
rect 2237 8449 2271 8483
rect 3065 8449 3099 8483
rect 4813 8449 4847 8483
rect 6193 8449 6227 8483
rect 7490 8449 7524 8483
rect 11253 8449 11287 8483
rect 12173 8449 12207 8483
rect 12909 8449 12943 8483
rect 13645 8449 13679 8483
rect 14105 8449 14139 8483
rect 16129 8449 16163 8483
rect 19257 8449 19291 8483
rect 19533 8449 19567 8483
rect 19901 8449 19935 8483
rect 21465 8449 21499 8483
rect 2421 8381 2455 8415
rect 2789 8381 2823 8415
rect 2973 8381 3007 8415
rect 4077 8381 4111 8415
rect 4905 8381 4939 8415
rect 5733 8381 5767 8415
rect 7757 8381 7791 8415
rect 8401 8381 8435 8415
rect 8585 8381 8619 8415
rect 9321 8381 9355 8415
rect 10977 8381 11011 8415
rect 12265 8381 12299 8415
rect 12357 8381 12391 8415
rect 13553 8381 13587 8415
rect 14289 8381 14323 8415
rect 15025 8381 15059 8415
rect 15945 8381 15979 8415
rect 16865 8381 16899 8415
rect 19717 8381 19751 8415
rect 20545 8381 20579 8415
rect 20637 8381 20671 8415
rect 3525 8313 3559 8347
rect 13093 8313 13127 8347
rect 13829 8313 13863 8347
rect 17877 8313 17911 8347
rect 1869 8245 1903 8279
rect 6009 8245 6043 8279
rect 11805 8245 11839 8279
rect 13921 8245 13955 8279
rect 21373 8245 21407 8279
rect 2421 8041 2455 8075
rect 2881 8041 2915 8075
rect 5273 8041 5307 8075
rect 6101 8041 6135 8075
rect 7205 8041 7239 8075
rect 11437 8041 11471 8075
rect 16313 8041 16347 8075
rect 16589 8041 16623 8075
rect 19257 8041 19291 8075
rect 20177 8041 20211 8075
rect 21373 8041 21407 8075
rect 21465 8041 21499 8075
rect 2789 7973 2823 8007
rect 6929 7973 6963 8007
rect 8769 7973 8803 8007
rect 10517 7973 10551 8007
rect 13921 7973 13955 8007
rect 16773 7973 16807 8007
rect 17601 7973 17635 8007
rect 19073 7973 19107 8007
rect 20269 7973 20303 8007
rect 1777 7905 1811 7939
rect 1961 7905 1995 7939
rect 3525 7905 3559 7939
rect 5825 7905 5859 7939
rect 6653 7905 6687 7939
rect 8125 7905 8159 7939
rect 9505 7905 9539 7939
rect 9873 7905 9907 7939
rect 11161 7905 11195 7939
rect 12817 7905 12851 7939
rect 13461 7905 13495 7939
rect 14749 7905 14783 7939
rect 15577 7905 15611 7939
rect 17049 7905 17083 7939
rect 17693 7905 17727 7939
rect 19809 7905 19843 7939
rect 20729 7905 20763 7939
rect 1409 7837 1443 7871
rect 2605 7837 2639 7871
rect 4914 7837 4948 7871
rect 5181 7837 5215 7871
rect 7113 7837 7147 7871
rect 7849 7837 7883 7871
rect 8309 7837 8343 7871
rect 8401 7837 8435 7871
rect 9321 7837 9355 7871
rect 10149 7837 10183 7871
rect 11069 7837 11103 7871
rect 13277 7837 13311 7871
rect 13737 7837 13771 7871
rect 14565 7837 14599 7871
rect 15485 7837 15519 7871
rect 17233 7837 17267 7871
rect 20453 7837 20487 7871
rect 3249 7769 3283 7803
rect 6469 7769 6503 7803
rect 10057 7769 10091 7803
rect 12572 7769 12606 7803
rect 15853 7769 15887 7803
rect 16221 7769 16255 7803
rect 17960 7769 17994 7803
rect 20913 7769 20947 7803
rect 1593 7701 1627 7735
rect 2053 7701 2087 7735
rect 3341 7701 3375 7735
rect 3801 7701 3835 7735
rect 5641 7701 5675 7735
rect 5733 7701 5767 7735
rect 6561 7701 6595 7735
rect 7573 7701 7607 7735
rect 7757 7701 7791 7735
rect 8953 7701 8987 7735
rect 9413 7701 9447 7735
rect 10609 7701 10643 7735
rect 10977 7701 11011 7735
rect 12909 7701 12943 7735
rect 13369 7701 13403 7735
rect 14197 7701 14231 7735
rect 14657 7701 14691 7735
rect 15025 7701 15059 7735
rect 15393 7701 15427 7735
rect 17141 7701 17175 7735
rect 19625 7701 19659 7735
rect 19717 7701 19751 7735
rect 21005 7701 21039 7735
rect 1961 7497 1995 7531
rect 2421 7497 2455 7531
rect 2789 7497 2823 7531
rect 4261 7497 4295 7531
rect 4721 7497 4755 7531
rect 6193 7497 6227 7531
rect 7113 7497 7147 7531
rect 7573 7497 7607 7531
rect 9965 7497 9999 7531
rect 10333 7497 10367 7531
rect 11345 7497 11379 7531
rect 11897 7497 11931 7531
rect 12173 7497 12207 7531
rect 12633 7497 12667 7531
rect 15301 7497 15335 7531
rect 16313 7497 16347 7531
rect 19349 7497 19383 7531
rect 19441 7497 19475 7531
rect 20361 7497 20395 7531
rect 20453 7497 20487 7531
rect 1501 7429 1535 7463
rect 2329 7429 2363 7463
rect 8289 7429 8323 7463
rect 10885 7429 10919 7463
rect 10977 7429 11011 7463
rect 11621 7429 11655 7463
rect 16129 7429 16163 7463
rect 17049 7429 17083 7463
rect 20913 7429 20947 7463
rect 3902 7361 3936 7395
rect 4169 7361 4203 7395
rect 4445 7361 4479 7395
rect 4537 7361 4571 7395
rect 5069 7361 5103 7395
rect 6377 7361 6411 7395
rect 6653 7361 6687 7395
rect 6929 7361 6963 7395
rect 7665 7361 7699 7395
rect 8033 7361 8067 7395
rect 9873 7361 9907 7395
rect 12541 7361 12575 7395
rect 13820 7361 13854 7395
rect 15393 7361 15427 7395
rect 17141 7361 17175 7395
rect 17408 7361 17442 7395
rect 18981 7361 19015 7395
rect 19809 7361 19843 7395
rect 20821 7361 20855 7395
rect 21465 7361 21499 7395
rect 2513 7293 2547 7327
rect 4813 7293 4847 7327
rect 7849 7293 7883 7327
rect 10057 7293 10091 7327
rect 10701 7293 10735 7327
rect 12725 7293 12759 7327
rect 13001 7293 13035 7327
rect 13553 7293 13587 7327
rect 15117 7293 15151 7327
rect 16405 7293 16439 7327
rect 18705 7293 18739 7327
rect 18889 7293 18923 7327
rect 19901 7293 19935 7327
rect 19993 7293 20027 7327
rect 21005 7293 21039 7327
rect 1685 7225 1719 7259
rect 9505 7225 9539 7259
rect 15945 7225 15979 7259
rect 18521 7225 18555 7259
rect 21281 7225 21315 7259
rect 1777 7157 1811 7191
rect 6561 7157 6595 7191
rect 6837 7157 6871 7191
rect 7205 7157 7239 7191
rect 9413 7157 9447 7191
rect 11713 7157 11747 7191
rect 13185 7157 13219 7191
rect 13369 7157 13403 7191
rect 14933 7157 14967 7191
rect 15761 7157 15795 7191
rect 16681 7157 16715 7191
rect 2421 6953 2455 6987
rect 11805 6953 11839 6987
rect 15669 6953 15703 6987
rect 18981 6953 19015 6987
rect 3249 6885 3283 6919
rect 3617 6885 3651 6919
rect 5365 6885 5399 6919
rect 1869 6817 1903 6851
rect 2697 6817 2731 6851
rect 4905 6817 4939 6851
rect 6101 6817 6135 6851
rect 6929 6817 6963 6851
rect 10885 6817 10919 6851
rect 11529 6817 11563 6851
rect 12357 6817 12391 6851
rect 12725 6817 12759 6851
rect 13553 6817 13587 6851
rect 14197 6817 14231 6851
rect 15025 6817 15059 6851
rect 15209 6817 15243 6851
rect 18061 6817 18095 6851
rect 18429 6817 18463 6851
rect 21005 6817 21039 6851
rect 1409 6749 1443 6783
rect 1961 6749 1995 6783
rect 2881 6749 2915 6783
rect 3801 6749 3835 6783
rect 4077 6749 4111 6783
rect 4721 6749 4755 6783
rect 5181 6749 5215 6783
rect 8585 6749 8619 6783
rect 8953 6749 8987 6783
rect 9413 6749 9447 6783
rect 12173 6749 12207 6783
rect 12265 6749 12299 6783
rect 13737 6749 13771 6783
rect 14473 6749 14507 6783
rect 15853 6749 15887 6783
rect 17058 6749 17092 6783
rect 17325 6749 17359 6783
rect 18521 6749 18555 6783
rect 18613 6749 18647 6783
rect 19257 6749 19291 6783
rect 19524 6749 19558 6783
rect 20729 6749 20763 6783
rect 2053 6681 2087 6715
rect 3433 6681 3467 6715
rect 6837 6681 6871 6715
rect 8340 6681 8374 6715
rect 10618 6681 10652 6715
rect 13001 6681 13035 6715
rect 14381 6681 14415 6715
rect 15301 6681 15335 6715
rect 1593 6613 1627 6647
rect 2789 6613 2823 6647
rect 4261 6613 4295 6647
rect 4353 6613 4387 6647
rect 4813 6613 4847 6647
rect 5549 6613 5583 6647
rect 5917 6613 5951 6647
rect 6009 6613 6043 6647
rect 6377 6613 6411 6647
rect 6745 6613 6779 6647
rect 7205 6613 7239 6647
rect 8769 6613 8803 6647
rect 9137 6613 9171 6647
rect 9229 6613 9263 6647
rect 9505 6613 9539 6647
rect 10977 6613 11011 6647
rect 11345 6613 11379 6647
rect 11437 6613 11471 6647
rect 12909 6613 12943 6647
rect 13369 6613 13403 6647
rect 13829 6613 13863 6647
rect 14841 6613 14875 6647
rect 15945 6613 15979 6647
rect 17417 6613 17451 6647
rect 17785 6613 17819 6647
rect 17877 6613 17911 6647
rect 20637 6613 20671 6647
rect 1593 6409 1627 6443
rect 6009 6409 6043 6443
rect 6745 6409 6779 6443
rect 6837 6409 6871 6443
rect 7205 6409 7239 6443
rect 7665 6409 7699 6443
rect 8401 6409 8435 6443
rect 8493 6409 8527 6443
rect 9321 6409 9355 6443
rect 9781 6409 9815 6443
rect 10241 6409 10275 6443
rect 10609 6409 10643 6443
rect 10977 6409 11011 6443
rect 11069 6409 11103 6443
rect 11529 6409 11563 6443
rect 11989 6409 12023 6443
rect 13277 6409 13311 6443
rect 13553 6409 13587 6443
rect 15577 6409 15611 6443
rect 16957 6409 16991 6443
rect 17049 6409 17083 6443
rect 17509 6409 17543 6443
rect 18705 6409 18739 6443
rect 18981 6409 19015 6443
rect 19349 6409 19383 6443
rect 19809 6409 19843 6443
rect 20269 6409 20303 6443
rect 21005 6409 21039 6443
rect 21373 6409 21407 6443
rect 2706 6341 2740 6375
rect 3608 6341 3642 6375
rect 7573 6341 7607 6375
rect 10149 6341 10183 6375
rect 14096 6341 14130 6375
rect 15669 6341 15703 6375
rect 20177 6341 20211 6375
rect 3065 6273 3099 6307
rect 3341 6273 3375 6307
rect 5733 6273 5767 6307
rect 6193 6273 6227 6307
rect 11897 6273 11931 6307
rect 12357 6273 12391 6307
rect 16221 6273 16255 6307
rect 17877 6273 17911 6307
rect 18529 6273 18563 6307
rect 18797 6273 18831 6307
rect 2973 6205 3007 6239
rect 4813 6205 4847 6239
rect 5089 6205 5123 6239
rect 7021 6205 7055 6239
rect 7757 6205 7791 6239
rect 8585 6205 8619 6239
rect 9045 6205 9079 6239
rect 9229 6205 9263 6239
rect 10425 6205 10459 6239
rect 11161 6205 11195 6239
rect 12081 6205 12115 6239
rect 13829 6205 13863 6239
rect 15393 6205 15427 6239
rect 16497 6205 16531 6239
rect 16865 6205 16899 6239
rect 17969 6205 18003 6239
rect 18153 6205 18187 6239
rect 19441 6205 19475 6239
rect 19625 6205 19659 6239
rect 20361 6205 20395 6239
rect 20729 6205 20763 6239
rect 20913 6205 20947 6239
rect 21465 6205 21499 6239
rect 12817 6137 12851 6171
rect 15209 6137 15243 6171
rect 1501 6069 1535 6103
rect 4721 6069 4755 6103
rect 5917 6069 5951 6103
rect 6377 6069 6411 6103
rect 8033 6069 8067 6103
rect 9689 6069 9723 6103
rect 12725 6069 12759 6103
rect 13093 6069 13127 6103
rect 13369 6069 13403 6103
rect 16037 6069 16071 6103
rect 17417 6069 17451 6103
rect 18337 6069 18371 6103
rect 1961 5865 1995 5899
rect 3617 5865 3651 5899
rect 5825 5865 5859 5899
rect 6377 5865 6411 5899
rect 10333 5865 10367 5899
rect 10793 5865 10827 5899
rect 11161 5865 11195 5899
rect 16497 5865 16531 5899
rect 18705 5865 18739 5899
rect 20637 5865 20671 5899
rect 7205 5797 7239 5831
rect 13829 5797 13863 5831
rect 15577 5797 15611 5831
rect 2145 5729 2179 5763
rect 3065 5729 3099 5763
rect 4445 5729 4479 5763
rect 6929 5729 6963 5763
rect 7757 5729 7791 5763
rect 8677 5729 8711 5763
rect 8953 5729 8987 5763
rect 11713 5729 11747 5763
rect 13093 5729 13127 5763
rect 13277 5729 13311 5763
rect 15945 5729 15979 5763
rect 16037 5729 16071 5763
rect 17049 5729 17083 5763
rect 17233 5729 17267 5763
rect 17877 5729 17911 5763
rect 21281 5729 21315 5763
rect 1777 5661 1811 5695
rect 3249 5661 3283 5695
rect 3801 5661 3835 5695
rect 4169 5661 4203 5695
rect 4712 5661 4746 5695
rect 5917 5661 5951 5695
rect 6837 5661 6871 5695
rect 8493 5661 8527 5695
rect 9209 5661 9243 5695
rect 10609 5661 10643 5695
rect 11621 5661 11655 5695
rect 12173 5661 12207 5695
rect 13001 5661 13035 5695
rect 13645 5661 13679 5695
rect 15218 5661 15252 5695
rect 15485 5661 15519 5695
rect 17417 5661 17451 5695
rect 19257 5661 19291 5695
rect 21189 5661 21223 5695
rect 1501 5593 1535 5627
rect 1685 5593 1719 5627
rect 2329 5593 2363 5627
rect 7573 5593 7607 5627
rect 8401 5593 8435 5627
rect 11989 5593 12023 5627
rect 17601 5593 17635 5627
rect 18797 5593 18831 5627
rect 18981 5593 19015 5627
rect 19524 5593 19558 5627
rect 2421 5525 2455 5559
rect 2789 5525 2823 5559
rect 3157 5525 3191 5559
rect 3985 5525 4019 5559
rect 4353 5525 4387 5559
rect 6101 5525 6135 5559
rect 6285 5525 6319 5559
rect 6745 5525 6779 5559
rect 7665 5525 7699 5559
rect 8033 5525 8067 5559
rect 10425 5525 10459 5559
rect 11069 5525 11103 5559
rect 11529 5525 11563 5559
rect 12357 5525 12391 5559
rect 12633 5525 12667 5559
rect 13461 5525 13495 5559
rect 14105 5525 14139 5559
rect 16129 5525 16163 5559
rect 16589 5525 16623 5559
rect 16957 5525 16991 5559
rect 18061 5525 18095 5559
rect 18153 5525 18187 5559
rect 18521 5525 18555 5559
rect 20729 5525 20763 5559
rect 21097 5525 21131 5559
rect 4353 5321 4387 5355
rect 4721 5321 4755 5355
rect 5457 5321 5491 5355
rect 7205 5321 7239 5355
rect 7573 5321 7607 5355
rect 8217 5321 8251 5355
rect 8309 5321 8343 5355
rect 8677 5321 8711 5355
rect 10149 5321 10183 5355
rect 11345 5321 11379 5355
rect 12081 5321 12115 5355
rect 12449 5321 12483 5355
rect 14565 5321 14599 5355
rect 14749 5321 14783 5355
rect 15025 5321 15059 5355
rect 15209 5321 15243 5355
rect 16037 5321 16071 5355
rect 16681 5321 16715 5355
rect 20177 5321 20211 5355
rect 2697 5253 2731 5287
rect 5917 5253 5951 5287
rect 15485 5253 15519 5287
rect 16129 5253 16163 5287
rect 17049 5253 17083 5287
rect 20269 5253 20303 5287
rect 1961 5185 1995 5219
rect 2421 5185 2455 5219
rect 3137 5185 3171 5219
rect 5181 5185 5215 5219
rect 5825 5185 5859 5219
rect 6745 5185 6779 5219
rect 7389 5185 7423 5219
rect 7849 5185 7883 5219
rect 8769 5185 8803 5219
rect 9036 5185 9070 5219
rect 10241 5185 10275 5219
rect 10977 5185 11011 5219
rect 11713 5185 11747 5219
rect 12541 5185 12575 5219
rect 14114 5185 14148 5219
rect 14381 5185 14415 5219
rect 15669 5185 15703 5219
rect 17877 5185 17911 5219
rect 18593 5185 18627 5219
rect 21557 5185 21591 5219
rect 2237 5117 2271 5151
rect 2881 5117 2915 5151
rect 4813 5117 4847 5151
rect 4905 5117 4939 5151
rect 6009 5117 6043 5151
rect 6837 5117 6871 5151
rect 6929 5117 6963 5151
rect 8125 5117 8159 5151
rect 10793 5117 10827 5151
rect 10885 5117 10919 5151
rect 12357 5117 12391 5151
rect 15945 5117 15979 5151
rect 17141 5117 17175 5151
rect 17233 5117 17267 5151
rect 17693 5117 17727 5151
rect 17785 5117 17819 5151
rect 18337 5117 18371 5151
rect 20453 5117 20487 5151
rect 21281 5117 21315 5151
rect 4261 5049 4295 5083
rect 5365 5049 5399 5083
rect 11529 5049 11563 5083
rect 12909 5049 12943 5083
rect 14841 5049 14875 5083
rect 16497 5049 16531 5083
rect 19809 5049 19843 5083
rect 2513 4981 2547 5015
rect 6377 4981 6411 5015
rect 7665 4981 7699 5015
rect 10425 4981 10459 5015
rect 11897 4981 11931 5015
rect 13001 4981 13035 5015
rect 18245 4981 18279 5015
rect 19717 4981 19751 5015
rect 1593 4777 1627 4811
rect 1961 4777 1995 4811
rect 3433 4777 3467 4811
rect 5365 4777 5399 4811
rect 8953 4777 8987 4811
rect 9781 4777 9815 4811
rect 11713 4777 11747 4811
rect 12909 4777 12943 4811
rect 16773 4777 16807 4811
rect 18337 4777 18371 4811
rect 20637 4777 20671 4811
rect 1869 4709 1903 4743
rect 8677 4709 8711 4743
rect 18245 4709 18279 4743
rect 19993 4709 20027 4743
rect 4169 4641 4203 4675
rect 4721 4641 4755 4675
rect 5825 4641 5859 4675
rect 5917 4641 5951 4675
rect 6653 4641 6687 4675
rect 6929 4641 6963 4675
rect 8125 4641 8159 4675
rect 9413 4641 9447 4675
rect 9597 4641 9631 4675
rect 10241 4641 10275 4675
rect 10425 4641 10459 4675
rect 11161 4641 11195 4675
rect 12357 4641 12391 4675
rect 13645 4641 13679 4675
rect 13921 4641 13955 4675
rect 14657 4641 14691 4675
rect 18889 4641 18923 4675
rect 19441 4641 19475 4675
rect 20729 4641 20763 4675
rect 1501 4573 1535 4607
rect 3341 4573 3375 4607
rect 3617 4573 3651 4607
rect 4445 4573 4479 4607
rect 5733 4573 5767 4607
rect 6285 4573 6319 4607
rect 8493 4573 8527 4607
rect 9321 4573 9355 4607
rect 10149 4573 10183 4607
rect 10609 4573 10643 4607
rect 11805 4573 11839 4607
rect 14841 4573 14875 4607
rect 15393 4573 15427 4607
rect 16865 4573 16899 4607
rect 17121 4573 17155 4607
rect 19533 4573 19567 4607
rect 20085 4573 20119 4607
rect 20453 4573 20487 4607
rect 21005 4573 21039 4607
rect 3074 4505 3108 4539
rect 7941 4505 7975 4539
rect 11253 4505 11287 4539
rect 11345 4505 11379 4539
rect 12541 4505 12575 4539
rect 13461 4505 13495 4539
rect 14749 4505 14783 4539
rect 15660 4505 15694 4539
rect 19625 4505 19659 4539
rect 3985 4437 4019 4471
rect 4261 4437 4295 4471
rect 4813 4437 4847 4471
rect 4905 4437 4939 4471
rect 5273 4437 5307 4471
rect 6377 4437 6411 4471
rect 7573 4437 7607 4471
rect 8033 4437 8067 4471
rect 10793 4437 10827 4471
rect 11989 4437 12023 4471
rect 12449 4437 12483 4471
rect 13001 4437 13035 4471
rect 13369 4437 13403 4471
rect 14381 4437 14415 4471
rect 15209 4437 15243 4471
rect 18705 4437 18739 4471
rect 18797 4437 18831 4471
rect 20269 4437 20303 4471
rect 1869 4233 1903 4267
rect 2329 4233 2363 4267
rect 2697 4233 2731 4267
rect 3249 4233 3283 4267
rect 9137 4233 9171 4267
rect 9505 4233 9539 4267
rect 11345 4233 11379 4267
rect 13185 4233 13219 4267
rect 14841 4233 14875 4267
rect 15301 4233 15335 4267
rect 16865 4233 16899 4267
rect 17785 4233 17819 4267
rect 20545 4233 20579 4267
rect 5825 4165 5859 4199
rect 6653 4165 6687 4199
rect 6837 4165 6871 4199
rect 9689 4165 9723 4199
rect 15669 4165 15703 4199
rect 18613 4165 18647 4199
rect 19073 4165 19107 4199
rect 21097 4165 21131 4199
rect 21465 4165 21499 4199
rect 1961 4097 1995 4131
rect 2789 4097 2823 4131
rect 4373 4097 4407 4131
rect 5181 4097 5215 4131
rect 7196 4097 7230 4131
rect 8493 4097 8527 4131
rect 10221 4097 10255 4131
rect 11529 4097 11563 4131
rect 11805 4097 11839 4131
rect 12173 4097 12207 4131
rect 12633 4097 12667 4131
rect 13093 4097 13127 4131
rect 14013 4097 14047 4131
rect 16313 4097 16347 4131
rect 16681 4097 16715 4131
rect 17049 4097 17083 4131
rect 17693 4097 17727 4131
rect 19809 4097 19843 4131
rect 20085 4097 20119 4131
rect 20361 4097 20395 4131
rect 20821 4097 20855 4131
rect 1685 4029 1719 4063
rect 2605 4029 2639 4063
rect 4629 4029 4663 4063
rect 4721 4029 4755 4063
rect 5917 4029 5951 4063
rect 6101 4029 6135 4063
rect 6377 4029 6411 4063
rect 6929 4029 6963 4063
rect 8953 4029 8987 4063
rect 9045 4029 9079 4063
rect 9965 4029 9999 4063
rect 12909 4029 12943 4063
rect 14105 4029 14139 4063
rect 14197 4029 14231 4063
rect 14933 4029 14967 4063
rect 15025 4029 15059 4063
rect 15761 4029 15795 4063
rect 15945 4029 15979 4063
rect 17601 4029 17635 4063
rect 18705 4029 18739 4063
rect 18797 4029 18831 4063
rect 20913 4029 20947 4063
rect 3157 3961 3191 3995
rect 5365 3961 5399 3995
rect 11989 3961 12023 3995
rect 13553 3961 13587 3995
rect 17325 3961 17359 3995
rect 18153 3961 18187 3995
rect 18245 3961 18279 3995
rect 19625 3961 19659 3995
rect 19993 3961 20027 3995
rect 20269 3961 20303 3995
rect 1501 3893 1535 3927
rect 4997 3893 5031 3927
rect 5457 3893 5491 3927
rect 8309 3893 8343 3927
rect 8585 3893 8619 3927
rect 9781 3893 9815 3927
rect 11713 3893 11747 3927
rect 12357 3893 12391 3927
rect 12449 3893 12483 3927
rect 13645 3893 13679 3927
rect 14473 3893 14507 3927
rect 16221 3893 16255 3927
rect 19441 3893 19475 3927
rect 20637 3893 20671 3927
rect 21373 3893 21407 3927
rect 1961 3689 1995 3723
rect 3893 3689 3927 3723
rect 6193 3689 6227 3723
rect 7113 3689 7147 3723
rect 8769 3689 8803 3723
rect 10149 3689 10183 3723
rect 11713 3689 11747 3723
rect 11897 3689 11931 3723
rect 15117 3689 15151 3723
rect 16497 3689 16531 3723
rect 16865 3689 16899 3723
rect 18153 3689 18187 3723
rect 18981 3689 19015 3723
rect 19993 3689 20027 3723
rect 1685 3621 1719 3655
rect 19349 3621 19383 3655
rect 19625 3621 19659 3655
rect 2605 3553 2639 3587
rect 3433 3553 3467 3587
rect 4169 3553 4203 3587
rect 6469 3553 6503 3587
rect 6653 3553 6687 3587
rect 7297 3553 7331 3587
rect 8217 3553 8251 3587
rect 8309 3553 8343 3587
rect 12541 3553 12575 3587
rect 14565 3553 14599 3587
rect 14749 3553 14783 3587
rect 15761 3553 15795 3587
rect 16773 3553 16807 3587
rect 17509 3553 17543 3587
rect 18337 3553 18371 3587
rect 18521 3553 18555 3587
rect 1501 3485 1535 3519
rect 1777 3485 1811 3519
rect 2421 3485 2455 3519
rect 4261 3485 4295 3519
rect 4813 3485 4847 3519
rect 5080 3485 5114 3519
rect 6745 3485 6779 3519
rect 7481 3485 7515 3519
rect 8953 3485 8987 3519
rect 9229 3485 9263 3519
rect 10333 3485 10367 3519
rect 12265 3485 12299 3519
rect 14933 3485 14967 3519
rect 15485 3485 15519 3519
rect 15945 3485 15979 3519
rect 16221 3485 16255 3519
rect 17141 3485 17175 3519
rect 17785 3485 17819 3519
rect 18613 3485 18647 3519
rect 19441 3485 19475 3519
rect 19717 3485 19751 3519
rect 20177 3485 20211 3519
rect 20637 3485 20671 3519
rect 20729 3485 20763 3519
rect 21005 3485 21039 3519
rect 8401 3417 8435 3451
rect 10057 3417 10091 3451
rect 10600 3417 10634 3451
rect 11989 3417 12023 3451
rect 12808 3417 12842 3451
rect 15577 3417 15611 3451
rect 2053 3349 2087 3383
rect 2513 3349 2547 3383
rect 2881 3349 2915 3383
rect 3249 3349 3283 3383
rect 3341 3349 3375 3383
rect 4353 3349 4387 3383
rect 4721 3349 4755 3383
rect 7573 3349 7607 3383
rect 7941 3349 7975 3383
rect 12449 3349 12483 3383
rect 13921 3349 13955 3383
rect 14105 3349 14139 3383
rect 14473 3349 14507 3383
rect 16129 3349 16163 3383
rect 16405 3349 16439 3383
rect 17325 3349 17359 3383
rect 17693 3349 17727 3383
rect 19901 3349 19935 3383
rect 20453 3349 20487 3383
rect 2421 3145 2455 3179
rect 2697 3145 2731 3179
rect 2973 3145 3007 3179
rect 5365 3145 5399 3179
rect 5733 3145 5767 3179
rect 5825 3145 5859 3179
rect 6377 3145 6411 3179
rect 9689 3145 9723 3179
rect 10057 3145 10091 3179
rect 10149 3145 10183 3179
rect 10517 3145 10551 3179
rect 10977 3145 11011 3179
rect 11897 3145 11931 3179
rect 13921 3145 13955 3179
rect 14289 3145 14323 3179
rect 15485 3145 15519 3179
rect 17417 3145 17451 3179
rect 18705 3145 18739 3179
rect 3433 3077 3467 3111
rect 7849 3077 7883 3111
rect 8033 3077 8067 3111
rect 8462 3077 8496 3111
rect 11989 3077 12023 3111
rect 13562 3077 13596 3111
rect 1961 3009 1995 3043
rect 2513 3009 2547 3043
rect 2789 3009 2823 3043
rect 3893 3009 3927 3043
rect 4160 3009 4194 3043
rect 7501 3009 7535 3043
rect 8217 3009 8251 3043
rect 10885 3009 10919 3043
rect 14933 3009 14967 3043
rect 15025 3009 15059 3043
rect 15301 3009 15335 3043
rect 15577 3009 15611 3043
rect 16129 3009 16163 3043
rect 16221 3009 16255 3043
rect 16681 3009 16715 3043
rect 16957 3009 16991 3043
rect 17233 3009 17267 3043
rect 17509 3009 17543 3043
rect 17785 3009 17819 3043
rect 18153 3009 18187 3043
rect 18521 3009 18555 3043
rect 18889 3009 18923 3043
rect 19257 3009 19291 3043
rect 19625 3009 19659 3043
rect 20269 3009 20303 3043
rect 20361 3009 20395 3043
rect 20729 3009 20763 3043
rect 2237 2941 2271 2975
rect 3249 2941 3283 2975
rect 3341 2941 3375 2975
rect 5917 2941 5951 2975
rect 7757 2941 7791 2975
rect 10333 2941 10367 2975
rect 11069 2941 11103 2975
rect 12081 2941 12115 2975
rect 13829 2941 13863 2975
rect 14381 2941 14415 2975
rect 14565 2941 14599 2975
rect 21005 2941 21039 2975
rect 9597 2873 9631 2907
rect 12449 2873 12483 2907
rect 16865 2873 16899 2907
rect 17693 2873 17727 2907
rect 18337 2873 18371 2907
rect 20085 2873 20119 2907
rect 3801 2805 3835 2839
rect 5273 2805 5307 2839
rect 11529 2805 11563 2839
rect 14749 2805 14783 2839
rect 15209 2805 15243 2839
rect 15761 2805 15795 2839
rect 15945 2805 15979 2839
rect 16405 2805 16439 2839
rect 17141 2805 17175 2839
rect 17969 2805 18003 2839
rect 19073 2805 19107 2839
rect 19441 2805 19475 2839
rect 19809 2805 19843 2839
rect 20545 2805 20579 2839
rect 5089 2601 5123 2635
rect 7113 2601 7147 2635
rect 7941 2601 7975 2635
rect 9045 2601 9079 2635
rect 11713 2601 11747 2635
rect 12541 2601 12575 2635
rect 15025 2601 15059 2635
rect 17233 2601 17267 2635
rect 18705 2601 18739 2635
rect 19073 2601 19107 2635
rect 19717 2601 19751 2635
rect 3617 2533 3651 2567
rect 14565 2533 14599 2567
rect 17969 2533 18003 2567
rect 19441 2533 19475 2567
rect 1961 2465 1995 2499
rect 3157 2465 3191 2499
rect 4629 2465 4663 2499
rect 4813 2465 4847 2499
rect 5733 2465 5767 2499
rect 5917 2465 5951 2499
rect 6561 2465 6595 2499
rect 7389 2465 7423 2499
rect 8585 2465 8619 2499
rect 10793 2465 10827 2499
rect 13093 2465 13127 2499
rect 20729 2465 20763 2499
rect 21005 2465 21039 2499
rect 2237 2397 2271 2431
rect 2881 2397 2915 2431
rect 4353 2397 4387 2431
rect 6745 2397 6779 2431
rect 7481 2397 7515 2431
rect 7573 2397 7607 2431
rect 9229 2397 9263 2431
rect 9873 2397 9907 2431
rect 10149 2397 10183 2431
rect 10701 2397 10735 2431
rect 11529 2397 11563 2431
rect 12081 2397 12115 2431
rect 12173 2397 12207 2431
rect 12909 2397 12943 2431
rect 13001 2397 13035 2431
rect 13369 2397 13403 2431
rect 13737 2397 13771 2431
rect 14105 2397 14139 2431
rect 14749 2397 14783 2431
rect 14841 2397 14875 2431
rect 15209 2397 15243 2431
rect 15577 2397 15611 2431
rect 15945 2397 15979 2431
rect 16313 2397 16347 2431
rect 16681 2397 16715 2431
rect 17049 2397 17083 2431
rect 17417 2397 17451 2431
rect 17785 2397 17819 2431
rect 18153 2397 18187 2431
rect 18521 2397 18555 2431
rect 18889 2397 18923 2431
rect 19257 2397 19291 2431
rect 20361 2397 20395 2431
rect 20637 2397 20671 2431
rect 3433 2329 3467 2363
rect 4997 2329 5031 2363
rect 6653 2329 6687 2363
rect 8401 2329 8435 2363
rect 11253 2329 11287 2363
rect 5273 2261 5307 2295
rect 5641 2261 5675 2295
rect 6193 2261 6227 2295
rect 8033 2261 8067 2295
rect 8493 2261 8527 2295
rect 10241 2261 10275 2295
rect 10609 2261 10643 2295
rect 11161 2261 11195 2295
rect 11897 2261 11931 2295
rect 12357 2261 12391 2295
rect 13553 2261 13587 2295
rect 13921 2261 13955 2295
rect 14289 2261 14323 2295
rect 15393 2261 15427 2295
rect 15761 2261 15795 2295
rect 16129 2261 16163 2295
rect 16497 2261 16531 2295
rect 16865 2261 16899 2295
rect 17601 2261 17635 2295
rect 18337 2261 18371 2295
<< metal1 >>
rect 1026 21088 1032 21140
rect 1084 21128 1090 21140
rect 11054 21128 11060 21140
rect 1084 21100 11060 21128
rect 1084 21088 1090 21100
rect 11054 21088 11060 21100
rect 11112 21088 11118 21140
rect 1670 21020 1676 21072
rect 1728 21060 1734 21072
rect 17770 21060 17776 21072
rect 1728 21032 17776 21060
rect 1728 21020 1734 21032
rect 17770 21020 17776 21032
rect 17828 21020 17834 21072
rect 4522 20884 4528 20936
rect 4580 20924 4586 20936
rect 11146 20924 11152 20936
rect 4580 20896 11152 20924
rect 4580 20884 4586 20896
rect 11146 20884 11152 20896
rect 11204 20884 11210 20936
rect 2130 20816 2136 20868
rect 2188 20856 2194 20868
rect 17218 20856 17224 20868
rect 2188 20828 17224 20856
rect 2188 20816 2194 20828
rect 17218 20816 17224 20828
rect 17276 20816 17282 20868
rect 3970 20748 3976 20800
rect 4028 20788 4034 20800
rect 6730 20788 6736 20800
rect 4028 20760 6736 20788
rect 4028 20748 4034 20760
rect 6730 20748 6736 20760
rect 6788 20788 6794 20800
rect 10042 20788 10048 20800
rect 6788 20760 10048 20788
rect 6788 20748 6794 20760
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 1854 20584 1860 20596
rect 1815 20556 1860 20584
rect 1854 20544 1860 20556
rect 1912 20544 1918 20596
rect 2222 20584 2228 20596
rect 2183 20556 2228 20584
rect 2222 20544 2228 20556
rect 2280 20544 2286 20596
rect 2700 20556 4108 20584
rect 2700 20525 2728 20556
rect 2685 20519 2743 20525
rect 2685 20485 2697 20519
rect 2731 20485 2743 20519
rect 2685 20479 2743 20485
rect 3053 20519 3111 20525
rect 3053 20485 3065 20519
rect 3099 20516 3111 20519
rect 3970 20516 3976 20528
rect 3099 20488 3976 20516
rect 3099 20485 3111 20488
rect 3053 20479 3111 20485
rect 3970 20476 3976 20488
rect 4028 20476 4034 20528
rect 4080 20516 4108 20556
rect 4338 20544 4344 20596
rect 4396 20584 4402 20596
rect 5810 20584 5816 20596
rect 4396 20556 5816 20584
rect 4396 20544 4402 20556
rect 5810 20544 5816 20556
rect 5868 20584 5874 20596
rect 6822 20584 6828 20596
rect 5868 20556 6828 20584
rect 5868 20544 5874 20556
rect 6822 20544 6828 20556
rect 6880 20544 6886 20596
rect 10321 20587 10379 20593
rect 10321 20553 10333 20587
rect 10367 20584 10379 20587
rect 10870 20584 10876 20596
rect 10367 20556 10876 20584
rect 10367 20553 10379 20556
rect 10321 20547 10379 20553
rect 10870 20544 10876 20556
rect 10928 20544 10934 20596
rect 11698 20544 11704 20596
rect 11756 20584 11762 20596
rect 11885 20587 11943 20593
rect 11885 20584 11897 20587
rect 11756 20556 11897 20584
rect 11756 20544 11762 20556
rect 11885 20553 11897 20556
rect 11931 20553 11943 20587
rect 11885 20547 11943 20553
rect 11974 20544 11980 20596
rect 12032 20584 12038 20596
rect 12253 20587 12311 20593
rect 12253 20584 12265 20587
rect 12032 20556 12265 20584
rect 12032 20544 12038 20556
rect 12253 20553 12265 20556
rect 12299 20553 12311 20587
rect 12253 20547 12311 20553
rect 12434 20544 12440 20596
rect 12492 20584 12498 20596
rect 12621 20587 12679 20593
rect 12621 20584 12633 20587
rect 12492 20556 12633 20584
rect 12492 20544 12498 20556
rect 12621 20553 12633 20556
rect 12667 20553 12679 20587
rect 12621 20547 12679 20553
rect 12710 20544 12716 20596
rect 12768 20584 12774 20596
rect 12897 20587 12955 20593
rect 12897 20584 12909 20587
rect 12768 20556 12909 20584
rect 12768 20544 12774 20556
rect 12897 20553 12909 20556
rect 12943 20553 12955 20587
rect 12897 20547 12955 20553
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 13357 20587 13415 20593
rect 13357 20584 13369 20587
rect 13136 20556 13369 20584
rect 13136 20544 13142 20556
rect 13357 20553 13369 20556
rect 13403 20553 13415 20587
rect 13357 20547 13415 20553
rect 13446 20544 13452 20596
rect 13504 20584 13510 20596
rect 13633 20587 13691 20593
rect 13633 20584 13645 20587
rect 13504 20556 13645 20584
rect 13504 20544 13510 20556
rect 13633 20553 13645 20556
rect 13679 20553 13691 20587
rect 13633 20547 13691 20553
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 13872 20556 14289 20584
rect 13872 20544 13878 20556
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 14550 20544 14556 20596
rect 14608 20584 14614 20596
rect 15013 20587 15071 20593
rect 15013 20584 15025 20587
rect 14608 20556 15025 20584
rect 14608 20544 14614 20556
rect 15013 20553 15025 20556
rect 15059 20553 15071 20587
rect 15013 20547 15071 20553
rect 15194 20544 15200 20596
rect 15252 20584 15258 20596
rect 15381 20587 15439 20593
rect 15381 20584 15393 20587
rect 15252 20556 15393 20584
rect 15252 20544 15258 20556
rect 15381 20553 15393 20556
rect 15427 20553 15439 20587
rect 15381 20547 15439 20553
rect 15654 20544 15660 20596
rect 15712 20584 15718 20596
rect 16117 20587 16175 20593
rect 16117 20584 16129 20587
rect 15712 20556 16129 20584
rect 15712 20544 15718 20556
rect 16117 20553 16129 20556
rect 16163 20553 16175 20587
rect 16117 20547 16175 20553
rect 16574 20544 16580 20596
rect 16632 20584 16638 20596
rect 16853 20587 16911 20593
rect 16853 20584 16865 20587
rect 16632 20556 16865 20584
rect 16632 20544 16638 20556
rect 16853 20553 16865 20556
rect 16899 20553 16911 20587
rect 16853 20547 16911 20553
rect 16942 20544 16948 20596
rect 17000 20584 17006 20596
rect 17221 20587 17279 20593
rect 17221 20584 17233 20587
rect 17000 20556 17233 20584
rect 17000 20544 17006 20556
rect 17221 20553 17233 20556
rect 17267 20553 17279 20587
rect 17221 20547 17279 20553
rect 17957 20587 18015 20593
rect 17957 20553 17969 20587
rect 18003 20553 18015 20587
rect 19518 20584 19524 20596
rect 19479 20556 19524 20584
rect 17957 20547 18015 20553
rect 5166 20516 5172 20528
rect 4080 20488 5172 20516
rect 5166 20476 5172 20488
rect 5224 20476 5230 20528
rect 5258 20476 5264 20528
rect 5316 20516 5322 20528
rect 6638 20516 6644 20528
rect 5316 20488 6644 20516
rect 5316 20476 5322 20488
rect 6638 20476 6644 20488
rect 6696 20476 6702 20528
rect 7282 20516 7288 20528
rect 6748 20488 7288 20516
rect 1670 20448 1676 20460
rect 1631 20420 1676 20448
rect 1670 20408 1676 20420
rect 1728 20408 1734 20460
rect 2041 20451 2099 20457
rect 2041 20417 2053 20451
rect 2087 20448 2099 20451
rect 2130 20448 2136 20460
rect 2087 20420 2136 20448
rect 2087 20417 2099 20420
rect 2041 20411 2099 20417
rect 2130 20408 2136 20420
rect 2188 20408 2194 20460
rect 2406 20448 2412 20460
rect 2367 20420 2412 20448
rect 2406 20408 2412 20420
rect 2464 20408 2470 20460
rect 3510 20448 3516 20460
rect 3471 20420 3516 20448
rect 3510 20408 3516 20420
rect 3568 20408 3574 20460
rect 3602 20408 3608 20460
rect 3660 20448 3666 20460
rect 4062 20448 4068 20460
rect 3660 20420 4068 20448
rect 3660 20408 3666 20420
rect 4062 20408 4068 20420
rect 4120 20448 4126 20460
rect 4617 20451 4675 20457
rect 4617 20448 4629 20451
rect 4120 20420 4629 20448
rect 4120 20408 4126 20420
rect 4617 20417 4629 20420
rect 4663 20417 4675 20451
rect 4617 20411 4675 20417
rect 4709 20451 4767 20457
rect 4709 20417 4721 20451
rect 4755 20417 4767 20451
rect 5074 20448 5080 20460
rect 5035 20420 5080 20448
rect 4709 20411 4767 20417
rect 4341 20383 4399 20389
rect 4341 20349 4353 20383
rect 4387 20380 4399 20383
rect 4522 20380 4528 20392
rect 4387 20352 4528 20380
rect 4387 20349 4399 20352
rect 4341 20343 4399 20349
rect 4522 20340 4528 20352
rect 4580 20340 4586 20392
rect 4724 20380 4752 20411
rect 5074 20408 5080 20420
rect 5132 20408 5138 20460
rect 5350 20408 5356 20460
rect 5408 20448 5414 20460
rect 6549 20451 6607 20457
rect 5408 20420 6224 20448
rect 5408 20408 5414 20420
rect 5442 20380 5448 20392
rect 4724 20352 5448 20380
rect 5442 20340 5448 20352
rect 5500 20340 5506 20392
rect 6196 20389 6224 20420
rect 6549 20417 6561 20451
rect 6595 20448 6607 20451
rect 6748 20448 6776 20488
rect 7282 20476 7288 20488
rect 7340 20476 7346 20528
rect 7466 20476 7472 20528
rect 7524 20516 7530 20528
rect 9033 20519 9091 20525
rect 7524 20488 8524 20516
rect 7524 20476 7530 20488
rect 6595 20420 6776 20448
rect 6595 20417 6607 20420
rect 6549 20411 6607 20417
rect 6822 20408 6828 20460
rect 6880 20448 6886 20460
rect 6917 20451 6975 20457
rect 6917 20448 6929 20451
rect 6880 20420 6929 20448
rect 6880 20408 6886 20420
rect 6917 20417 6929 20420
rect 6963 20417 6975 20451
rect 6917 20411 6975 20417
rect 7009 20451 7067 20457
rect 7009 20417 7021 20451
rect 7055 20448 7067 20451
rect 7374 20448 7380 20460
rect 7055 20420 7380 20448
rect 7055 20417 7067 20420
rect 7009 20411 7067 20417
rect 7374 20408 7380 20420
rect 7432 20408 7438 20460
rect 7561 20451 7619 20457
rect 7561 20417 7573 20451
rect 7607 20448 7619 20451
rect 7650 20448 7656 20460
rect 7607 20420 7656 20448
rect 7607 20417 7619 20420
rect 7561 20411 7619 20417
rect 7650 20408 7656 20420
rect 7708 20408 7714 20460
rect 7745 20451 7803 20457
rect 7745 20417 7757 20451
rect 7791 20448 7803 20451
rect 8202 20448 8208 20460
rect 7791 20420 8208 20448
rect 7791 20417 7803 20420
rect 7745 20411 7803 20417
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 8496 20457 8524 20488
rect 9033 20485 9045 20519
rect 9079 20516 9091 20519
rect 9079 20488 10548 20516
rect 9079 20485 9091 20488
rect 9033 20479 9091 20485
rect 10520 20460 10548 20488
rect 15746 20476 15752 20528
rect 15804 20516 15810 20528
rect 15804 20488 16528 20516
rect 15804 20476 15810 20488
rect 8481 20451 8539 20457
rect 8481 20417 8493 20451
rect 8527 20417 8539 20451
rect 8481 20411 8539 20417
rect 9306 20408 9312 20460
rect 9364 20448 9370 20460
rect 9953 20451 10011 20457
rect 9953 20448 9965 20451
rect 9364 20420 9965 20448
rect 9364 20408 9370 20420
rect 9953 20417 9965 20420
rect 9999 20417 10011 20451
rect 10134 20448 10140 20460
rect 10095 20420 10140 20448
rect 9953 20411 10011 20417
rect 5905 20383 5963 20389
rect 5905 20349 5917 20383
rect 5951 20349 5963 20383
rect 5905 20343 5963 20349
rect 6181 20383 6239 20389
rect 6181 20349 6193 20383
rect 6227 20380 6239 20383
rect 6638 20380 6644 20392
rect 6227 20352 6644 20380
rect 6227 20349 6239 20352
rect 6181 20343 6239 20349
rect 2866 20272 2872 20324
rect 2924 20312 2930 20324
rect 3970 20312 3976 20324
rect 2924 20284 3976 20312
rect 2924 20272 2930 20284
rect 3970 20272 3976 20284
rect 4028 20272 4034 20324
rect 4890 20312 4896 20324
rect 4851 20284 4896 20312
rect 4890 20272 4896 20284
rect 4948 20272 4954 20324
rect 5261 20315 5319 20321
rect 5261 20281 5273 20315
rect 5307 20312 5319 20315
rect 5350 20312 5356 20324
rect 5307 20284 5356 20312
rect 5307 20281 5319 20284
rect 5261 20275 5319 20281
rect 5350 20272 5356 20284
rect 5408 20272 5414 20324
rect 5920 20312 5948 20343
rect 6638 20340 6644 20352
rect 6696 20340 6702 20392
rect 6733 20383 6791 20389
rect 6733 20349 6745 20383
rect 6779 20380 6791 20383
rect 6779 20352 7052 20380
rect 6779 20349 6791 20352
rect 6733 20343 6791 20349
rect 6822 20312 6828 20324
rect 5920 20284 6828 20312
rect 6822 20272 6828 20284
rect 6880 20272 6886 20324
rect 1486 20244 1492 20256
rect 1447 20216 1492 20244
rect 1486 20204 1492 20216
rect 1544 20204 1550 20256
rect 2774 20204 2780 20256
rect 2832 20244 2838 20256
rect 2832 20216 2877 20244
rect 2832 20204 2838 20216
rect 2958 20204 2964 20256
rect 3016 20244 3022 20256
rect 3145 20247 3203 20253
rect 3145 20244 3157 20247
rect 3016 20216 3157 20244
rect 3016 20204 3022 20216
rect 3145 20213 3157 20216
rect 3191 20213 3203 20247
rect 3418 20244 3424 20256
rect 3379 20216 3424 20244
rect 3145 20207 3203 20213
rect 3418 20204 3424 20216
rect 3476 20204 3482 20256
rect 5718 20204 5724 20256
rect 5776 20244 5782 20256
rect 6365 20247 6423 20253
rect 6365 20244 6377 20247
rect 5776 20216 6377 20244
rect 5776 20204 5782 20216
rect 6365 20213 6377 20216
rect 6411 20213 6423 20247
rect 7024 20244 7052 20352
rect 7098 20340 7104 20392
rect 7156 20380 7162 20392
rect 7156 20352 8616 20380
rect 7156 20340 7162 20352
rect 7377 20315 7435 20321
rect 7377 20281 7389 20315
rect 7423 20312 7435 20315
rect 7423 20284 8524 20312
rect 7423 20281 7435 20284
rect 7377 20275 7435 20281
rect 8496 20256 8524 20284
rect 8386 20244 8392 20256
rect 7024 20216 8392 20244
rect 6365 20207 6423 20213
rect 8386 20204 8392 20216
rect 8444 20204 8450 20256
rect 8478 20204 8484 20256
rect 8536 20204 8542 20256
rect 8588 20244 8616 20352
rect 8662 20340 8668 20392
rect 8720 20380 8726 20392
rect 8757 20383 8815 20389
rect 8757 20380 8769 20383
rect 8720 20352 8769 20380
rect 8720 20340 8726 20352
rect 8757 20349 8769 20352
rect 8803 20380 8815 20383
rect 9122 20380 9128 20392
rect 8803 20352 9128 20380
rect 8803 20349 8815 20352
rect 8757 20343 8815 20349
rect 9122 20340 9128 20352
rect 9180 20340 9186 20392
rect 9674 20380 9680 20392
rect 9635 20352 9680 20380
rect 9674 20340 9680 20352
rect 9732 20340 9738 20392
rect 9968 20312 9996 20411
rect 10134 20408 10140 20420
rect 10192 20408 10198 20460
rect 10502 20448 10508 20460
rect 10463 20420 10508 20448
rect 10502 20408 10508 20420
rect 10560 20408 10566 20460
rect 10594 20408 10600 20460
rect 10652 20448 10658 20460
rect 11701 20451 11759 20457
rect 11701 20448 11713 20451
rect 10652 20420 11713 20448
rect 10652 20408 10658 20420
rect 11701 20417 11713 20420
rect 11747 20417 11759 20451
rect 12066 20448 12072 20460
rect 12027 20420 12072 20448
rect 11701 20411 11759 20417
rect 12066 20408 12072 20420
rect 12124 20408 12130 20460
rect 12158 20408 12164 20460
rect 12216 20448 12222 20460
rect 12437 20451 12495 20457
rect 12437 20448 12449 20451
rect 12216 20420 12449 20448
rect 12216 20408 12222 20420
rect 12437 20417 12449 20420
rect 12483 20417 12495 20451
rect 13078 20448 13084 20460
rect 13039 20420 13084 20448
rect 12437 20411 12495 20417
rect 13078 20408 13084 20420
rect 13136 20408 13142 20460
rect 13170 20408 13176 20460
rect 13228 20448 13234 20460
rect 13228 20420 13273 20448
rect 13228 20408 13234 20420
rect 13630 20408 13636 20460
rect 13688 20448 13694 20460
rect 13817 20451 13875 20457
rect 13817 20448 13829 20451
rect 13688 20420 13829 20448
rect 13688 20408 13694 20420
rect 13817 20417 13829 20420
rect 13863 20417 13875 20451
rect 13817 20411 13875 20417
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20417 14151 20451
rect 14093 20411 14151 20417
rect 10781 20383 10839 20389
rect 10781 20349 10793 20383
rect 10827 20380 10839 20383
rect 10827 20352 12434 20380
rect 10827 20349 10839 20352
rect 10781 20343 10839 20349
rect 10962 20312 10968 20324
rect 9968 20284 10968 20312
rect 10962 20272 10968 20284
rect 11020 20272 11026 20324
rect 12406 20312 12434 20352
rect 13354 20340 13360 20392
rect 13412 20380 13418 20392
rect 14108 20380 14136 20411
rect 14274 20408 14280 20460
rect 14332 20448 14338 20460
rect 14461 20451 14519 20457
rect 14461 20448 14473 20451
rect 14332 20420 14473 20448
rect 14332 20408 14338 20420
rect 14461 20417 14473 20420
rect 14507 20417 14519 20451
rect 14461 20411 14519 20417
rect 14642 20408 14648 20460
rect 14700 20448 14706 20460
rect 14829 20451 14887 20457
rect 14829 20448 14841 20451
rect 14700 20420 14841 20448
rect 14700 20408 14706 20420
rect 14829 20417 14841 20420
rect 14875 20417 14887 20451
rect 14829 20411 14887 20417
rect 14918 20408 14924 20460
rect 14976 20448 14982 20460
rect 15197 20451 15255 20457
rect 15197 20448 15209 20451
rect 14976 20420 15209 20448
rect 14976 20408 14982 20420
rect 15197 20417 15209 20420
rect 15243 20417 15255 20451
rect 15562 20448 15568 20460
rect 15523 20420 15568 20448
rect 15197 20411 15255 20417
rect 15562 20408 15568 20420
rect 15620 20408 15626 20460
rect 15930 20448 15936 20460
rect 15891 20420 15936 20448
rect 15930 20408 15936 20420
rect 15988 20408 15994 20460
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20417 16359 20451
rect 16301 20411 16359 20417
rect 13412 20352 14136 20380
rect 13412 20340 13418 20352
rect 13538 20312 13544 20324
rect 11532 20284 12020 20312
rect 12406 20284 13544 20312
rect 11532 20244 11560 20284
rect 8588 20216 11560 20244
rect 11609 20247 11667 20253
rect 11609 20213 11621 20247
rect 11655 20244 11667 20247
rect 11882 20244 11888 20256
rect 11655 20216 11888 20244
rect 11655 20213 11667 20216
rect 11609 20207 11667 20213
rect 11882 20204 11888 20216
rect 11940 20204 11946 20256
rect 11992 20244 12020 20284
rect 13538 20272 13544 20284
rect 13596 20272 13602 20324
rect 14182 20272 14188 20324
rect 14240 20312 14246 20324
rect 14645 20315 14703 20321
rect 14645 20312 14657 20315
rect 14240 20284 14657 20312
rect 14240 20272 14246 20284
rect 14645 20281 14657 20284
rect 14691 20281 14703 20315
rect 14645 20275 14703 20281
rect 15286 20272 15292 20324
rect 15344 20312 15350 20324
rect 15749 20315 15807 20321
rect 15749 20312 15761 20315
rect 15344 20284 15761 20312
rect 15344 20272 15350 20284
rect 15749 20281 15761 20284
rect 15795 20281 15807 20315
rect 16316 20312 16344 20411
rect 16500 20380 16528 20488
rect 17126 20476 17132 20528
rect 17184 20516 17190 20528
rect 17972 20516 18000 20547
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 19978 20584 19984 20596
rect 19939 20556 19984 20584
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 20346 20584 20352 20596
rect 20307 20556 20352 20584
rect 20346 20544 20352 20556
rect 20404 20544 20410 20596
rect 21174 20544 21180 20596
rect 21232 20584 21238 20596
rect 21453 20587 21511 20593
rect 21453 20584 21465 20587
rect 21232 20556 21465 20584
rect 21232 20544 21238 20556
rect 21453 20553 21465 20556
rect 21499 20553 21511 20587
rect 21453 20547 21511 20553
rect 17184 20488 18000 20516
rect 18984 20488 19840 20516
rect 17184 20476 17190 20488
rect 16666 20448 16672 20460
rect 16627 20420 16672 20448
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 16942 20408 16948 20460
rect 17000 20448 17006 20460
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 17000 20420 17049 20448
rect 17000 20408 17006 20420
rect 17037 20417 17049 20420
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 17405 20451 17463 20457
rect 17405 20417 17417 20451
rect 17451 20417 17463 20451
rect 17405 20411 17463 20417
rect 17420 20380 17448 20411
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 17773 20451 17831 20457
rect 17773 20448 17785 20451
rect 17644 20420 17785 20448
rect 17644 20408 17650 20420
rect 17773 20417 17785 20420
rect 17819 20417 17831 20451
rect 17773 20411 17831 20417
rect 17954 20408 17960 20460
rect 18012 20448 18018 20460
rect 18141 20451 18199 20457
rect 18141 20448 18153 20451
rect 18012 20420 18153 20448
rect 18012 20408 18018 20420
rect 18141 20417 18153 20420
rect 18187 20417 18199 20451
rect 18141 20411 18199 20417
rect 18230 20408 18236 20460
rect 18288 20448 18294 20460
rect 18509 20451 18567 20457
rect 18509 20448 18521 20451
rect 18288 20420 18521 20448
rect 18288 20408 18294 20420
rect 18509 20417 18521 20420
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 18690 20408 18696 20460
rect 18748 20448 18754 20460
rect 18877 20451 18935 20457
rect 18877 20448 18889 20451
rect 18748 20420 18889 20448
rect 18748 20408 18754 20420
rect 18877 20417 18889 20420
rect 18923 20417 18935 20451
rect 18877 20411 18935 20417
rect 16500 20352 17448 20380
rect 16316 20284 16620 20312
rect 15749 20275 15807 20281
rect 13814 20244 13820 20256
rect 11992 20216 13820 20244
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 16390 20204 16396 20256
rect 16448 20244 16454 20256
rect 16485 20247 16543 20253
rect 16485 20244 16497 20247
rect 16448 20216 16497 20244
rect 16448 20204 16454 20216
rect 16485 20213 16497 20216
rect 16531 20213 16543 20247
rect 16592 20244 16620 20284
rect 17034 20272 17040 20324
rect 17092 20312 17098 20324
rect 17589 20315 17647 20321
rect 17589 20312 17601 20315
rect 17092 20284 17601 20312
rect 17092 20272 17098 20284
rect 17589 20281 17601 20284
rect 17635 20281 17647 20315
rect 17589 20275 17647 20281
rect 17862 20272 17868 20324
rect 17920 20312 17926 20324
rect 18693 20315 18751 20321
rect 18693 20312 18705 20315
rect 17920 20284 18705 20312
rect 17920 20272 17926 20284
rect 18693 20281 18705 20284
rect 18739 20281 18751 20315
rect 18693 20275 18751 20281
rect 18874 20272 18880 20324
rect 18932 20312 18938 20324
rect 18984 20312 19012 20488
rect 19702 20448 19708 20460
rect 19663 20420 19708 20448
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 19812 20457 19840 20488
rect 19797 20451 19855 20457
rect 19797 20417 19809 20451
rect 19843 20417 19855 20451
rect 19797 20411 19855 20417
rect 20165 20451 20223 20457
rect 20165 20417 20177 20451
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20417 20591 20451
rect 20533 20411 20591 20417
rect 20901 20451 20959 20457
rect 20901 20417 20913 20451
rect 20947 20417 20959 20451
rect 20901 20411 20959 20417
rect 20180 20380 20208 20411
rect 20548 20380 20576 20411
rect 19076 20352 20208 20380
rect 20272 20352 20576 20380
rect 20916 20380 20944 20411
rect 20990 20408 20996 20460
rect 21048 20448 21054 20460
rect 21269 20451 21327 20457
rect 21269 20448 21281 20451
rect 21048 20420 21281 20448
rect 21048 20408 21054 20420
rect 21269 20417 21281 20420
rect 21315 20417 21327 20451
rect 21269 20411 21327 20417
rect 21358 20380 21364 20392
rect 20916 20352 21364 20380
rect 19076 20321 19104 20352
rect 18932 20284 19012 20312
rect 19061 20315 19119 20321
rect 18932 20272 18938 20284
rect 19061 20281 19073 20315
rect 19107 20281 19119 20315
rect 19061 20275 19119 20281
rect 19337 20315 19395 20321
rect 19337 20281 19349 20315
rect 19383 20312 19395 20315
rect 19610 20312 19616 20324
rect 19383 20284 19616 20312
rect 19383 20281 19395 20284
rect 19337 20275 19395 20281
rect 19610 20272 19616 20284
rect 19668 20272 19674 20324
rect 17402 20244 17408 20256
rect 16592 20216 17408 20244
rect 16485 20207 16543 20213
rect 17402 20204 17408 20216
rect 17460 20204 17466 20256
rect 17494 20204 17500 20256
rect 17552 20244 17558 20256
rect 18325 20247 18383 20253
rect 18325 20244 18337 20247
rect 17552 20216 18337 20244
rect 17552 20204 17558 20216
rect 18325 20213 18337 20216
rect 18371 20213 18383 20247
rect 18325 20207 18383 20213
rect 18414 20204 18420 20256
rect 18472 20244 18478 20256
rect 20272 20244 20300 20352
rect 21358 20340 21364 20352
rect 21416 20340 21422 20392
rect 20717 20315 20775 20321
rect 20717 20281 20729 20315
rect 20763 20312 20775 20315
rect 21542 20312 21548 20324
rect 20763 20284 21548 20312
rect 20763 20281 20775 20284
rect 20717 20275 20775 20281
rect 21542 20272 21548 20284
rect 21600 20272 21606 20324
rect 21082 20244 21088 20256
rect 18472 20216 20300 20244
rect 21043 20216 21088 20244
rect 18472 20204 18478 20216
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 1946 20000 1952 20052
rect 2004 20040 2010 20052
rect 2225 20043 2283 20049
rect 2225 20040 2237 20043
rect 2004 20012 2237 20040
rect 2004 20000 2010 20012
rect 2225 20009 2237 20012
rect 2271 20009 2283 20043
rect 2225 20003 2283 20009
rect 2593 20043 2651 20049
rect 2593 20009 2605 20043
rect 2639 20040 2651 20043
rect 3878 20040 3884 20052
rect 2639 20012 3884 20040
rect 2639 20009 2651 20012
rect 2593 20003 2651 20009
rect 3878 20000 3884 20012
rect 3936 20000 3942 20052
rect 4065 20043 4123 20049
rect 4065 20009 4077 20043
rect 4111 20040 4123 20043
rect 4111 20012 5488 20040
rect 4111 20009 4123 20012
rect 4065 20003 4123 20009
rect 2866 19972 2872 19984
rect 2827 19944 2872 19972
rect 2866 19932 2872 19944
rect 2924 19932 2930 19984
rect 3234 19972 3240 19984
rect 3195 19944 3240 19972
rect 3234 19932 3240 19944
rect 3292 19932 3298 19984
rect 3326 19932 3332 19984
rect 3384 19972 3390 19984
rect 3605 19975 3663 19981
rect 3605 19972 3617 19975
rect 3384 19944 3617 19972
rect 3384 19932 3390 19944
rect 3605 19941 3617 19944
rect 3651 19941 3663 19975
rect 3605 19935 3663 19941
rect 5460 19904 5488 20012
rect 5534 20000 5540 20052
rect 5592 20040 5598 20052
rect 6730 20040 6736 20052
rect 5592 20012 6736 20040
rect 5592 20000 5598 20012
rect 6730 20000 6736 20012
rect 6788 20040 6794 20052
rect 7101 20043 7159 20049
rect 7101 20040 7113 20043
rect 6788 20012 7113 20040
rect 6788 20000 6794 20012
rect 7101 20009 7113 20012
rect 7147 20009 7159 20043
rect 7101 20003 7159 20009
rect 9125 20043 9183 20049
rect 9125 20009 9137 20043
rect 9171 20040 9183 20043
rect 10594 20040 10600 20052
rect 9171 20012 10600 20040
rect 9171 20009 9183 20012
rect 9125 20003 9183 20009
rect 10594 20000 10600 20012
rect 10652 20000 10658 20052
rect 11238 20000 11244 20052
rect 11296 20040 11302 20052
rect 11425 20043 11483 20049
rect 11425 20040 11437 20043
rect 11296 20012 11437 20040
rect 11296 20000 11302 20012
rect 11425 20009 11437 20012
rect 11471 20009 11483 20043
rect 12066 20040 12072 20052
rect 12027 20012 12072 20040
rect 11425 20003 11483 20009
rect 12066 20000 12072 20012
rect 12124 20000 12130 20052
rect 12529 20043 12587 20049
rect 12529 20009 12541 20043
rect 12575 20040 12587 20043
rect 13078 20040 13084 20052
rect 12575 20012 12664 20040
rect 13039 20012 13084 20040
rect 12575 20009 12587 20012
rect 12529 20003 12587 20009
rect 8386 19932 8392 19984
rect 8444 19972 8450 19984
rect 8570 19972 8576 19984
rect 8444 19944 8576 19972
rect 8444 19932 8450 19944
rect 8570 19932 8576 19944
rect 8628 19972 8634 19984
rect 9585 19975 9643 19981
rect 9585 19972 9597 19975
rect 8628 19944 9597 19972
rect 8628 19932 8634 19944
rect 9585 19941 9597 19944
rect 9631 19941 9643 19975
rect 12434 19972 12440 19984
rect 9585 19935 9643 19941
rect 10980 19944 12440 19972
rect 7742 19904 7748 19916
rect 5460 19876 5856 19904
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19836 1731 19839
rect 1762 19836 1768 19848
rect 1719 19808 1768 19836
rect 1719 19805 1731 19808
rect 1673 19799 1731 19805
rect 1762 19796 1768 19808
rect 1820 19796 1826 19848
rect 2041 19839 2099 19845
rect 2041 19805 2053 19839
rect 2087 19805 2099 19839
rect 2406 19836 2412 19848
rect 2367 19808 2412 19836
rect 2041 19799 2099 19805
rect 1394 19728 1400 19780
rect 1452 19768 1458 19780
rect 2056 19768 2084 19799
rect 2406 19796 2412 19808
rect 2464 19796 2470 19848
rect 2590 19796 2596 19848
rect 2648 19836 2654 19848
rect 2685 19839 2743 19845
rect 2685 19836 2697 19839
rect 2648 19808 2697 19836
rect 2648 19796 2654 19808
rect 2685 19805 2697 19808
rect 2731 19805 2743 19839
rect 2685 19799 2743 19805
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19836 3111 19839
rect 4249 19839 4307 19845
rect 3099 19808 3924 19836
rect 3099 19805 3111 19808
rect 3053 19799 3111 19805
rect 1452 19740 2084 19768
rect 1452 19728 1458 19740
rect 2222 19728 2228 19780
rect 2280 19768 2286 19780
rect 3326 19768 3332 19780
rect 2280 19740 3332 19768
rect 2280 19728 2286 19740
rect 3326 19728 3332 19740
rect 3384 19728 3390 19780
rect 3421 19771 3479 19777
rect 3421 19737 3433 19771
rect 3467 19768 3479 19771
rect 3602 19768 3608 19780
rect 3467 19740 3608 19768
rect 3467 19737 3479 19740
rect 3421 19731 3479 19737
rect 3602 19728 3608 19740
rect 3660 19728 3666 19780
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 1854 19700 1860 19712
rect 1815 19672 1860 19700
rect 1854 19660 1860 19672
rect 1912 19660 1918 19712
rect 3896 19700 3924 19808
rect 4249 19805 4261 19839
rect 4295 19836 4307 19839
rect 5718 19836 5724 19848
rect 4295 19808 5724 19836
rect 4295 19805 4307 19808
rect 4249 19799 4307 19805
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 5828 19836 5856 19876
rect 6840 19876 7748 19904
rect 5828 19808 6684 19836
rect 3973 19771 4031 19777
rect 3973 19737 3985 19771
rect 4019 19768 4031 19771
rect 4516 19771 4574 19777
rect 4019 19740 4476 19768
rect 4019 19737 4031 19740
rect 3973 19731 4031 19737
rect 4246 19700 4252 19712
rect 3896 19672 4252 19700
rect 4246 19660 4252 19672
rect 4304 19660 4310 19712
rect 4448 19700 4476 19740
rect 4516 19737 4528 19771
rect 4562 19768 4574 19771
rect 4706 19768 4712 19780
rect 4562 19740 4712 19768
rect 4562 19737 4574 19740
rect 4516 19731 4574 19737
rect 4706 19728 4712 19740
rect 4764 19728 4770 19780
rect 5534 19768 5540 19780
rect 5460 19740 5540 19768
rect 5460 19700 5488 19740
rect 5534 19728 5540 19740
rect 5592 19728 5598 19780
rect 5966 19771 6024 19777
rect 5966 19768 5978 19771
rect 5644 19740 5978 19768
rect 5644 19712 5672 19740
rect 5966 19737 5978 19740
rect 6012 19737 6024 19771
rect 6656 19768 6684 19808
rect 6840 19768 6868 19876
rect 7742 19864 7748 19876
rect 7800 19904 7806 19916
rect 7837 19907 7895 19913
rect 7837 19904 7849 19907
rect 7800 19876 7849 19904
rect 7800 19864 7806 19876
rect 7837 19873 7849 19876
rect 7883 19873 7895 19907
rect 7837 19867 7895 19873
rect 8205 19907 8263 19913
rect 8205 19873 8217 19907
rect 8251 19904 8263 19907
rect 8662 19904 8668 19916
rect 8251 19876 8668 19904
rect 8251 19873 8263 19876
rect 8205 19867 8263 19873
rect 8662 19864 8668 19876
rect 8720 19864 8726 19916
rect 10980 19913 11008 19944
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 12636 19972 12664 20012
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 13354 20040 13360 20052
rect 13315 20012 13360 20040
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 13630 20040 13636 20052
rect 13591 20012 13636 20040
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 14274 20040 14280 20052
rect 14235 20012 14280 20040
rect 14274 20000 14280 20012
rect 14332 20000 14338 20052
rect 14642 20040 14648 20052
rect 14603 20012 14648 20040
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 14918 20040 14924 20052
rect 14879 20012 14924 20040
rect 14918 20000 14924 20012
rect 14976 20000 14982 20052
rect 15197 20043 15255 20049
rect 15197 20009 15209 20043
rect 15243 20040 15255 20043
rect 15562 20040 15568 20052
rect 15243 20012 15568 20040
rect 15243 20009 15255 20012
rect 15197 20003 15255 20009
rect 15562 20000 15568 20012
rect 15620 20000 15626 20052
rect 15746 20040 15752 20052
rect 15707 20012 15752 20040
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 16025 20043 16083 20049
rect 16025 20009 16037 20043
rect 16071 20040 16083 20043
rect 16666 20040 16672 20052
rect 16071 20012 16672 20040
rect 16071 20009 16083 20012
rect 16025 20003 16083 20009
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 16761 20043 16819 20049
rect 16761 20009 16773 20043
rect 16807 20040 16819 20043
rect 17218 20040 17224 20052
rect 16807 20012 17224 20040
rect 16807 20009 16819 20012
rect 16761 20003 16819 20009
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 17402 20000 17408 20052
rect 17460 20040 17466 20052
rect 18046 20040 18052 20052
rect 17460 20012 18052 20040
rect 17460 20000 17466 20012
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 18230 20040 18236 20052
rect 18191 20012 18236 20040
rect 18230 20000 18236 20012
rect 18288 20000 18294 20052
rect 18322 20000 18328 20052
rect 18380 20040 18386 20052
rect 18417 20043 18475 20049
rect 18417 20040 18429 20043
rect 18380 20012 18429 20040
rect 18380 20000 18386 20012
rect 18417 20009 18429 20012
rect 18463 20009 18475 20043
rect 18417 20003 18475 20009
rect 18506 20000 18512 20052
rect 18564 20040 18570 20052
rect 18693 20043 18751 20049
rect 18693 20040 18705 20043
rect 18564 20012 18705 20040
rect 18564 20000 18570 20012
rect 18693 20009 18705 20012
rect 18739 20009 18751 20043
rect 18693 20003 18751 20009
rect 18966 20000 18972 20052
rect 19024 20040 19030 20052
rect 19334 20040 19340 20052
rect 19024 20012 19340 20040
rect 19024 20000 19030 20012
rect 19334 20000 19340 20012
rect 19392 20040 19398 20052
rect 19521 20043 19579 20049
rect 19521 20040 19533 20043
rect 19392 20012 19533 20040
rect 19392 20000 19398 20012
rect 19521 20009 19533 20012
rect 19567 20009 19579 20043
rect 20530 20040 20536 20052
rect 20491 20012 20536 20040
rect 19521 20003 19579 20009
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 12805 19975 12863 19981
rect 12636 19944 12756 19972
rect 10965 19907 11023 19913
rect 10965 19873 10977 19907
rect 11011 19873 11023 19907
rect 10965 19867 11023 19873
rect 12161 19907 12219 19913
rect 12161 19873 12173 19907
rect 12207 19904 12219 19907
rect 12250 19904 12256 19916
rect 12207 19876 12256 19904
rect 12207 19873 12219 19876
rect 12161 19867 12219 19873
rect 8941 19839 8999 19845
rect 7852 19808 8524 19836
rect 6656 19740 6868 19768
rect 5966 19731 6024 19737
rect 6914 19728 6920 19780
rect 6972 19768 6978 19780
rect 7852 19768 7880 19808
rect 6972 19740 7880 19768
rect 6972 19728 6978 19740
rect 8202 19728 8208 19780
rect 8260 19768 8266 19780
rect 8389 19771 8447 19777
rect 8389 19768 8401 19771
rect 8260 19740 8401 19768
rect 8260 19728 8266 19740
rect 8389 19737 8401 19740
rect 8435 19737 8447 19771
rect 8496 19768 8524 19808
rect 8941 19805 8953 19839
rect 8987 19836 8999 19839
rect 10318 19836 10324 19848
rect 8987 19808 10324 19836
rect 8987 19805 8999 19808
rect 8941 19799 8999 19805
rect 10318 19796 10324 19808
rect 10376 19796 10382 19848
rect 10980 19836 11008 19867
rect 12250 19864 12256 19876
rect 12308 19864 12314 19916
rect 12728 19904 12756 19944
rect 12805 19941 12817 19975
rect 12851 19972 12863 19975
rect 13170 19972 13176 19984
rect 12851 19944 13176 19972
rect 12851 19941 12863 19944
rect 12805 19935 12863 19941
rect 13170 19932 13176 19944
rect 13228 19932 13234 19984
rect 13722 19972 13728 19984
rect 13683 19944 13728 19972
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 15473 19975 15531 19981
rect 15473 19941 15485 19975
rect 15519 19972 15531 19975
rect 15930 19972 15936 19984
rect 15519 19944 15936 19972
rect 15519 19941 15531 19944
rect 15473 19935 15531 19941
rect 15930 19932 15936 19944
rect 15988 19932 15994 19984
rect 16850 19932 16856 19984
rect 16908 19972 16914 19984
rect 17037 19975 17095 19981
rect 17037 19972 17049 19975
rect 16908 19944 17049 19972
rect 16908 19932 16914 19944
rect 17037 19941 17049 19944
rect 17083 19941 17095 19975
rect 17770 19972 17776 19984
rect 17731 19944 17776 19972
rect 17037 19935 17095 19941
rect 17770 19932 17776 19944
rect 17828 19932 17834 19984
rect 18598 19932 18604 19984
rect 18656 19972 18662 19984
rect 19242 19972 19248 19984
rect 18656 19944 19248 19972
rect 18656 19932 18662 19944
rect 19242 19932 19248 19944
rect 19300 19932 19306 19984
rect 18322 19904 18328 19916
rect 12728 19876 13216 19904
rect 10796 19808 11008 19836
rect 11057 19839 11115 19845
rect 9217 19771 9275 19777
rect 9217 19768 9229 19771
rect 8496 19740 9229 19768
rect 8389 19731 8447 19737
rect 9217 19737 9229 19740
rect 9263 19737 9275 19771
rect 9217 19731 9275 19737
rect 9401 19771 9459 19777
rect 9401 19737 9413 19771
rect 9447 19768 9459 19771
rect 9582 19768 9588 19780
rect 9447 19740 9588 19768
rect 9447 19737 9459 19740
rect 9401 19731 9459 19737
rect 9582 19728 9588 19740
rect 9640 19728 9646 19780
rect 10410 19728 10416 19780
rect 10468 19768 10474 19780
rect 10698 19771 10756 19777
rect 10698 19768 10710 19771
rect 10468 19740 10710 19768
rect 10468 19728 10474 19740
rect 10698 19737 10710 19740
rect 10744 19737 10756 19771
rect 10698 19731 10756 19737
rect 5626 19700 5632 19712
rect 4448 19672 5488 19700
rect 5587 19672 5632 19700
rect 5626 19660 5632 19672
rect 5684 19660 5690 19712
rect 6086 19660 6092 19712
rect 6144 19700 6150 19712
rect 7098 19700 7104 19712
rect 6144 19672 7104 19700
rect 6144 19660 6150 19672
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 7190 19660 7196 19712
rect 7248 19700 7254 19712
rect 7248 19672 7293 19700
rect 7248 19660 7254 19672
rect 7374 19660 7380 19712
rect 7432 19700 7438 19712
rect 7561 19703 7619 19709
rect 7561 19700 7573 19703
rect 7432 19672 7573 19700
rect 7432 19660 7438 19672
rect 7561 19669 7573 19672
rect 7607 19669 7619 19703
rect 7561 19663 7619 19669
rect 7653 19703 7711 19709
rect 7653 19669 7665 19703
rect 7699 19700 7711 19703
rect 8110 19700 8116 19712
rect 7699 19672 8116 19700
rect 7699 19669 7711 19672
rect 7653 19663 7711 19669
rect 8110 19660 8116 19672
rect 8168 19660 8174 19712
rect 8294 19700 8300 19712
rect 8255 19672 8300 19700
rect 8294 19660 8300 19672
rect 8352 19660 8358 19712
rect 8754 19700 8760 19712
rect 8715 19672 8760 19700
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 8846 19660 8852 19712
rect 8904 19700 8910 19712
rect 10796 19700 10824 19808
rect 11057 19805 11069 19839
rect 11103 19805 11115 19839
rect 11606 19836 11612 19848
rect 11567 19808 11612 19836
rect 11057 19799 11115 19805
rect 10870 19728 10876 19780
rect 10928 19768 10934 19780
rect 11072 19768 11100 19799
rect 11606 19796 11612 19808
rect 11664 19796 11670 19848
rect 11882 19836 11888 19848
rect 11843 19808 11888 19836
rect 11882 19796 11888 19808
rect 11940 19796 11946 19848
rect 12066 19796 12072 19848
rect 12124 19836 12130 19848
rect 12613 19839 12671 19845
rect 12124 19812 12296 19836
rect 12345 19815 12403 19821
rect 12345 19812 12357 19815
rect 12124 19808 12357 19812
rect 12124 19796 12130 19808
rect 12268 19784 12357 19808
rect 12345 19781 12357 19784
rect 12391 19781 12403 19815
rect 12613 19805 12625 19839
rect 12659 19812 12671 19839
rect 12894 19836 12900 19848
rect 12659 19805 12756 19812
rect 12855 19808 12900 19836
rect 12613 19799 12756 19805
rect 12636 19784 12756 19799
rect 12894 19796 12900 19808
rect 12952 19796 12958 19848
rect 13188 19845 13216 19876
rect 16960 19876 18328 19904
rect 13173 19839 13231 19845
rect 13173 19805 13185 19839
rect 13219 19805 13231 19839
rect 13173 19799 13231 19805
rect 13262 19796 13268 19848
rect 13320 19836 13326 19848
rect 13449 19839 13507 19845
rect 13449 19836 13461 19839
rect 13320 19808 13461 19836
rect 13320 19796 13326 19808
rect 13449 19805 13461 19808
rect 13495 19805 13507 19839
rect 13449 19799 13507 19805
rect 13909 19839 13967 19845
rect 13909 19805 13921 19839
rect 13955 19805 13967 19839
rect 14090 19836 14096 19848
rect 14051 19808 14096 19836
rect 13909 19799 13967 19805
rect 12158 19768 12164 19780
rect 10928 19740 11100 19768
rect 11256 19740 12164 19768
rect 10928 19728 10934 19740
rect 11256 19709 11284 19740
rect 12158 19728 12164 19740
rect 12216 19728 12222 19780
rect 12345 19775 12403 19781
rect 12728 19768 12756 19784
rect 12802 19768 12808 19780
rect 12728 19740 12808 19768
rect 12802 19728 12808 19740
rect 12860 19728 12866 19780
rect 8904 19672 10824 19700
rect 11241 19703 11299 19709
rect 8904 19660 8910 19672
rect 11241 19669 11253 19703
rect 11287 19669 11299 19703
rect 11790 19700 11796 19712
rect 11751 19672 11796 19700
rect 11241 19663 11299 19669
rect 11790 19660 11796 19672
rect 11848 19660 11854 19712
rect 12618 19660 12624 19712
rect 12676 19700 12682 19712
rect 13924 19700 13952 19799
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14458 19836 14464 19848
rect 14419 19808 14464 19836
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 14734 19836 14740 19848
rect 14695 19808 14740 19836
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 15010 19836 15016 19848
rect 14971 19808 15016 19836
rect 15010 19796 15016 19808
rect 15068 19796 15074 19848
rect 15194 19796 15200 19848
rect 15252 19836 15258 19848
rect 15289 19839 15347 19845
rect 15289 19836 15301 19839
rect 15252 19808 15301 19836
rect 15252 19796 15258 19808
rect 15289 19805 15301 19808
rect 15335 19805 15347 19839
rect 15562 19836 15568 19848
rect 15523 19808 15568 19836
rect 15289 19799 15347 19805
rect 15562 19796 15568 19808
rect 15620 19796 15626 19848
rect 15746 19796 15752 19848
rect 15804 19836 15810 19848
rect 16960 19845 16988 19876
rect 18322 19864 18328 19876
rect 18380 19864 18386 19916
rect 18969 19907 19027 19913
rect 18969 19904 18981 19907
rect 18432 19876 18981 19904
rect 15841 19839 15899 19845
rect 15841 19836 15853 19839
rect 15804 19808 15853 19836
rect 15804 19796 15810 19808
rect 15841 19805 15853 19808
rect 15887 19836 15899 19839
rect 16117 19839 16175 19845
rect 16117 19836 16129 19839
rect 15887 19808 16129 19836
rect 15887 19805 15899 19808
rect 15841 19799 15899 19805
rect 16117 19805 16129 19808
rect 16163 19805 16175 19839
rect 16485 19839 16543 19845
rect 16485 19836 16497 19839
rect 16117 19799 16175 19805
rect 16316 19808 16497 19836
rect 16316 19712 16344 19808
rect 16485 19805 16497 19808
rect 16531 19805 16543 19839
rect 16485 19799 16543 19805
rect 16945 19839 17003 19845
rect 16945 19805 16957 19839
rect 16991 19805 17003 19839
rect 16945 19799 17003 19805
rect 17221 19839 17279 19845
rect 17221 19805 17233 19839
rect 17267 19836 17279 19839
rect 17310 19836 17316 19848
rect 17267 19808 17316 19836
rect 17267 19805 17279 19808
rect 17221 19799 17279 19805
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19836 17739 19839
rect 17862 19836 17868 19848
rect 17727 19808 17868 19836
rect 17727 19805 17739 19808
rect 17681 19799 17739 19805
rect 17862 19796 17868 19808
rect 17920 19796 17926 19848
rect 17957 19839 18015 19845
rect 17957 19805 17969 19839
rect 18003 19805 18015 19839
rect 17957 19799 18015 19805
rect 18049 19839 18107 19845
rect 18049 19805 18061 19839
rect 18095 19836 18107 19839
rect 18138 19836 18144 19848
rect 18095 19808 18144 19836
rect 18095 19805 18107 19808
rect 18049 19799 18107 19805
rect 17586 19768 17592 19780
rect 16684 19740 17592 19768
rect 16298 19700 16304 19712
rect 12676 19672 13952 19700
rect 16259 19672 16304 19700
rect 12676 19660 12682 19672
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 16684 19709 16712 19740
rect 17586 19728 17592 19740
rect 17644 19728 17650 19780
rect 17972 19768 18000 19799
rect 18138 19796 18144 19808
rect 18196 19836 18202 19848
rect 18432 19836 18460 19876
rect 18969 19873 18981 19876
rect 19015 19873 19027 19907
rect 18969 19867 19027 19873
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 20438 19904 20444 19916
rect 19668 19876 20444 19904
rect 19668 19864 19674 19876
rect 18196 19808 18460 19836
rect 18601 19839 18659 19845
rect 18196 19796 18202 19808
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 18782 19836 18788 19848
rect 18647 19808 18788 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 18782 19796 18788 19808
rect 18840 19796 18846 19848
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19429 19839 19487 19845
rect 18923 19808 19380 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 18690 19768 18696 19780
rect 17972 19740 18696 19768
rect 18690 19728 18696 19740
rect 18748 19768 18754 19780
rect 18966 19768 18972 19780
rect 18748 19740 18972 19768
rect 18748 19728 18754 19740
rect 18966 19728 18972 19740
rect 19024 19728 19030 19780
rect 19352 19768 19380 19808
rect 19429 19805 19441 19839
rect 19475 19836 19487 19839
rect 19794 19836 19800 19848
rect 19475 19808 19800 19836
rect 19475 19805 19487 19808
rect 19429 19799 19487 19805
rect 19794 19796 19800 19808
rect 19852 19796 19858 19848
rect 20180 19845 20208 19876
rect 20438 19864 20444 19876
rect 20496 19864 20502 19916
rect 20165 19839 20223 19845
rect 20165 19805 20177 19839
rect 20211 19805 20223 19839
rect 20346 19836 20352 19848
rect 20307 19808 20352 19836
rect 20165 19799 20223 19805
rect 20346 19796 20352 19808
rect 20404 19796 20410 19848
rect 20456 19836 20484 19864
rect 20717 19839 20775 19845
rect 20717 19836 20729 19839
rect 20456 19808 20729 19836
rect 20717 19805 20729 19808
rect 20763 19805 20775 19839
rect 21266 19836 21272 19848
rect 21227 19808 21272 19836
rect 20717 19799 20775 19805
rect 21266 19796 21272 19808
rect 21324 19796 21330 19848
rect 19610 19768 19616 19780
rect 19352 19740 19616 19768
rect 19610 19728 19616 19740
rect 19668 19728 19674 19780
rect 19886 19768 19892 19780
rect 19847 19740 19892 19768
rect 19886 19728 19892 19740
rect 19944 19728 19950 19780
rect 20070 19728 20076 19780
rect 20128 19768 20134 19780
rect 20993 19771 21051 19777
rect 20993 19768 21005 19771
rect 20128 19740 21005 19768
rect 20128 19728 20134 19740
rect 20993 19737 21005 19740
rect 21039 19737 21051 19771
rect 20993 19731 21051 19737
rect 16669 19703 16727 19709
rect 16669 19669 16681 19703
rect 16715 19669 16727 19703
rect 17494 19700 17500 19712
rect 17455 19672 17500 19700
rect 16669 19663 16727 19669
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 18046 19660 18052 19712
rect 18104 19700 18110 19712
rect 19245 19703 19303 19709
rect 19245 19700 19257 19703
rect 18104 19672 19257 19700
rect 18104 19660 18110 19672
rect 19245 19669 19257 19672
rect 19291 19669 19303 19703
rect 21450 19700 21456 19712
rect 21411 19672 21456 19700
rect 19245 19663 19303 19669
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 1578 19456 1584 19508
rect 1636 19496 1642 19508
rect 1857 19499 1915 19505
rect 1857 19496 1869 19499
rect 1636 19468 1869 19496
rect 1636 19456 1642 19468
rect 1857 19465 1869 19468
rect 1903 19465 1915 19499
rect 1857 19459 1915 19465
rect 2317 19499 2375 19505
rect 2317 19465 2329 19499
rect 2363 19496 2375 19499
rect 2866 19496 2872 19508
rect 2363 19468 2872 19496
rect 2363 19465 2375 19468
rect 2317 19459 2375 19465
rect 2866 19456 2872 19468
rect 2924 19456 2930 19508
rect 3326 19456 3332 19508
rect 3384 19496 3390 19508
rect 3697 19499 3755 19505
rect 3697 19496 3709 19499
rect 3384 19468 3709 19496
rect 3384 19456 3390 19468
rect 3697 19465 3709 19468
rect 3743 19465 3755 19499
rect 3697 19459 3755 19465
rect 106 19388 112 19440
rect 164 19428 170 19440
rect 934 19428 940 19440
rect 164 19400 940 19428
rect 164 19388 170 19400
rect 934 19388 940 19400
rect 992 19388 998 19440
rect 3142 19428 3148 19440
rect 2148 19400 3148 19428
rect 198 19320 204 19372
rect 256 19360 262 19372
rect 1302 19360 1308 19372
rect 256 19332 1308 19360
rect 256 19320 262 19332
rect 1302 19320 1308 19332
rect 1360 19320 1366 19372
rect 1670 19360 1676 19372
rect 1631 19332 1676 19360
rect 1670 19320 1676 19332
rect 1728 19320 1734 19372
rect 1946 19320 1952 19372
rect 2004 19360 2010 19372
rect 2148 19369 2176 19400
rect 3142 19388 3148 19400
rect 3200 19388 3206 19440
rect 3712 19428 3740 19459
rect 3786 19456 3792 19508
rect 3844 19496 3850 19508
rect 4893 19499 4951 19505
rect 4893 19496 4905 19499
rect 3844 19468 4905 19496
rect 3844 19456 3850 19468
rect 4893 19465 4905 19468
rect 4939 19496 4951 19499
rect 5258 19496 5264 19508
rect 4939 19468 5264 19496
rect 4939 19465 4951 19468
rect 4893 19459 4951 19465
rect 5258 19456 5264 19468
rect 5316 19456 5322 19508
rect 5353 19499 5411 19505
rect 5353 19465 5365 19499
rect 5399 19496 5411 19499
rect 5721 19499 5779 19505
rect 5721 19496 5733 19499
rect 5399 19468 5733 19496
rect 5399 19465 5411 19468
rect 5353 19459 5411 19465
rect 5721 19465 5733 19468
rect 5767 19465 5779 19499
rect 5721 19459 5779 19465
rect 5813 19499 5871 19505
rect 5813 19465 5825 19499
rect 5859 19496 5871 19499
rect 5994 19496 6000 19508
rect 5859 19468 6000 19496
rect 5859 19465 5871 19468
rect 5813 19459 5871 19465
rect 5994 19456 6000 19468
rect 6052 19456 6058 19508
rect 6181 19499 6239 19505
rect 6181 19465 6193 19499
rect 6227 19496 6239 19499
rect 6733 19499 6791 19505
rect 6733 19496 6745 19499
rect 6227 19468 6745 19496
rect 6227 19465 6239 19468
rect 6181 19459 6239 19465
rect 6733 19465 6745 19468
rect 6779 19465 6791 19499
rect 6733 19459 6791 19465
rect 6825 19499 6883 19505
rect 6825 19465 6837 19499
rect 6871 19496 6883 19499
rect 7190 19496 7196 19508
rect 6871 19468 7196 19496
rect 6871 19465 6883 19468
rect 6825 19459 6883 19465
rect 7190 19456 7196 19468
rect 7248 19456 7254 19508
rect 8662 19496 8668 19508
rect 8623 19468 8668 19496
rect 8662 19456 8668 19468
rect 8720 19456 8726 19508
rect 8754 19456 8760 19508
rect 8812 19496 8818 19508
rect 10505 19499 10563 19505
rect 10505 19496 10517 19499
rect 8812 19468 10517 19496
rect 8812 19456 8818 19468
rect 10505 19465 10517 19468
rect 10551 19465 10563 19499
rect 10505 19459 10563 19465
rect 10594 19456 10600 19508
rect 10652 19496 10658 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 10652 19468 10977 19496
rect 10652 19456 10658 19468
rect 10965 19465 10977 19468
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 12066 19456 12072 19508
rect 12124 19496 12130 19508
rect 12434 19496 12440 19508
rect 12124 19468 12440 19496
rect 12124 19456 12130 19468
rect 12434 19456 12440 19468
rect 12492 19456 12498 19508
rect 12526 19456 12532 19508
rect 12584 19496 12590 19508
rect 12989 19499 13047 19505
rect 12989 19496 13001 19499
rect 12584 19468 13001 19496
rect 12584 19456 12590 19468
rect 12989 19465 13001 19468
rect 13035 19465 13047 19499
rect 12989 19459 13047 19465
rect 14001 19499 14059 19505
rect 14001 19465 14013 19499
rect 14047 19496 14059 19499
rect 14090 19496 14096 19508
rect 14047 19468 14096 19496
rect 14047 19465 14059 19468
rect 14001 19459 14059 19465
rect 14090 19456 14096 19468
rect 14148 19456 14154 19508
rect 14369 19499 14427 19505
rect 14369 19465 14381 19499
rect 14415 19496 14427 19499
rect 15010 19496 15016 19508
rect 14415 19468 15016 19496
rect 14415 19465 14427 19468
rect 14369 19459 14427 19465
rect 15010 19456 15016 19468
rect 15068 19456 15074 19508
rect 16485 19499 16543 19505
rect 16485 19465 16497 19499
rect 16531 19496 16543 19499
rect 16942 19496 16948 19508
rect 16531 19468 16948 19496
rect 16531 19465 16543 19468
rect 16485 19459 16543 19465
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 17221 19499 17279 19505
rect 17221 19465 17233 19499
rect 17267 19496 17279 19499
rect 17954 19496 17960 19508
rect 17267 19468 17960 19496
rect 17267 19465 17279 19468
rect 17221 19459 17279 19465
rect 17954 19456 17960 19468
rect 18012 19456 18018 19508
rect 18141 19499 18199 19505
rect 18141 19465 18153 19499
rect 18187 19465 18199 19499
rect 18414 19496 18420 19508
rect 18375 19468 18420 19496
rect 18141 19459 18199 19465
rect 8680 19428 8708 19456
rect 9002 19431 9060 19437
rect 9002 19428 9014 19431
rect 3712 19400 7144 19428
rect 2041 19363 2099 19369
rect 2041 19360 2053 19363
rect 2004 19332 2053 19360
rect 2004 19320 2010 19332
rect 2041 19329 2053 19332
rect 2087 19329 2099 19363
rect 2041 19323 2099 19329
rect 2133 19363 2191 19369
rect 2133 19329 2145 19363
rect 2179 19329 2191 19363
rect 2133 19323 2191 19329
rect 2777 19363 2835 19369
rect 2777 19329 2789 19363
rect 2823 19360 2835 19363
rect 2958 19360 2964 19372
rect 2823 19332 2964 19360
rect 2823 19329 2835 19332
rect 2777 19323 2835 19329
rect 2958 19320 2964 19332
rect 3016 19320 3022 19372
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19360 3663 19363
rect 4338 19360 4344 19372
rect 3651 19332 4200 19360
rect 4299 19332 4344 19360
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 2593 19295 2651 19301
rect 2593 19261 2605 19295
rect 2639 19261 2651 19295
rect 2593 19255 2651 19261
rect 2685 19295 2743 19301
rect 2685 19261 2697 19295
rect 2731 19292 2743 19295
rect 3326 19292 3332 19304
rect 2731 19264 3332 19292
rect 2731 19261 2743 19264
rect 2685 19255 2743 19261
rect 2608 19224 2636 19255
rect 3326 19252 3332 19264
rect 3384 19292 3390 19304
rect 3694 19292 3700 19304
rect 3384 19264 3700 19292
rect 3384 19252 3390 19264
rect 3694 19252 3700 19264
rect 3752 19252 3758 19304
rect 3878 19292 3884 19304
rect 3839 19264 3884 19292
rect 3878 19252 3884 19264
rect 3936 19252 3942 19304
rect 4172 19292 4200 19332
rect 4338 19320 4344 19332
rect 4396 19320 4402 19372
rect 4430 19320 4436 19372
rect 4488 19360 4494 19372
rect 4985 19363 5043 19369
rect 4985 19360 4997 19363
rect 4488 19332 4997 19360
rect 4488 19320 4494 19332
rect 4985 19329 4997 19332
rect 5031 19329 5043 19363
rect 4985 19323 5043 19329
rect 4614 19292 4620 19304
rect 4172 19264 4620 19292
rect 4614 19252 4620 19264
rect 4672 19252 4678 19304
rect 4801 19295 4859 19301
rect 4801 19261 4813 19295
rect 4847 19261 4859 19295
rect 5534 19292 5540 19304
rect 5495 19264 5540 19292
rect 4801 19255 4859 19261
rect 3896 19224 3924 19252
rect 2608 19196 3924 19224
rect 4157 19227 4215 19233
rect 4157 19193 4169 19227
rect 4203 19224 4215 19227
rect 4816 19224 4844 19255
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19261 6699 19295
rect 6641 19255 6699 19261
rect 5626 19224 5632 19236
rect 4203 19196 4752 19224
rect 4816 19196 5632 19224
rect 4203 19193 4215 19196
rect 4157 19187 4215 19193
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 3142 19156 3148 19168
rect 3103 19128 3148 19156
rect 3142 19116 3148 19128
rect 3200 19116 3206 19168
rect 3234 19116 3240 19168
rect 3292 19156 3298 19168
rect 3292 19128 3337 19156
rect 3292 19116 3298 19128
rect 4246 19116 4252 19168
rect 4304 19156 4310 19168
rect 4433 19159 4491 19165
rect 4433 19156 4445 19159
rect 4304 19128 4445 19156
rect 4304 19116 4310 19128
rect 4433 19125 4445 19128
rect 4479 19125 4491 19159
rect 4724 19156 4752 19196
rect 5626 19184 5632 19196
rect 5684 19184 5690 19236
rect 6270 19156 6276 19168
rect 4724 19128 6276 19156
rect 4433 19119 4491 19125
rect 6270 19116 6276 19128
rect 6328 19116 6334 19168
rect 6656 19156 6684 19255
rect 7116 19236 7144 19400
rect 7484 19400 8064 19428
rect 8680 19400 9014 19428
rect 7190 19320 7196 19372
rect 7248 19320 7254 19372
rect 7484 19360 7512 19400
rect 7558 19369 7564 19372
rect 7098 19184 7104 19236
rect 7156 19184 7162 19236
rect 7208 19233 7236 19320
rect 7282 19294 7288 19346
rect 7340 19334 7346 19346
rect 7392 19334 7512 19360
rect 7340 19332 7512 19334
rect 7340 19306 7420 19332
rect 7552 19323 7564 19369
rect 7616 19360 7622 19372
rect 8036 19360 8064 19400
rect 9002 19397 9014 19400
rect 9048 19397 9060 19431
rect 9002 19391 9060 19397
rect 10226 19388 10232 19440
rect 10284 19428 10290 19440
rect 11149 19431 11207 19437
rect 11149 19428 11161 19431
rect 10284 19400 11161 19428
rect 10284 19388 10290 19400
rect 11149 19397 11161 19400
rect 11195 19397 11207 19431
rect 11149 19391 11207 19397
rect 11532 19400 11928 19428
rect 8757 19363 8815 19369
rect 8757 19360 8769 19363
rect 7616 19332 7652 19360
rect 8036 19332 8769 19360
rect 7558 19320 7564 19323
rect 7616 19320 7622 19332
rect 8757 19329 8769 19332
rect 8803 19360 8815 19363
rect 8846 19360 8852 19372
rect 8803 19332 8852 19360
rect 8803 19329 8815 19332
rect 8757 19323 8815 19329
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 9766 19320 9772 19372
rect 9824 19360 9830 19372
rect 11532 19369 11560 19400
rect 10597 19363 10655 19369
rect 10597 19360 10609 19363
rect 9824 19332 10609 19360
rect 9824 19320 9830 19332
rect 10597 19329 10609 19332
rect 10643 19329 10655 19363
rect 10597 19323 10655 19329
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19329 11575 19363
rect 11517 19323 11575 19329
rect 11606 19320 11612 19372
rect 11664 19360 11670 19372
rect 11784 19363 11842 19369
rect 11784 19360 11796 19363
rect 11664 19332 11796 19360
rect 11664 19320 11670 19332
rect 11784 19329 11796 19332
rect 11830 19329 11842 19363
rect 11900 19360 11928 19400
rect 12250 19388 12256 19440
rect 12308 19428 12314 19440
rect 12894 19428 12900 19440
rect 12308 19400 12900 19428
rect 12308 19388 12314 19400
rect 12894 19388 12900 19400
rect 12952 19388 12958 19440
rect 14734 19388 14740 19440
rect 14792 19428 14798 19440
rect 14918 19428 14924 19440
rect 14792 19400 14924 19428
rect 14792 19388 14798 19400
rect 14918 19388 14924 19400
rect 14976 19388 14982 19440
rect 16390 19388 16396 19440
rect 16448 19428 16454 19440
rect 16448 19400 17172 19428
rect 16448 19388 16454 19400
rect 12066 19360 12072 19372
rect 11900 19332 12072 19360
rect 11784 19323 11842 19329
rect 12066 19320 12072 19332
rect 12124 19360 12130 19372
rect 13173 19363 13231 19369
rect 12124 19332 12572 19360
rect 12124 19320 12130 19332
rect 7340 19294 7346 19306
rect 7285 19261 7297 19294
rect 7331 19261 7343 19294
rect 10410 19292 10416 19304
rect 7285 19255 7343 19261
rect 10152 19264 10416 19292
rect 10152 19233 10180 19264
rect 10410 19252 10416 19264
rect 10468 19252 10474 19304
rect 12544 19292 12572 19332
rect 13173 19329 13185 19363
rect 13219 19329 13231 19363
rect 13173 19323 13231 19329
rect 14185 19363 14243 19369
rect 14185 19329 14197 19363
rect 14231 19360 14243 19363
rect 14366 19360 14372 19372
rect 14231 19332 14372 19360
rect 14231 19329 14243 19332
rect 14185 19323 14243 19329
rect 13078 19292 13084 19304
rect 12544 19264 13084 19292
rect 13078 19252 13084 19264
rect 13136 19292 13142 19304
rect 13188 19292 13216 19323
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19360 14519 19363
rect 14550 19360 14556 19372
rect 14507 19332 14556 19360
rect 14507 19329 14519 19332
rect 14461 19323 14519 19329
rect 14550 19320 14556 19332
rect 14608 19320 14614 19372
rect 15562 19360 15568 19372
rect 14660 19332 15568 19360
rect 13136 19264 13216 19292
rect 13136 19252 13142 19264
rect 14660 19233 14688 19332
rect 15562 19320 15568 19332
rect 15620 19320 15626 19372
rect 16114 19320 16120 19372
rect 16172 19360 16178 19372
rect 16301 19363 16359 19369
rect 16301 19360 16313 19363
rect 16172 19332 16313 19360
rect 16172 19320 16178 19332
rect 16301 19329 16313 19332
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 16850 19320 16856 19372
rect 16908 19360 16914 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16908 19332 17049 19360
rect 16908 19320 16914 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17144 19360 17172 19400
rect 17310 19388 17316 19440
rect 17368 19428 17374 19440
rect 18156 19428 18184 19459
rect 18414 19456 18420 19468
rect 18472 19456 18478 19508
rect 18782 19496 18788 19508
rect 18743 19468 18788 19496
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 18966 19456 18972 19508
rect 19024 19496 19030 19508
rect 19061 19499 19119 19505
rect 19061 19496 19073 19499
rect 19024 19468 19073 19496
rect 19024 19456 19030 19468
rect 19061 19465 19073 19468
rect 19107 19465 19119 19499
rect 19061 19459 19119 19465
rect 19426 19456 19432 19508
rect 19484 19496 19490 19508
rect 19797 19499 19855 19505
rect 19797 19496 19809 19499
rect 19484 19468 19809 19496
rect 19484 19456 19490 19468
rect 19797 19465 19809 19468
rect 19843 19465 19855 19499
rect 19797 19459 19855 19465
rect 20165 19499 20223 19505
rect 20165 19465 20177 19499
rect 20211 19496 20223 19499
rect 22278 19496 22284 19508
rect 20211 19468 22284 19496
rect 20211 19465 20223 19468
rect 20165 19459 20223 19465
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 17368 19400 18092 19428
rect 18156 19400 20392 19428
rect 17368 19388 17374 19400
rect 17954 19360 17960 19372
rect 17144 19332 17960 19360
rect 17037 19323 17095 19329
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 18064 19360 18092 19400
rect 18230 19360 18236 19372
rect 18064 19332 18236 19360
rect 18230 19320 18236 19332
rect 18288 19320 18294 19372
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 18509 19363 18567 19369
rect 18509 19360 18521 19363
rect 18380 19332 18521 19360
rect 18380 19320 18386 19332
rect 18509 19329 18521 19332
rect 18555 19329 18567 19363
rect 18509 19323 18567 19329
rect 18690 19320 18696 19372
rect 18748 19360 18754 19372
rect 18969 19363 19027 19369
rect 18969 19360 18981 19363
rect 18748 19332 18981 19360
rect 18748 19320 18754 19332
rect 18969 19329 18981 19332
rect 19015 19329 19027 19363
rect 19242 19360 19248 19372
rect 19203 19332 19248 19360
rect 18969 19323 19027 19329
rect 19242 19320 19248 19332
rect 19300 19320 19306 19372
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 19392 19332 19437 19360
rect 19392 19320 19398 19332
rect 19518 19320 19524 19372
rect 19576 19360 19582 19372
rect 19613 19363 19671 19369
rect 19613 19360 19625 19363
rect 19576 19332 19625 19360
rect 19576 19320 19582 19332
rect 19613 19329 19625 19332
rect 19659 19329 19671 19363
rect 19978 19360 19984 19372
rect 19939 19332 19984 19360
rect 19613 19323 19671 19329
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 20364 19369 20392 19400
rect 20349 19363 20407 19369
rect 20349 19329 20361 19363
rect 20395 19329 20407 19363
rect 20349 19323 20407 19329
rect 20438 19320 20444 19372
rect 20496 19360 20502 19372
rect 20622 19360 20628 19372
rect 20496 19332 20628 19360
rect 20496 19320 20502 19332
rect 20622 19320 20628 19332
rect 20680 19360 20686 19372
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 20680 19332 20729 19360
rect 20680 19320 20686 19332
rect 20717 19329 20729 19332
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 21174 19320 21180 19372
rect 21232 19360 21238 19372
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 21232 19332 21281 19360
rect 21232 19320 21238 19332
rect 21269 19329 21281 19332
rect 21315 19329 21327 19363
rect 21269 19323 21327 19329
rect 17865 19295 17923 19301
rect 17865 19261 17877 19295
rect 17911 19292 17923 19295
rect 20456 19292 20484 19320
rect 17911 19264 20484 19292
rect 17911 19261 17923 19264
rect 17865 19255 17923 19261
rect 20806 19252 20812 19304
rect 20864 19292 20870 19304
rect 20901 19295 20959 19301
rect 20901 19292 20913 19295
rect 20864 19264 20913 19292
rect 20864 19252 20870 19264
rect 20901 19261 20913 19264
rect 20947 19261 20959 19295
rect 20901 19255 20959 19261
rect 7193 19227 7251 19233
rect 7193 19193 7205 19227
rect 7239 19193 7251 19227
rect 7193 19187 7251 19193
rect 10137 19227 10195 19233
rect 10137 19193 10149 19227
rect 10183 19193 10195 19227
rect 13449 19227 13507 19233
rect 13449 19224 13461 19227
rect 10137 19187 10195 19193
rect 11072 19196 11367 19224
rect 7558 19156 7564 19168
rect 6656 19128 7564 19156
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 11072 19156 11100 19196
rect 11238 19156 11244 19168
rect 9732 19128 11100 19156
rect 11199 19128 11244 19156
rect 9732 19116 9738 19128
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 11339 19156 11367 19196
rect 12820 19196 13461 19224
rect 12820 19156 12848 19196
rect 13449 19193 13461 19196
rect 13495 19193 13507 19227
rect 13449 19187 13507 19193
rect 14645 19227 14703 19233
rect 14645 19193 14657 19227
rect 14691 19193 14703 19227
rect 15286 19224 15292 19236
rect 15247 19196 15292 19224
rect 14645 19187 14703 19193
rect 15286 19184 15292 19196
rect 15344 19184 15350 19236
rect 18693 19227 18751 19233
rect 18693 19193 18705 19227
rect 18739 19224 18751 19227
rect 18874 19224 18880 19236
rect 18739 19196 18880 19224
rect 18739 19193 18751 19196
rect 18693 19187 18751 19193
rect 18874 19184 18880 19196
rect 18932 19184 18938 19236
rect 19521 19227 19579 19233
rect 19521 19193 19533 19227
rect 19567 19224 19579 19227
rect 20254 19224 20260 19236
rect 19567 19196 20260 19224
rect 19567 19193 19579 19196
rect 19521 19187 19579 19193
rect 11339 19128 12848 19156
rect 12894 19116 12900 19168
rect 12952 19156 12958 19168
rect 12952 19128 12997 19156
rect 12952 19116 12958 19128
rect 13170 19116 13176 19168
rect 13228 19156 13234 19168
rect 13265 19159 13323 19165
rect 13265 19156 13277 19159
rect 13228 19128 13277 19156
rect 13228 19116 13234 19128
rect 13265 19125 13277 19128
rect 13311 19125 13323 19159
rect 13265 19119 13323 19125
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 13633 19159 13691 19165
rect 13633 19156 13645 19159
rect 13412 19128 13645 19156
rect 13412 19116 13418 19128
rect 13633 19125 13645 19128
rect 13679 19125 13691 19159
rect 13633 19119 13691 19125
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 14090 19156 14096 19168
rect 13780 19128 14096 19156
rect 13780 19116 13786 19128
rect 14090 19116 14096 19128
rect 14148 19116 14154 19168
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 14829 19159 14887 19165
rect 14829 19156 14841 19159
rect 14516 19128 14841 19156
rect 14516 19116 14522 19128
rect 14829 19125 14841 19128
rect 14875 19156 14887 19159
rect 15010 19156 15016 19168
rect 14875 19128 15016 19156
rect 14875 19125 14887 19128
rect 14829 19119 14887 19125
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 15194 19156 15200 19168
rect 15155 19128 15200 19156
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 15470 19156 15476 19168
rect 15431 19128 15476 19156
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 15654 19156 15660 19168
rect 15615 19128 15660 19156
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 16114 19156 16120 19168
rect 16075 19128 16120 19156
rect 16114 19116 16120 19128
rect 16172 19116 16178 19168
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 16850 19156 16856 19168
rect 16448 19128 16856 19156
rect 16448 19116 16454 19128
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 18322 19116 18328 19168
rect 18380 19156 18386 19168
rect 19536 19156 19564 19187
rect 20254 19184 20260 19196
rect 20312 19184 20318 19236
rect 20530 19224 20536 19236
rect 20491 19196 20536 19224
rect 20530 19184 20536 19196
rect 20588 19184 20594 19236
rect 18380 19128 19564 19156
rect 18380 19116 18386 19128
rect 19886 19116 19892 19168
rect 19944 19156 19950 19168
rect 20162 19156 20168 19168
rect 19944 19128 20168 19156
rect 19944 19116 19950 19128
rect 20162 19116 20168 19128
rect 20220 19116 20226 19168
rect 21450 19156 21456 19168
rect 21411 19128 21456 19156
rect 21450 19116 21456 19128
rect 21508 19116 21514 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 2133 18955 2191 18961
rect 2133 18952 2145 18955
rect 1728 18924 2145 18952
rect 1728 18912 1734 18924
rect 2133 18921 2145 18924
rect 2179 18921 2191 18955
rect 2133 18915 2191 18921
rect 2498 18912 2504 18964
rect 2556 18952 2562 18964
rect 2682 18952 2688 18964
rect 2556 18924 2688 18952
rect 2556 18912 2562 18924
rect 2682 18912 2688 18924
rect 2740 18952 2746 18964
rect 2777 18955 2835 18961
rect 2777 18952 2789 18955
rect 2740 18924 2789 18952
rect 2740 18912 2746 18924
rect 2777 18921 2789 18924
rect 2823 18921 2835 18955
rect 2777 18915 2835 18921
rect 2866 18912 2872 18964
rect 2924 18952 2930 18964
rect 5442 18952 5448 18964
rect 2924 18924 5448 18952
rect 2924 18912 2930 18924
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 5902 18912 5908 18964
rect 5960 18952 5966 18964
rect 5960 18924 7420 18952
rect 5960 18912 5966 18924
rect 1762 18844 1768 18896
rect 1820 18884 1826 18896
rect 2409 18887 2467 18893
rect 2409 18884 2421 18887
rect 1820 18856 2421 18884
rect 1820 18844 1826 18856
rect 2409 18853 2421 18856
rect 2455 18853 2467 18887
rect 2409 18847 2467 18853
rect 2958 18844 2964 18896
rect 3016 18884 3022 18896
rect 3881 18887 3939 18893
rect 3016 18856 3464 18884
rect 3016 18844 3022 18856
rect 3142 18776 3148 18828
rect 3200 18816 3206 18828
rect 3436 18825 3464 18856
rect 3881 18853 3893 18887
rect 3927 18853 3939 18887
rect 3881 18847 3939 18853
rect 3329 18819 3387 18825
rect 3329 18816 3341 18819
rect 3200 18788 3341 18816
rect 3200 18776 3206 18788
rect 3329 18785 3341 18788
rect 3375 18785 3387 18819
rect 3329 18779 3387 18785
rect 3421 18819 3479 18825
rect 3421 18785 3433 18819
rect 3467 18785 3479 18819
rect 3421 18779 3479 18785
rect 3694 18776 3700 18828
rect 3752 18816 3758 18828
rect 3896 18816 3924 18847
rect 5718 18844 5724 18896
rect 5776 18884 5782 18896
rect 7392 18884 7420 18924
rect 7558 18912 7564 18964
rect 7616 18952 7622 18964
rect 7837 18955 7895 18961
rect 7837 18952 7849 18955
rect 7616 18924 7849 18952
rect 7616 18912 7622 18924
rect 7837 18921 7849 18924
rect 7883 18921 7895 18955
rect 7837 18915 7895 18921
rect 9677 18955 9735 18961
rect 9677 18921 9689 18955
rect 9723 18952 9735 18955
rect 9766 18952 9772 18964
rect 9723 18924 9772 18952
rect 9723 18921 9735 18924
rect 9677 18915 9735 18921
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 10226 18952 10232 18964
rect 10187 18924 10232 18952
rect 10226 18912 10232 18924
rect 10284 18912 10290 18964
rect 10505 18955 10563 18961
rect 10505 18921 10517 18955
rect 10551 18952 10563 18955
rect 10870 18952 10876 18964
rect 10551 18924 10876 18952
rect 10551 18921 10563 18924
rect 10505 18915 10563 18921
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 10962 18912 10968 18964
rect 11020 18952 11026 18964
rect 13725 18955 13783 18961
rect 13725 18952 13737 18955
rect 11020 18924 12296 18952
rect 11020 18912 11026 18924
rect 5776 18856 6500 18884
rect 7392 18856 10088 18884
rect 5776 18844 5782 18856
rect 4157 18819 4215 18825
rect 4157 18816 4169 18819
rect 3752 18788 4169 18816
rect 3752 18776 3758 18788
rect 4157 18785 4169 18788
rect 4203 18785 4215 18819
rect 4157 18779 4215 18785
rect 1670 18748 1676 18760
rect 1631 18720 1676 18748
rect 1670 18708 1676 18720
rect 1728 18708 1734 18760
rect 1762 18708 1768 18760
rect 1820 18748 1826 18760
rect 2317 18751 2375 18757
rect 1820 18720 1865 18748
rect 1820 18708 1826 18720
rect 2317 18717 2329 18751
rect 2363 18717 2375 18751
rect 2590 18748 2596 18760
rect 2551 18720 2596 18748
rect 2317 18711 2375 18717
rect 2332 18680 2360 18711
rect 2590 18708 2596 18720
rect 2648 18708 2654 18760
rect 3234 18748 3240 18760
rect 3195 18720 3240 18748
rect 3234 18708 3240 18720
rect 3292 18708 3298 18760
rect 4065 18751 4123 18757
rect 4065 18717 4077 18751
rect 4111 18748 4123 18751
rect 5736 18748 5764 18844
rect 6472 18825 6500 18856
rect 6181 18819 6239 18825
rect 6181 18785 6193 18819
rect 6227 18785 6239 18819
rect 6181 18779 6239 18785
rect 6457 18819 6515 18825
rect 6457 18785 6469 18819
rect 6503 18785 6515 18819
rect 6457 18779 6515 18785
rect 4111 18720 5764 18748
rect 4111 18717 4123 18720
rect 4065 18711 4123 18717
rect 5994 18708 6000 18760
rect 6052 18748 6058 18760
rect 6089 18751 6147 18757
rect 6089 18748 6101 18751
rect 6052 18720 6101 18748
rect 6052 18708 6058 18720
rect 6089 18717 6101 18720
rect 6135 18717 6147 18751
rect 6089 18711 6147 18717
rect 2498 18680 2504 18692
rect 2332 18652 2504 18680
rect 2498 18640 2504 18652
rect 2556 18640 2562 18692
rect 4424 18683 4482 18689
rect 4424 18649 4436 18683
rect 4470 18680 4482 18683
rect 5902 18680 5908 18692
rect 4470 18652 5908 18680
rect 4470 18649 4482 18652
rect 4424 18643 4482 18649
rect 5902 18640 5908 18652
rect 5960 18680 5966 18692
rect 6196 18680 6224 18779
rect 7742 18776 7748 18828
rect 7800 18816 7806 18828
rect 8481 18819 8539 18825
rect 8481 18816 8493 18819
rect 7800 18788 8493 18816
rect 7800 18776 7806 18788
rect 8481 18785 8493 18788
rect 8527 18785 8539 18819
rect 8481 18779 8539 18785
rect 8662 18776 8668 18828
rect 8720 18816 8726 18828
rect 9033 18819 9091 18825
rect 9033 18816 9045 18819
rect 8720 18788 9045 18816
rect 8720 18776 8726 18788
rect 9033 18785 9045 18788
rect 9079 18785 9091 18819
rect 9033 18779 9091 18785
rect 6730 18757 6736 18760
rect 6724 18748 6736 18757
rect 6691 18720 6736 18748
rect 6724 18711 6736 18720
rect 6730 18708 6736 18711
rect 6788 18708 6794 18760
rect 8294 18748 8300 18760
rect 6840 18720 8300 18748
rect 5960 18652 6224 18680
rect 5960 18640 5966 18652
rect 6270 18640 6276 18692
rect 6328 18680 6334 18692
rect 6840 18680 6868 18720
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 9398 18708 9404 18760
rect 9456 18748 9462 18760
rect 9953 18751 10011 18757
rect 9953 18748 9965 18751
rect 9456 18720 9965 18748
rect 9456 18708 9462 18720
rect 9953 18717 9965 18720
rect 9999 18717 10011 18751
rect 9953 18711 10011 18717
rect 6328 18652 6868 18680
rect 6328 18640 6334 18652
rect 7006 18640 7012 18692
rect 7064 18680 7070 18692
rect 8389 18683 8447 18689
rect 8389 18680 8401 18683
rect 7064 18652 8401 18680
rect 7064 18640 7070 18652
rect 8389 18649 8401 18652
rect 8435 18649 8447 18683
rect 9766 18680 9772 18692
rect 8389 18643 8447 18649
rect 8496 18652 9536 18680
rect 9727 18652 9772 18680
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 1946 18612 1952 18624
rect 1907 18584 1952 18612
rect 1946 18572 1952 18584
rect 2004 18572 2010 18624
rect 2866 18612 2872 18624
rect 2827 18584 2872 18612
rect 2866 18572 2872 18584
rect 2924 18572 2930 18624
rect 3326 18572 3332 18624
rect 3384 18612 3390 18624
rect 4062 18612 4068 18624
rect 3384 18584 4068 18612
rect 3384 18572 3390 18584
rect 4062 18572 4068 18584
rect 4120 18572 4126 18624
rect 4706 18572 4712 18624
rect 4764 18612 4770 18624
rect 5537 18615 5595 18621
rect 5537 18612 5549 18615
rect 4764 18584 5549 18612
rect 4764 18572 4770 18584
rect 5537 18581 5549 18584
rect 5583 18581 5595 18615
rect 5537 18575 5595 18581
rect 5626 18572 5632 18624
rect 5684 18612 5690 18624
rect 5684 18584 5729 18612
rect 5684 18572 5690 18584
rect 5810 18572 5816 18624
rect 5868 18612 5874 18624
rect 5997 18615 6055 18621
rect 5997 18612 6009 18615
rect 5868 18584 6009 18612
rect 5868 18572 5874 18584
rect 5997 18581 6009 18584
rect 6043 18581 6055 18615
rect 5997 18575 6055 18581
rect 7926 18572 7932 18624
rect 7984 18612 7990 18624
rect 8294 18612 8300 18624
rect 7984 18584 8029 18612
rect 8207 18584 8300 18612
rect 7984 18572 7990 18584
rect 8294 18572 8300 18584
rect 8352 18612 8358 18624
rect 8496 18612 8524 18652
rect 8352 18584 8524 18612
rect 8352 18572 8358 18584
rect 9030 18572 9036 18624
rect 9088 18612 9094 18624
rect 9217 18615 9275 18621
rect 9217 18612 9229 18615
rect 9088 18584 9229 18612
rect 9088 18572 9094 18584
rect 9217 18581 9229 18584
rect 9263 18581 9275 18615
rect 9217 18575 9275 18581
rect 9306 18572 9312 18624
rect 9364 18612 9370 18624
rect 9508 18612 9536 18652
rect 9766 18640 9772 18652
rect 9824 18640 9830 18692
rect 10060 18680 10088 18856
rect 11977 18819 12035 18825
rect 11977 18785 11989 18819
rect 12023 18816 12035 18819
rect 12066 18816 12072 18828
rect 12023 18788 12072 18816
rect 12023 18785 12035 18788
rect 11977 18779 12035 18785
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 12161 18819 12219 18825
rect 12161 18785 12173 18819
rect 12207 18785 12219 18819
rect 12268 18816 12296 18924
rect 12406 18924 13737 18952
rect 12406 18896 12434 18924
rect 13725 18921 13737 18924
rect 13771 18921 13783 18955
rect 13725 18915 13783 18921
rect 18598 18912 18604 18964
rect 18656 18952 18662 18964
rect 19337 18955 19395 18961
rect 19337 18952 19349 18955
rect 18656 18924 19349 18952
rect 18656 18912 18662 18924
rect 19337 18921 19349 18924
rect 19383 18921 19395 18955
rect 19610 18952 19616 18964
rect 19571 18924 19616 18952
rect 19337 18915 19395 18921
rect 19610 18912 19616 18924
rect 19668 18912 19674 18964
rect 19889 18955 19947 18961
rect 19889 18921 19901 18955
rect 19935 18952 19947 18955
rect 20990 18952 20996 18964
rect 19935 18924 20996 18952
rect 19935 18921 19947 18924
rect 19889 18915 19947 18921
rect 20990 18912 20996 18924
rect 21048 18912 21054 18964
rect 12342 18844 12348 18896
rect 12400 18856 12434 18896
rect 12400 18844 12406 18856
rect 12526 18844 12532 18896
rect 12584 18884 12590 18896
rect 12897 18887 12955 18893
rect 12897 18884 12909 18887
rect 12584 18856 12909 18884
rect 12584 18844 12590 18856
rect 12897 18853 12909 18856
rect 12943 18853 12955 18887
rect 12897 18847 12955 18853
rect 19061 18887 19119 18893
rect 19061 18853 19073 18887
rect 19107 18853 19119 18887
rect 19061 18847 19119 18853
rect 13354 18816 13360 18828
rect 12268 18788 13360 18816
rect 12161 18779 12219 18785
rect 10318 18748 10324 18760
rect 10279 18720 10324 18748
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 10686 18708 10692 18760
rect 10744 18748 10750 18760
rect 12176 18748 12204 18779
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 13449 18819 13507 18825
rect 13449 18785 13461 18819
rect 13495 18785 13507 18819
rect 14274 18816 14280 18828
rect 14235 18788 14280 18816
rect 13449 18779 13507 18785
rect 10744 18720 12204 18748
rect 12345 18751 12403 18757
rect 10744 18708 10750 18720
rect 11624 18692 11652 18720
rect 12345 18717 12357 18751
rect 12391 18748 12403 18751
rect 12434 18748 12440 18760
rect 12391 18720 12440 18748
rect 12391 18717 12403 18720
rect 12345 18711 12403 18717
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 12894 18708 12900 18760
rect 12952 18748 12958 18760
rect 13464 18748 13492 18779
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 18785 18819 18843 18825
rect 18785 18785 18797 18819
rect 18831 18816 18843 18819
rect 19076 18816 19104 18847
rect 19426 18844 19432 18896
rect 19484 18884 19490 18896
rect 19484 18856 19564 18884
rect 19484 18844 19490 18856
rect 19334 18816 19340 18828
rect 18831 18788 19012 18816
rect 19076 18788 19340 18816
rect 18831 18785 18843 18788
rect 18785 18779 18843 18785
rect 12952 18720 13492 18748
rect 12952 18708 12958 18720
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14369 18751 14427 18757
rect 14369 18748 14381 18751
rect 13872 18720 14381 18748
rect 13872 18708 13878 18720
rect 14369 18717 14381 18720
rect 14415 18717 14427 18751
rect 18874 18748 18880 18760
rect 18835 18720 18880 18748
rect 14369 18711 14427 18717
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 18984 18748 19012 18788
rect 19334 18776 19340 18788
rect 19392 18776 19398 18828
rect 19426 18748 19432 18760
rect 18984 18720 19432 18748
rect 19426 18708 19432 18720
rect 19484 18708 19490 18760
rect 19536 18724 19564 18856
rect 19702 18844 19708 18896
rect 19760 18884 19766 18896
rect 19981 18887 20039 18893
rect 19981 18884 19993 18887
rect 19760 18856 19993 18884
rect 19760 18844 19766 18856
rect 19981 18853 19993 18856
rect 20027 18853 20039 18887
rect 19981 18847 20039 18853
rect 20257 18887 20315 18893
rect 20257 18853 20269 18887
rect 20303 18884 20315 18887
rect 20530 18884 20536 18896
rect 20303 18856 20536 18884
rect 20303 18853 20315 18856
rect 20257 18847 20315 18853
rect 20530 18844 20536 18856
rect 20588 18844 20594 18896
rect 20165 18751 20223 18757
rect 19705 18727 19763 18733
rect 19705 18724 19717 18727
rect 19536 18696 19717 18724
rect 19705 18693 19717 18696
rect 19751 18693 19763 18727
rect 20165 18717 20177 18751
rect 20211 18717 20223 18751
rect 20438 18748 20444 18760
rect 20399 18720 20444 18748
rect 20165 18711 20223 18717
rect 10060 18652 10824 18680
rect 10502 18612 10508 18624
rect 9364 18584 9409 18612
rect 9508 18584 10508 18612
rect 9364 18572 9370 18584
rect 10502 18572 10508 18584
rect 10560 18572 10566 18624
rect 10597 18615 10655 18621
rect 10597 18581 10609 18615
rect 10643 18612 10655 18615
rect 10686 18612 10692 18624
rect 10643 18584 10692 18612
rect 10643 18581 10655 18584
rect 10597 18575 10655 18581
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 10796 18612 10824 18652
rect 11606 18640 11612 18692
rect 11664 18640 11670 18692
rect 11732 18683 11790 18689
rect 11732 18649 11744 18683
rect 11778 18680 11790 18683
rect 11974 18680 11980 18692
rect 11778 18652 11980 18680
rect 11778 18649 11790 18652
rect 11732 18643 11790 18649
rect 11974 18640 11980 18652
rect 12032 18640 12038 18692
rect 13357 18683 13415 18689
rect 13357 18680 13369 18683
rect 12820 18652 13369 18680
rect 12342 18612 12348 18624
rect 10796 18584 12348 18612
rect 12342 18572 12348 18584
rect 12400 18572 12406 18624
rect 12437 18615 12495 18621
rect 12437 18581 12449 18615
rect 12483 18612 12495 18615
rect 12618 18612 12624 18624
rect 12483 18584 12624 18612
rect 12483 18581 12495 18584
rect 12437 18575 12495 18581
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 12820 18621 12848 18652
rect 13357 18649 13369 18652
rect 13403 18649 13415 18683
rect 13357 18643 13415 18649
rect 13446 18640 13452 18692
rect 13504 18680 13510 18692
rect 14461 18683 14519 18689
rect 14461 18680 14473 18683
rect 13504 18652 14473 18680
rect 13504 18640 13510 18652
rect 14461 18649 14473 18652
rect 14507 18649 14519 18683
rect 14461 18643 14519 18649
rect 18601 18683 18659 18689
rect 19705 18687 19763 18693
rect 18601 18649 18613 18683
rect 18647 18680 18659 18683
rect 18647 18652 19472 18680
rect 18647 18649 18659 18652
rect 18601 18643 18659 18649
rect 12805 18615 12863 18621
rect 12805 18581 12817 18615
rect 12851 18581 12863 18615
rect 13262 18612 13268 18624
rect 13223 18584 13268 18612
rect 12805 18575 12863 18581
rect 13262 18572 13268 18584
rect 13320 18572 13326 18624
rect 14826 18612 14832 18624
rect 14787 18584 14832 18612
rect 14826 18572 14832 18584
rect 14884 18572 14890 18624
rect 18417 18615 18475 18621
rect 18417 18581 18429 18615
rect 18463 18612 18475 18615
rect 19334 18612 19340 18624
rect 18463 18584 19340 18612
rect 18463 18581 18475 18584
rect 18417 18575 18475 18581
rect 19334 18572 19340 18584
rect 19392 18572 19398 18624
rect 19444 18612 19472 18652
rect 19518 18612 19524 18624
rect 19444 18584 19524 18612
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 20180 18612 20208 18711
rect 20438 18708 20444 18720
rect 20496 18708 20502 18760
rect 20622 18748 20628 18760
rect 20583 18720 20628 18748
rect 20622 18708 20628 18720
rect 20680 18708 20686 18760
rect 21269 18751 21327 18757
rect 21269 18748 21281 18751
rect 20732 18720 21281 18748
rect 20254 18640 20260 18692
rect 20312 18680 20318 18692
rect 20732 18680 20760 18720
rect 21269 18717 21281 18720
rect 21315 18717 21327 18751
rect 21269 18711 21327 18717
rect 20898 18680 20904 18692
rect 20312 18652 20760 18680
rect 20859 18652 20904 18680
rect 20312 18640 20318 18652
rect 20898 18640 20904 18652
rect 20956 18640 20962 18692
rect 20346 18612 20352 18624
rect 20180 18584 20352 18612
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 21450 18612 21456 18624
rect 21411 18584 21456 18612
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 1762 18408 1768 18420
rect 1723 18380 1768 18408
rect 1762 18368 1768 18380
rect 1820 18368 1826 18420
rect 4893 18411 4951 18417
rect 4893 18377 4905 18411
rect 4939 18408 4951 18411
rect 5626 18408 5632 18420
rect 4939 18380 5632 18408
rect 4939 18377 4951 18380
rect 4893 18371 4951 18377
rect 5626 18368 5632 18380
rect 5684 18368 5690 18420
rect 5994 18368 6000 18420
rect 6052 18408 6058 18420
rect 6181 18411 6239 18417
rect 6181 18408 6193 18411
rect 6052 18380 6193 18408
rect 6052 18368 6058 18380
rect 6181 18377 6193 18380
rect 6227 18377 6239 18411
rect 6181 18371 6239 18377
rect 6365 18411 6423 18417
rect 6365 18377 6377 18411
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 1210 18300 1216 18352
rect 1268 18340 1274 18352
rect 2774 18340 2780 18352
rect 1268 18312 2780 18340
rect 1268 18300 1274 18312
rect 2774 18300 2780 18312
rect 2832 18300 2838 18352
rect 2958 18300 2964 18352
rect 3016 18340 3022 18352
rect 3154 18343 3212 18349
rect 3154 18340 3166 18343
rect 3016 18312 3166 18340
rect 3016 18300 3022 18312
rect 3154 18309 3166 18312
rect 3200 18309 3212 18343
rect 3154 18303 3212 18309
rect 3326 18300 3332 18352
rect 3384 18340 3390 18352
rect 3789 18343 3847 18349
rect 3789 18340 3801 18343
rect 3384 18312 3801 18340
rect 3384 18300 3390 18312
rect 3789 18309 3801 18312
rect 3835 18309 3847 18343
rect 3789 18303 3847 18309
rect 5074 18300 5080 18352
rect 5132 18340 5138 18352
rect 5721 18343 5779 18349
rect 5721 18340 5733 18343
rect 5132 18312 5733 18340
rect 5132 18300 5138 18312
rect 5721 18309 5733 18312
rect 5767 18309 5779 18343
rect 5721 18303 5779 18309
rect 5813 18343 5871 18349
rect 5813 18309 5825 18343
rect 5859 18340 5871 18343
rect 6380 18340 6408 18371
rect 7282 18368 7288 18420
rect 7340 18408 7346 18420
rect 7377 18411 7435 18417
rect 7377 18408 7389 18411
rect 7340 18380 7389 18408
rect 7340 18368 7346 18380
rect 7377 18377 7389 18380
rect 7423 18377 7435 18411
rect 7377 18371 7435 18377
rect 7745 18411 7803 18417
rect 7745 18377 7757 18411
rect 7791 18408 7803 18411
rect 7926 18408 7932 18420
rect 7791 18380 7932 18408
rect 7791 18377 7803 18380
rect 7745 18371 7803 18377
rect 7926 18368 7932 18380
rect 7984 18368 7990 18420
rect 8202 18408 8208 18420
rect 8163 18380 8208 18408
rect 8202 18368 8208 18380
rect 8260 18368 8266 18420
rect 8665 18411 8723 18417
rect 8665 18377 8677 18411
rect 8711 18408 8723 18411
rect 9125 18411 9183 18417
rect 9125 18408 9137 18411
rect 8711 18380 9137 18408
rect 8711 18377 8723 18380
rect 8665 18371 8723 18377
rect 9125 18377 9137 18380
rect 9171 18377 9183 18411
rect 9125 18371 9183 18377
rect 9398 18368 9404 18420
rect 9456 18408 9462 18420
rect 11333 18411 11391 18417
rect 9456 18380 10456 18408
rect 9456 18368 9462 18380
rect 5859 18312 6408 18340
rect 5859 18309 5871 18312
rect 5813 18303 5871 18309
rect 6546 18300 6552 18352
rect 6604 18340 6610 18352
rect 10428 18340 10456 18380
rect 11333 18377 11345 18411
rect 11379 18408 11391 18411
rect 12618 18408 12624 18420
rect 11379 18380 12434 18408
rect 12579 18380 12624 18408
rect 11379 18377 11391 18380
rect 11333 18371 11391 18377
rect 6604 18312 7236 18340
rect 6604 18300 6610 18312
rect 7208 18284 7236 18312
rect 7300 18312 10364 18340
rect 10428 18312 11100 18340
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 1762 18272 1768 18284
rect 1719 18244 1768 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 1946 18272 1952 18284
rect 1907 18244 1952 18272
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 3421 18275 3479 18281
rect 3421 18241 3433 18275
rect 3467 18272 3479 18275
rect 3694 18272 3700 18284
rect 3467 18244 3700 18272
rect 3467 18241 3479 18244
rect 3421 18235 3479 18241
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 2041 18071 2099 18077
rect 2041 18037 2053 18071
rect 2087 18068 2099 18071
rect 2130 18068 2136 18080
rect 2087 18040 2136 18068
rect 2087 18037 2099 18040
rect 2041 18031 2099 18037
rect 2130 18028 2136 18040
rect 2188 18028 2194 18080
rect 3234 18028 3240 18080
rect 3292 18068 3298 18080
rect 3436 18068 3464 18235
rect 3694 18232 3700 18244
rect 3752 18232 3758 18284
rect 3878 18272 3884 18284
rect 3839 18244 3884 18272
rect 3878 18232 3884 18244
rect 3936 18232 3942 18284
rect 3970 18232 3976 18284
rect 4028 18272 4034 18284
rect 4341 18275 4399 18281
rect 4341 18272 4353 18275
rect 4028 18244 4353 18272
rect 4028 18232 4034 18244
rect 4341 18241 4353 18244
rect 4387 18241 4399 18275
rect 4982 18272 4988 18284
rect 4943 18244 4988 18272
rect 4341 18235 4399 18241
rect 4982 18232 4988 18244
rect 5040 18232 5046 18284
rect 5442 18232 5448 18284
rect 5500 18272 5506 18284
rect 6362 18272 6368 18284
rect 5500 18244 6368 18272
rect 5500 18232 5506 18244
rect 6362 18232 6368 18244
rect 6420 18272 6426 18284
rect 6733 18275 6791 18281
rect 6733 18272 6745 18275
rect 6420 18244 6745 18272
rect 6420 18232 6426 18244
rect 6733 18241 6745 18244
rect 6779 18241 6791 18275
rect 7006 18272 7012 18284
rect 6733 18235 6791 18241
rect 6840 18244 7012 18272
rect 3510 18164 3516 18216
rect 3568 18204 3574 18216
rect 3605 18207 3663 18213
rect 3605 18204 3617 18207
rect 3568 18176 3617 18204
rect 3568 18164 3574 18176
rect 3605 18173 3617 18176
rect 3651 18173 3663 18207
rect 4706 18204 4712 18216
rect 4667 18176 4712 18204
rect 3605 18167 3663 18173
rect 4706 18164 4712 18176
rect 4764 18164 4770 18216
rect 5534 18164 5540 18216
rect 5592 18204 5598 18216
rect 5629 18207 5687 18213
rect 5629 18204 5641 18207
rect 5592 18176 5641 18204
rect 5592 18164 5598 18176
rect 5629 18173 5641 18176
rect 5675 18173 5687 18207
rect 5629 18167 5687 18173
rect 6086 18164 6092 18216
rect 6144 18204 6150 18216
rect 6840 18213 6868 18244
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 7190 18272 7196 18284
rect 7103 18244 7196 18272
rect 7190 18232 7196 18244
rect 7248 18232 7254 18284
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6144 18176 6837 18204
rect 6144 18164 6150 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 6825 18167 6883 18173
rect 6917 18207 6975 18213
rect 6917 18173 6929 18207
rect 6963 18173 6975 18207
rect 6917 18167 6975 18173
rect 4249 18139 4307 18145
rect 4249 18105 4261 18139
rect 4295 18136 4307 18139
rect 5442 18136 5448 18148
rect 4295 18108 5448 18136
rect 4295 18105 4307 18108
rect 4249 18099 4307 18105
rect 5442 18096 5448 18108
rect 5500 18096 5506 18148
rect 6730 18096 6736 18148
rect 6788 18136 6794 18148
rect 6932 18136 6960 18167
rect 6788 18108 6960 18136
rect 6788 18096 6794 18108
rect 4522 18068 4528 18080
rect 3292 18040 3464 18068
rect 4483 18040 4528 18068
rect 3292 18028 3298 18040
rect 4522 18028 4528 18040
rect 4580 18028 4586 18080
rect 4614 18028 4620 18080
rect 4672 18068 4678 18080
rect 4890 18068 4896 18080
rect 4672 18040 4896 18068
rect 4672 18028 4678 18040
rect 4890 18028 4896 18040
rect 4948 18028 4954 18080
rect 5353 18071 5411 18077
rect 5353 18037 5365 18071
rect 5399 18068 5411 18071
rect 7300 18068 7328 18312
rect 7834 18272 7840 18284
rect 7795 18244 7840 18272
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 7926 18232 7932 18284
rect 7984 18272 7990 18284
rect 9490 18272 9496 18284
rect 7984 18244 9496 18272
rect 7984 18232 7990 18244
rect 9490 18232 9496 18244
rect 9548 18232 9554 18284
rect 10336 18281 10364 18312
rect 10137 18275 10195 18281
rect 10137 18272 10149 18275
rect 9692 18244 10149 18272
rect 7558 18204 7564 18216
rect 7519 18176 7564 18204
rect 7558 18164 7564 18176
rect 7616 18204 7622 18216
rect 8294 18204 8300 18216
rect 7616 18176 8300 18204
rect 7616 18164 7622 18176
rect 8294 18164 8300 18176
rect 8352 18204 8358 18216
rect 8389 18207 8447 18213
rect 8389 18204 8401 18207
rect 8352 18176 8401 18204
rect 8352 18164 8358 18176
rect 8389 18173 8401 18176
rect 8435 18173 8447 18207
rect 8570 18204 8576 18216
rect 8531 18176 8576 18204
rect 8389 18167 8447 18173
rect 8570 18164 8576 18176
rect 8628 18164 8634 18216
rect 9582 18204 9588 18216
rect 9543 18176 9588 18204
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 9692 18213 9720 18244
rect 10137 18241 10149 18244
rect 10183 18241 10195 18275
rect 10137 18235 10195 18241
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18241 10379 18275
rect 10321 18235 10379 18241
rect 10778 18232 10784 18284
rect 10836 18272 10842 18284
rect 10965 18275 11023 18281
rect 10965 18272 10977 18275
rect 10836 18244 10977 18272
rect 10836 18232 10842 18244
rect 10965 18241 10977 18244
rect 11011 18241 11023 18275
rect 10965 18235 11023 18241
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18173 9735 18207
rect 10686 18204 10692 18216
rect 10647 18176 10692 18204
rect 9677 18167 9735 18173
rect 9030 18136 9036 18148
rect 8991 18108 9036 18136
rect 9030 18096 9036 18108
rect 9088 18096 9094 18148
rect 9692 18136 9720 18167
rect 10686 18164 10692 18176
rect 10744 18164 10750 18216
rect 10870 18204 10876 18216
rect 10831 18176 10876 18204
rect 10870 18164 10876 18176
rect 10928 18164 10934 18216
rect 11072 18204 11100 18312
rect 11790 18300 11796 18352
rect 11848 18340 11854 18352
rect 12253 18343 12311 18349
rect 12253 18340 12265 18343
rect 11848 18312 12265 18340
rect 11848 18300 11854 18312
rect 12253 18309 12265 18312
rect 12299 18309 12311 18343
rect 12406 18340 12434 18380
rect 12618 18368 12624 18380
rect 12676 18368 12682 18420
rect 13262 18408 13268 18420
rect 12820 18380 13268 18408
rect 12820 18340 12848 18380
rect 13262 18368 13268 18380
rect 13320 18368 13326 18420
rect 17954 18368 17960 18420
rect 18012 18408 18018 18420
rect 19518 18408 19524 18420
rect 18012 18380 19524 18408
rect 18012 18368 18018 18380
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 19613 18411 19671 18417
rect 19613 18377 19625 18411
rect 19659 18408 19671 18411
rect 21634 18408 21640 18420
rect 19659 18380 21640 18408
rect 19659 18377 19671 18380
rect 19613 18371 19671 18377
rect 21634 18368 21640 18380
rect 21692 18368 21698 18420
rect 12406 18312 12848 18340
rect 12253 18303 12311 18309
rect 11606 18232 11612 18284
rect 11664 18232 11670 18284
rect 12268 18272 12296 18303
rect 12894 18300 12900 18352
rect 12952 18340 12958 18352
rect 13348 18343 13406 18349
rect 13348 18340 13360 18343
rect 12952 18312 13360 18340
rect 12952 18300 12958 18312
rect 13348 18309 13360 18312
rect 13394 18309 13406 18343
rect 16390 18340 16396 18352
rect 13348 18303 13406 18309
rect 14476 18312 16396 18340
rect 14476 18272 14504 18312
rect 16390 18300 16396 18312
rect 16448 18300 16454 18352
rect 20806 18340 20812 18352
rect 19444 18312 20812 18340
rect 12268 18244 14504 18272
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 19444 18281 19472 18312
rect 20806 18300 20812 18312
rect 20864 18300 20870 18352
rect 14737 18275 14795 18281
rect 14737 18272 14749 18275
rect 14608 18244 14749 18272
rect 14608 18232 14614 18244
rect 14737 18241 14749 18244
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 19429 18275 19487 18281
rect 19429 18241 19441 18275
rect 19475 18241 19487 18275
rect 19702 18272 19708 18284
rect 19663 18244 19708 18272
rect 19429 18235 19487 18241
rect 19702 18232 19708 18244
rect 19760 18232 19766 18284
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 20162 18272 20168 18284
rect 20027 18244 20168 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 20346 18272 20352 18284
rect 20307 18244 20352 18272
rect 20346 18232 20352 18244
rect 20404 18232 20410 18284
rect 20530 18232 20536 18284
rect 20588 18272 20594 18284
rect 20625 18275 20683 18281
rect 20625 18272 20637 18275
rect 20588 18244 20637 18272
rect 20588 18232 20594 18244
rect 20625 18241 20637 18244
rect 20671 18241 20683 18275
rect 20625 18235 20683 18241
rect 20714 18232 20720 18284
rect 20772 18272 20778 18284
rect 20901 18275 20959 18281
rect 20901 18272 20913 18275
rect 20772 18244 20913 18272
rect 20772 18232 20778 18244
rect 20901 18241 20913 18244
rect 20947 18241 20959 18275
rect 20901 18235 20959 18241
rect 20990 18232 20996 18284
rect 21048 18272 21054 18284
rect 21269 18275 21327 18281
rect 21269 18272 21281 18275
rect 21048 18244 21281 18272
rect 21048 18232 21054 18244
rect 21269 18241 21281 18244
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 11517 18207 11575 18213
rect 11517 18204 11529 18207
rect 11072 18176 11529 18204
rect 11517 18173 11529 18176
rect 11563 18173 11575 18207
rect 11624 18204 11652 18232
rect 11974 18204 11980 18216
rect 11624 18176 11980 18204
rect 11517 18167 11575 18173
rect 11974 18164 11980 18176
rect 12032 18164 12038 18216
rect 12158 18204 12164 18216
rect 12119 18176 12164 18204
rect 12158 18164 12164 18176
rect 12216 18164 12222 18216
rect 12710 18204 12716 18216
rect 12671 18176 12716 18204
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 13078 18204 13084 18216
rect 12991 18176 13084 18204
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 19334 18164 19340 18216
rect 19392 18204 19398 18216
rect 20438 18204 20444 18216
rect 19392 18176 20444 18204
rect 19392 18164 19398 18176
rect 20438 18164 20444 18176
rect 20496 18164 20502 18216
rect 21358 18204 21364 18216
rect 20732 18176 21364 18204
rect 9600 18108 9720 18136
rect 5399 18040 7328 18068
rect 5399 18037 5411 18040
rect 5353 18031 5411 18037
rect 7742 18028 7748 18080
rect 7800 18068 7806 18080
rect 9600 18068 9628 18108
rect 9858 18096 9864 18148
rect 9916 18136 9922 18148
rect 9953 18139 10011 18145
rect 9953 18136 9965 18139
rect 9916 18108 9965 18136
rect 9916 18096 9922 18108
rect 9953 18105 9965 18108
rect 9999 18105 10011 18139
rect 9953 18099 10011 18105
rect 10505 18139 10563 18145
rect 10505 18105 10517 18139
rect 10551 18136 10563 18139
rect 12526 18136 12532 18148
rect 10551 18108 12532 18136
rect 10551 18105 10563 18108
rect 10505 18099 10563 18105
rect 12526 18096 12532 18108
rect 12584 18096 12590 18148
rect 7800 18040 9628 18068
rect 7800 18028 7806 18040
rect 9674 18028 9680 18080
rect 9732 18068 9738 18080
rect 11054 18068 11060 18080
rect 9732 18040 11060 18068
rect 9732 18028 9738 18040
rect 11054 18028 11060 18040
rect 11112 18068 11118 18080
rect 11606 18068 11612 18080
rect 11112 18040 11612 18068
rect 11112 18028 11118 18040
rect 11606 18028 11612 18040
rect 11664 18028 11670 18080
rect 11698 18028 11704 18080
rect 11756 18068 11762 18080
rect 13096 18068 13124 18164
rect 14553 18139 14611 18145
rect 14553 18136 14565 18139
rect 14016 18108 14565 18136
rect 14016 18068 14044 18108
rect 14553 18105 14565 18108
rect 14599 18105 14611 18139
rect 14553 18099 14611 18105
rect 18969 18139 19027 18145
rect 18969 18105 18981 18139
rect 19015 18136 19027 18139
rect 19153 18139 19211 18145
rect 19153 18136 19165 18139
rect 19015 18108 19165 18136
rect 19015 18105 19027 18108
rect 18969 18099 19027 18105
rect 19153 18105 19165 18108
rect 19199 18136 19211 18139
rect 20622 18136 20628 18148
rect 19199 18108 20628 18136
rect 19199 18105 19211 18108
rect 19153 18099 19211 18105
rect 20622 18096 20628 18108
rect 20680 18096 20686 18148
rect 11756 18040 11801 18068
rect 13096 18040 14044 18068
rect 11756 18028 11762 18040
rect 14274 18028 14280 18080
rect 14332 18068 14338 18080
rect 14458 18068 14464 18080
rect 14332 18040 14464 18068
rect 14332 18028 14338 18040
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 15010 18028 15016 18080
rect 15068 18068 15074 18080
rect 15565 18071 15623 18077
rect 15565 18068 15577 18071
rect 15068 18040 15577 18068
rect 15068 18028 15074 18040
rect 15565 18037 15577 18040
rect 15611 18068 15623 18071
rect 16022 18068 16028 18080
rect 15611 18040 16028 18068
rect 15611 18037 15623 18040
rect 15565 18031 15623 18037
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 19337 18071 19395 18077
rect 19337 18037 19349 18071
rect 19383 18068 19395 18071
rect 19610 18068 19616 18080
rect 19383 18040 19616 18068
rect 19383 18037 19395 18040
rect 19337 18031 19395 18037
rect 19610 18028 19616 18040
rect 19668 18028 19674 18080
rect 19889 18071 19947 18077
rect 19889 18037 19901 18071
rect 19935 18068 19947 18071
rect 19978 18068 19984 18080
rect 19935 18040 19984 18068
rect 19935 18037 19947 18040
rect 19889 18031 19947 18037
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 20162 18068 20168 18080
rect 20123 18040 20168 18068
rect 20162 18028 20168 18040
rect 20220 18028 20226 18080
rect 20533 18071 20591 18077
rect 20533 18037 20545 18071
rect 20579 18068 20591 18071
rect 20732 18068 20760 18176
rect 21358 18164 21364 18176
rect 21416 18164 21422 18216
rect 21082 18136 21088 18148
rect 21043 18108 21088 18136
rect 21082 18096 21088 18108
rect 21140 18096 21146 18148
rect 20579 18040 20760 18068
rect 20809 18071 20867 18077
rect 20579 18037 20591 18040
rect 20533 18031 20591 18037
rect 20809 18037 20821 18071
rect 20855 18068 20867 18071
rect 21174 18068 21180 18080
rect 20855 18040 21180 18068
rect 20855 18037 20867 18040
rect 20809 18031 20867 18037
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 21450 18068 21456 18080
rect 21411 18040 21456 18068
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 1857 17867 1915 17873
rect 1857 17864 1869 17867
rect 1728 17836 1869 17864
rect 1728 17824 1734 17836
rect 1857 17833 1869 17836
rect 1903 17833 1915 17867
rect 1857 17827 1915 17833
rect 2406 17824 2412 17876
rect 2464 17864 2470 17876
rect 2464 17836 3372 17864
rect 2464 17824 2470 17836
rect 1670 17660 1676 17672
rect 1631 17632 1676 17660
rect 1670 17620 1676 17632
rect 1728 17620 1734 17672
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17629 2099 17663
rect 2041 17623 2099 17629
rect 2225 17663 2283 17669
rect 2225 17629 2237 17663
rect 2271 17660 2283 17663
rect 3234 17660 3240 17672
rect 2271 17632 3240 17660
rect 2271 17629 2283 17632
rect 2225 17623 2283 17629
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 2056 17524 2084 17623
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 2130 17552 2136 17604
rect 2188 17592 2194 17604
rect 2492 17595 2550 17601
rect 2492 17592 2504 17595
rect 2188 17564 2504 17592
rect 2188 17552 2194 17564
rect 2492 17561 2504 17564
rect 2538 17592 2550 17595
rect 3050 17592 3056 17604
rect 2538 17564 3056 17592
rect 2538 17561 2550 17564
rect 2492 17555 2550 17561
rect 3050 17552 3056 17564
rect 3108 17552 3114 17604
rect 3344 17592 3372 17836
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 3605 17867 3663 17873
rect 3605 17864 3617 17867
rect 3476 17836 3617 17864
rect 3476 17824 3482 17836
rect 3605 17833 3617 17836
rect 3651 17833 3663 17867
rect 4430 17864 4436 17876
rect 3605 17827 3663 17833
rect 3988 17836 4436 17864
rect 3510 17620 3516 17672
rect 3568 17660 3574 17672
rect 3988 17660 4016 17836
rect 4430 17824 4436 17836
rect 4488 17824 4494 17876
rect 4617 17867 4675 17873
rect 4617 17833 4629 17867
rect 4663 17864 4675 17867
rect 5074 17864 5080 17876
rect 4663 17836 5080 17864
rect 4663 17833 4675 17836
rect 4617 17827 4675 17833
rect 5074 17824 5080 17836
rect 5132 17824 5138 17876
rect 5902 17824 5908 17876
rect 5960 17864 5966 17876
rect 6089 17867 6147 17873
rect 6089 17864 6101 17867
rect 5960 17836 6101 17864
rect 5960 17824 5966 17836
rect 6089 17833 6101 17836
rect 6135 17833 6147 17867
rect 6089 17827 6147 17833
rect 6638 17824 6644 17876
rect 6696 17864 6702 17876
rect 7742 17864 7748 17876
rect 6696 17836 7748 17864
rect 6696 17824 6702 17836
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 8757 17867 8815 17873
rect 8757 17833 8769 17867
rect 8803 17864 8815 17867
rect 9306 17864 9312 17876
rect 8803 17836 9312 17864
rect 8803 17833 8815 17836
rect 8757 17827 8815 17833
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 9646 17836 10088 17864
rect 4448 17796 4476 17824
rect 4448 17768 4752 17796
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17728 4123 17731
rect 4430 17728 4436 17740
rect 4111 17700 4436 17728
rect 4111 17697 4123 17700
rect 4065 17691 4123 17697
rect 4430 17688 4436 17700
rect 4488 17688 4494 17740
rect 4724 17728 4752 17768
rect 6362 17756 6368 17808
rect 6420 17796 6426 17808
rect 9646 17796 9674 17836
rect 6420 17768 9674 17796
rect 9953 17799 10011 17805
rect 6420 17756 6426 17768
rect 4724 17700 4844 17728
rect 4157 17663 4215 17669
rect 4157 17660 4169 17663
rect 3568 17632 4169 17660
rect 3568 17620 3574 17632
rect 4157 17629 4169 17632
rect 4203 17629 4215 17663
rect 4157 17623 4215 17629
rect 4246 17620 4252 17672
rect 4304 17660 4310 17672
rect 4709 17663 4767 17669
rect 4709 17660 4721 17663
rect 4304 17632 4721 17660
rect 4304 17620 4310 17632
rect 4709 17629 4721 17632
rect 4755 17629 4767 17663
rect 4816 17660 4844 17700
rect 6546 17688 6552 17740
rect 6604 17728 6610 17740
rect 6733 17731 6791 17737
rect 6733 17728 6745 17731
rect 6604 17700 6745 17728
rect 6604 17688 6610 17700
rect 6733 17697 6745 17700
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 7193 17731 7251 17737
rect 7193 17697 7205 17731
rect 7239 17728 7251 17731
rect 8110 17728 8116 17740
rect 7239 17700 8116 17728
rect 7239 17697 7251 17700
rect 7193 17691 7251 17697
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 8205 17731 8263 17737
rect 8205 17697 8217 17731
rect 8251 17728 8263 17731
rect 8294 17728 8300 17740
rect 8251 17700 8300 17728
rect 8251 17697 8263 17700
rect 8205 17691 8263 17697
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 9416 17737 9444 17768
rect 9953 17765 9965 17799
rect 9999 17765 10011 17799
rect 10060 17796 10088 17836
rect 10134 17824 10140 17876
rect 10192 17864 10198 17876
rect 10410 17864 10416 17876
rect 10192 17836 10237 17864
rect 10371 17836 10416 17864
rect 10192 17824 10198 17836
rect 10410 17824 10416 17836
rect 10468 17824 10474 17876
rect 11054 17864 11060 17876
rect 11015 17836 11060 17864
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 12158 17824 12164 17876
rect 12216 17864 12222 17876
rect 12253 17867 12311 17873
rect 12253 17864 12265 17867
rect 12216 17836 12265 17864
rect 12216 17824 12222 17836
rect 12253 17833 12265 17836
rect 12299 17833 12311 17867
rect 12253 17827 12311 17833
rect 12342 17824 12348 17876
rect 12400 17864 12406 17876
rect 16298 17864 16304 17876
rect 12400 17836 16304 17864
rect 12400 17824 12406 17836
rect 16298 17824 16304 17836
rect 16356 17824 16362 17876
rect 19058 17824 19064 17876
rect 19116 17864 19122 17876
rect 20257 17867 20315 17873
rect 20257 17864 20269 17867
rect 19116 17836 20269 17864
rect 19116 17824 19122 17836
rect 20257 17833 20269 17836
rect 20303 17833 20315 17867
rect 20257 17827 20315 17833
rect 21177 17867 21235 17873
rect 21177 17833 21189 17867
rect 21223 17864 21235 17867
rect 21266 17864 21272 17876
rect 21223 17836 21272 17864
rect 21223 17833 21235 17836
rect 21177 17827 21235 17833
rect 21266 17824 21272 17836
rect 21324 17824 21330 17876
rect 10226 17796 10232 17808
rect 10060 17768 10232 17796
rect 9953 17759 10011 17765
rect 9401 17731 9459 17737
rect 9401 17697 9413 17731
rect 9447 17697 9459 17731
rect 9401 17691 9459 17697
rect 9585 17731 9643 17737
rect 9585 17697 9597 17731
rect 9631 17728 9643 17731
rect 9674 17728 9680 17740
rect 9631 17700 9680 17728
rect 9631 17697 9643 17700
rect 9585 17691 9643 17697
rect 9674 17688 9680 17700
rect 9732 17728 9738 17740
rect 9858 17728 9864 17740
rect 9732 17700 9864 17728
rect 9732 17688 9738 17700
rect 9858 17688 9864 17700
rect 9916 17688 9922 17740
rect 5258 17660 5264 17672
rect 4816 17632 5264 17660
rect 4709 17623 4767 17629
rect 5258 17620 5264 17632
rect 5316 17620 5322 17672
rect 5442 17620 5448 17672
rect 5500 17660 5506 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 5500 17632 9781 17660
rect 5500 17620 5506 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9968 17660 9996 17759
rect 10226 17756 10232 17768
rect 10284 17756 10290 17808
rect 12894 17756 12900 17808
rect 12952 17796 12958 17808
rect 13265 17799 13323 17805
rect 13265 17796 13277 17799
rect 12952 17768 13277 17796
rect 12952 17756 12958 17768
rect 13265 17765 13277 17768
rect 13311 17765 13323 17799
rect 13265 17759 13323 17765
rect 19702 17756 19708 17808
rect 19760 17796 19766 17808
rect 20717 17799 20775 17805
rect 19760 17768 20668 17796
rect 19760 17756 19766 17768
rect 10042 17688 10048 17740
rect 10100 17728 10106 17740
rect 10100 17700 11192 17728
rect 10100 17688 10106 17700
rect 10321 17663 10379 17669
rect 10321 17660 10333 17663
rect 9968 17632 10333 17660
rect 9769 17623 9827 17629
rect 10321 17629 10333 17632
rect 10367 17629 10379 17663
rect 10594 17660 10600 17672
rect 10555 17632 10600 17660
rect 10321 17623 10379 17629
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 11164 17660 11192 17700
rect 11238 17688 11244 17740
rect 11296 17728 11302 17740
rect 11514 17728 11520 17740
rect 11296 17700 11520 17728
rect 11296 17688 11302 17700
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 12158 17688 12164 17740
rect 12216 17728 12222 17740
rect 12805 17731 12863 17737
rect 12805 17728 12817 17731
rect 12216 17700 12817 17728
rect 12216 17688 12222 17700
rect 12805 17697 12817 17700
rect 12851 17697 12863 17731
rect 16298 17728 16304 17740
rect 16259 17700 16304 17728
rect 12805 17691 12863 17697
rect 16298 17688 16304 17700
rect 16356 17688 16362 17740
rect 18874 17688 18880 17740
rect 18932 17728 18938 17740
rect 20640 17728 20668 17768
rect 20717 17765 20729 17799
rect 20763 17796 20775 17799
rect 22094 17796 22100 17808
rect 20763 17768 22100 17796
rect 20763 17765 20775 17768
rect 20717 17759 20775 17765
rect 22094 17756 22100 17768
rect 22152 17756 22158 17808
rect 18932 17700 20576 17728
rect 20640 17700 20944 17728
rect 18932 17688 18938 17700
rect 11333 17663 11391 17669
rect 11333 17660 11345 17663
rect 11164 17632 11345 17660
rect 11333 17629 11345 17632
rect 11379 17660 11391 17663
rect 12621 17663 12679 17669
rect 12621 17660 12633 17663
rect 11379 17632 12633 17660
rect 11379 17629 11391 17632
rect 11333 17623 11391 17629
rect 12621 17629 12633 17632
rect 12667 17660 12679 17663
rect 13722 17660 13728 17672
rect 12667 17632 13728 17660
rect 12667 17629 12679 17632
rect 12621 17623 12679 17629
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 14182 17660 14188 17672
rect 14143 17632 14188 17660
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 14458 17669 14464 17672
rect 14452 17660 14464 17669
rect 14371 17632 14464 17660
rect 14452 17623 14464 17632
rect 14516 17660 14522 17672
rect 16316 17660 16344 17688
rect 14516 17632 16344 17660
rect 14458 17620 14464 17623
rect 14516 17620 14522 17632
rect 17402 17620 17408 17672
rect 17460 17660 17466 17672
rect 19702 17660 19708 17672
rect 17460 17632 19708 17660
rect 17460 17620 17466 17632
rect 19702 17620 19708 17632
rect 19760 17620 19766 17672
rect 20070 17660 20076 17672
rect 20031 17632 20076 17660
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 20548 17669 20576 17700
rect 20916 17669 20944 17700
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17629 20591 17663
rect 20533 17623 20591 17629
rect 20901 17663 20959 17669
rect 20901 17629 20913 17663
rect 20947 17629 20959 17663
rect 20901 17623 20959 17629
rect 20993 17663 21051 17669
rect 20993 17629 21005 17663
rect 21039 17629 21051 17663
rect 21266 17660 21272 17672
rect 21227 17632 21272 17660
rect 20993 17623 21051 17629
rect 4976 17595 5034 17601
rect 3344 17564 4936 17592
rect 2590 17524 2596 17536
rect 2056 17496 2596 17524
rect 2590 17484 2596 17496
rect 2648 17484 2654 17536
rect 2774 17484 2780 17536
rect 2832 17524 2838 17536
rect 3142 17524 3148 17536
rect 2832 17496 3148 17524
rect 2832 17484 2838 17496
rect 3142 17484 3148 17496
rect 3200 17524 3206 17536
rect 4062 17524 4068 17536
rect 3200 17496 4068 17524
rect 3200 17484 3206 17496
rect 4062 17484 4068 17496
rect 4120 17484 4126 17536
rect 4249 17527 4307 17533
rect 4249 17493 4261 17527
rect 4295 17524 4307 17527
rect 4522 17524 4528 17536
rect 4295 17496 4528 17524
rect 4295 17493 4307 17496
rect 4249 17487 4307 17493
rect 4522 17484 4528 17496
rect 4580 17484 4586 17536
rect 4908 17524 4936 17564
rect 4976 17561 4988 17595
rect 5022 17592 5034 17595
rect 5534 17592 5540 17604
rect 5022 17564 5540 17592
rect 5022 17561 5034 17564
rect 4976 17555 5034 17561
rect 5534 17552 5540 17564
rect 5592 17552 5598 17604
rect 5902 17552 5908 17604
rect 5960 17592 5966 17604
rect 5960 17564 6224 17592
rect 5960 17552 5966 17564
rect 6086 17524 6092 17536
rect 4908 17496 6092 17524
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 6196 17533 6224 17564
rect 6454 17552 6460 17604
rect 6512 17592 6518 17604
rect 6549 17595 6607 17601
rect 6549 17592 6561 17595
rect 6512 17564 6561 17592
rect 6512 17552 6518 17564
rect 6549 17561 6561 17564
rect 6595 17561 6607 17595
rect 6549 17555 6607 17561
rect 7006 17552 7012 17604
rect 7064 17592 7070 17604
rect 7377 17595 7435 17601
rect 7377 17592 7389 17595
rect 7064 17564 7389 17592
rect 7064 17552 7070 17564
rect 7377 17561 7389 17564
rect 7423 17561 7435 17595
rect 11701 17595 11759 17601
rect 11701 17592 11713 17595
rect 7377 17555 7435 17561
rect 7760 17564 10364 17592
rect 6181 17527 6239 17533
rect 6181 17493 6193 17527
rect 6227 17493 6239 17527
rect 6181 17487 6239 17493
rect 6638 17484 6644 17536
rect 6696 17524 6702 17536
rect 6696 17496 6741 17524
rect 6696 17484 6702 17496
rect 7098 17484 7104 17536
rect 7156 17524 7162 17536
rect 7760 17533 7788 17564
rect 7285 17527 7343 17533
rect 7285 17524 7297 17527
rect 7156 17496 7297 17524
rect 7156 17484 7162 17496
rect 7285 17493 7297 17496
rect 7331 17493 7343 17527
rect 7285 17487 7343 17493
rect 7745 17527 7803 17533
rect 7745 17493 7757 17527
rect 7791 17493 7803 17527
rect 7926 17524 7932 17536
rect 7887 17496 7932 17524
rect 7745 17487 7803 17493
rect 7926 17484 7932 17496
rect 7984 17484 7990 17536
rect 8202 17484 8208 17536
rect 8260 17524 8266 17536
rect 8297 17527 8355 17533
rect 8297 17524 8309 17527
rect 8260 17496 8309 17524
rect 8260 17484 8266 17496
rect 8297 17493 8309 17496
rect 8343 17493 8355 17527
rect 8297 17487 8355 17493
rect 8386 17484 8392 17536
rect 8444 17524 8450 17536
rect 8444 17496 8489 17524
rect 8444 17484 8450 17496
rect 8754 17484 8760 17536
rect 8812 17524 8818 17536
rect 8941 17527 8999 17533
rect 8941 17524 8953 17527
rect 8812 17496 8953 17524
rect 8812 17484 8818 17496
rect 8941 17493 8953 17496
rect 8987 17493 8999 17527
rect 8941 17487 8999 17493
rect 9309 17527 9367 17533
rect 9309 17493 9321 17527
rect 9355 17524 9367 17527
rect 9490 17524 9496 17536
rect 9355 17496 9496 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 9490 17484 9496 17496
rect 9548 17524 9554 17536
rect 10134 17524 10140 17536
rect 9548 17496 10140 17524
rect 9548 17484 9554 17496
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 10336 17524 10364 17564
rect 10520 17564 11713 17592
rect 10520 17524 10548 17564
rect 11701 17561 11713 17564
rect 11747 17561 11759 17595
rect 13446 17592 13452 17604
rect 13407 17564 13452 17592
rect 11701 17555 11759 17561
rect 13446 17552 13452 17564
rect 13504 17552 13510 17604
rect 13630 17552 13636 17604
rect 13688 17592 13694 17604
rect 19518 17592 19524 17604
rect 13688 17564 19524 17592
rect 13688 17552 13694 17564
rect 19518 17552 19524 17564
rect 19576 17592 19582 17604
rect 19889 17595 19947 17601
rect 19889 17592 19901 17595
rect 19576 17564 19901 17592
rect 19576 17552 19582 17564
rect 19889 17561 19901 17564
rect 19935 17592 19947 17595
rect 21008 17592 21036 17623
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 19935 17564 21036 17592
rect 19935 17561 19947 17564
rect 19889 17555 19947 17561
rect 10686 17524 10692 17536
rect 10336 17496 10548 17524
rect 10647 17496 10692 17524
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 10870 17524 10876 17536
rect 10831 17496 10876 17524
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 11790 17524 11796 17536
rect 11751 17496 11796 17524
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 12161 17527 12219 17533
rect 12161 17493 12173 17527
rect 12207 17524 12219 17527
rect 12434 17524 12440 17536
rect 12207 17496 12440 17524
rect 12207 17493 12219 17496
rect 12161 17487 12219 17493
rect 12434 17484 12440 17496
rect 12492 17484 12498 17536
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 12713 17527 12771 17533
rect 12713 17524 12725 17527
rect 12584 17496 12725 17524
rect 12584 17484 12590 17496
rect 12713 17493 12725 17496
rect 12759 17524 12771 17527
rect 13081 17527 13139 17533
rect 13081 17524 13093 17527
rect 12759 17496 13093 17524
rect 12759 17493 12771 17496
rect 12713 17487 12771 17493
rect 13081 17493 13093 17496
rect 13127 17524 13139 17527
rect 13722 17524 13728 17536
rect 13127 17496 13728 17524
rect 13127 17493 13139 17496
rect 13081 17487 13139 17493
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 14734 17484 14740 17536
rect 14792 17524 14798 17536
rect 15194 17524 15200 17536
rect 14792 17496 15200 17524
rect 14792 17484 14798 17496
rect 15194 17484 15200 17496
rect 15252 17484 15258 17536
rect 15286 17484 15292 17536
rect 15344 17524 15350 17536
rect 15565 17527 15623 17533
rect 15565 17524 15577 17527
rect 15344 17496 15577 17524
rect 15344 17484 15350 17496
rect 15565 17493 15577 17496
rect 15611 17493 15623 17527
rect 15565 17487 15623 17493
rect 15654 17484 15660 17536
rect 15712 17524 15718 17536
rect 16022 17524 16028 17536
rect 15712 17496 15757 17524
rect 15983 17496 16028 17524
rect 15712 17484 15718 17496
rect 16022 17484 16028 17496
rect 16080 17484 16086 17536
rect 16117 17527 16175 17533
rect 16117 17493 16129 17527
rect 16163 17524 16175 17527
rect 17862 17524 17868 17536
rect 16163 17496 17868 17524
rect 16163 17493 16175 17496
rect 16117 17487 16175 17493
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 20346 17524 20352 17536
rect 20307 17496 20352 17524
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 21450 17524 21456 17536
rect 21411 17496 21456 17524
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1762 17280 1768 17332
rect 1820 17320 1826 17332
rect 1857 17323 1915 17329
rect 1857 17320 1869 17323
rect 1820 17292 1869 17320
rect 1820 17280 1826 17292
rect 1857 17289 1869 17292
rect 1903 17289 1915 17323
rect 1857 17283 1915 17289
rect 1946 17280 1952 17332
rect 2004 17320 2010 17332
rect 2133 17323 2191 17329
rect 2133 17320 2145 17323
rect 2004 17292 2145 17320
rect 2004 17280 2010 17292
rect 2133 17289 2145 17292
rect 2179 17289 2191 17323
rect 2133 17283 2191 17289
rect 2685 17323 2743 17329
rect 2685 17289 2697 17323
rect 2731 17320 2743 17323
rect 2866 17320 2872 17332
rect 2731 17292 2872 17320
rect 2731 17289 2743 17292
rect 2685 17283 2743 17289
rect 2866 17280 2872 17292
rect 2924 17280 2930 17332
rect 3145 17323 3203 17329
rect 3145 17289 3157 17323
rect 3191 17320 3203 17323
rect 3326 17320 3332 17332
rect 3191 17292 3332 17320
rect 3191 17289 3203 17292
rect 3145 17283 3203 17289
rect 3326 17280 3332 17292
rect 3384 17280 3390 17332
rect 4617 17323 4675 17329
rect 4617 17289 4629 17323
rect 4663 17289 4675 17323
rect 4617 17283 4675 17289
rect 3418 17212 3424 17264
rect 3476 17261 3482 17264
rect 3476 17255 3540 17261
rect 3476 17221 3494 17255
rect 3528 17221 3540 17255
rect 3476 17215 3540 17221
rect 3476 17212 3482 17215
rect 4430 17212 4436 17264
rect 4488 17252 4494 17264
rect 4632 17252 4660 17283
rect 4982 17280 4988 17332
rect 5040 17320 5046 17332
rect 5445 17323 5503 17329
rect 5445 17320 5457 17323
rect 5040 17292 5457 17320
rect 5040 17280 5046 17292
rect 5445 17289 5457 17292
rect 5491 17289 5503 17323
rect 5902 17320 5908 17332
rect 5863 17292 5908 17320
rect 5445 17283 5503 17289
rect 5902 17280 5908 17292
rect 5960 17280 5966 17332
rect 6178 17280 6184 17332
rect 6236 17320 6242 17332
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 6236 17292 6837 17320
rect 6236 17280 6242 17292
rect 6825 17289 6837 17292
rect 6871 17289 6883 17323
rect 8202 17320 8208 17332
rect 8163 17292 8208 17320
rect 6825 17283 6883 17289
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 8570 17280 8576 17332
rect 8628 17320 8634 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8628 17292 9045 17320
rect 8628 17280 8634 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9033 17283 9091 17289
rect 9493 17323 9551 17329
rect 9493 17289 9505 17323
rect 9539 17320 9551 17323
rect 10134 17320 10140 17332
rect 9539 17292 10140 17320
rect 9539 17289 9551 17292
rect 9493 17283 9551 17289
rect 10134 17280 10140 17292
rect 10192 17320 10198 17332
rect 10686 17320 10692 17332
rect 10192 17292 10692 17320
rect 10192 17280 10198 17292
rect 10686 17280 10692 17292
rect 10744 17280 10750 17332
rect 10778 17280 10784 17332
rect 10836 17320 10842 17332
rect 11701 17323 11759 17329
rect 11701 17320 11713 17323
rect 10836 17292 11713 17320
rect 10836 17280 10842 17292
rect 11701 17289 11713 17292
rect 11747 17289 11759 17323
rect 11701 17283 11759 17289
rect 12069 17323 12127 17329
rect 12069 17289 12081 17323
rect 12115 17320 12127 17323
rect 12710 17320 12716 17332
rect 12115 17292 12716 17320
rect 12115 17289 12127 17292
rect 12069 17283 12127 17289
rect 12710 17280 12716 17292
rect 12768 17280 12774 17332
rect 12986 17320 12992 17332
rect 12947 17292 12992 17320
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 14185 17323 14243 17329
rect 14185 17289 14197 17323
rect 14231 17320 14243 17323
rect 14645 17323 14703 17329
rect 14645 17320 14657 17323
rect 14231 17292 14657 17320
rect 14231 17289 14243 17292
rect 14185 17283 14243 17289
rect 14645 17289 14657 17292
rect 14691 17289 14703 17323
rect 14645 17283 14703 17289
rect 14826 17280 14832 17332
rect 14884 17320 14890 17332
rect 15749 17323 15807 17329
rect 15749 17320 15761 17323
rect 14884 17292 15761 17320
rect 14884 17280 14890 17292
rect 15749 17289 15761 17292
rect 15795 17289 15807 17323
rect 15749 17283 15807 17289
rect 19981 17323 20039 17329
rect 19981 17289 19993 17323
rect 20027 17320 20039 17323
rect 20254 17320 20260 17332
rect 20027 17292 20260 17320
rect 20027 17289 20039 17292
rect 19981 17283 20039 17289
rect 20254 17280 20260 17292
rect 20312 17280 20318 17332
rect 20530 17280 20536 17332
rect 20588 17280 20594 17332
rect 20714 17320 20720 17332
rect 20675 17292 20720 17320
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 20990 17320 20996 17332
rect 20951 17292 20996 17320
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 6457 17255 6515 17261
rect 6457 17252 6469 17255
rect 4488 17224 6469 17252
rect 4488 17212 4494 17224
rect 6457 17221 6469 17224
rect 6503 17221 6515 17255
rect 6457 17215 6515 17221
rect 7285 17255 7343 17261
rect 7285 17221 7297 17255
rect 7331 17252 7343 17255
rect 7650 17252 7656 17264
rect 7331 17224 7656 17252
rect 7331 17221 7343 17224
rect 7285 17215 7343 17221
rect 7650 17212 7656 17224
rect 7708 17212 7714 17264
rect 8110 17212 8116 17264
rect 8168 17252 8174 17264
rect 8168 17224 10088 17252
rect 8168 17212 8174 17224
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 1762 17184 1768 17196
rect 1719 17156 1768 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 2041 17187 2099 17193
rect 2041 17153 2053 17187
rect 2087 17153 2099 17187
rect 2041 17147 2099 17153
rect 2056 17116 2084 17147
rect 2130 17144 2136 17196
rect 2188 17184 2194 17196
rect 2317 17187 2375 17193
rect 2317 17184 2329 17187
rect 2188 17156 2329 17184
rect 2188 17144 2194 17156
rect 2317 17153 2329 17156
rect 2363 17153 2375 17187
rect 2317 17147 2375 17153
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17184 2835 17187
rect 3142 17184 3148 17196
rect 2823 17156 3148 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 3142 17144 3148 17156
rect 3200 17144 3206 17196
rect 3234 17144 3240 17196
rect 3292 17184 3298 17196
rect 3292 17156 3337 17184
rect 3292 17144 3298 17156
rect 4062 17144 4068 17196
rect 4120 17184 4126 17196
rect 4709 17187 4767 17193
rect 4709 17184 4721 17187
rect 4120 17156 4721 17184
rect 4120 17144 4126 17156
rect 4709 17153 4721 17156
rect 4755 17153 4767 17187
rect 5169 17187 5227 17193
rect 5169 17184 5181 17187
rect 4709 17147 4767 17153
rect 4816 17156 5181 17184
rect 2222 17116 2228 17128
rect 2056 17088 2228 17116
rect 2222 17076 2228 17088
rect 2280 17076 2286 17128
rect 2593 17119 2651 17125
rect 2593 17085 2605 17119
rect 2639 17116 2651 17119
rect 3050 17116 3056 17128
rect 2639 17088 3056 17116
rect 2639 17085 2651 17088
rect 2593 17079 2651 17085
rect 3050 17076 3056 17088
rect 3108 17076 3114 17128
rect 4816 16992 4844 17156
rect 5169 17153 5181 17156
rect 5215 17153 5227 17187
rect 5350 17184 5356 17196
rect 5311 17156 5356 17184
rect 5169 17147 5227 17153
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 5902 17184 5908 17196
rect 5859 17156 5908 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 5902 17144 5908 17156
rect 5960 17144 5966 17196
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17184 7251 17187
rect 7558 17184 7564 17196
rect 7239 17156 7564 17184
rect 7239 17153 7251 17156
rect 7193 17147 7251 17153
rect 7558 17144 7564 17156
rect 7616 17144 7622 17196
rect 7834 17144 7840 17196
rect 7892 17184 7898 17196
rect 8573 17187 8631 17193
rect 8573 17184 8585 17187
rect 7892 17156 8585 17184
rect 7892 17144 7898 17156
rect 8573 17153 8585 17156
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 8662 17144 8668 17196
rect 8720 17184 8726 17196
rect 9398 17184 9404 17196
rect 8720 17156 8765 17184
rect 9359 17156 9404 17184
rect 8720 17144 8726 17156
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 10060 17184 10088 17224
rect 10226 17212 10232 17264
rect 10284 17252 10290 17264
rect 12897 17255 12955 17261
rect 12897 17252 12909 17255
rect 10284 17224 12909 17252
rect 10284 17212 10290 17224
rect 12897 17221 12909 17224
rect 12943 17221 12955 17255
rect 12897 17215 12955 17221
rect 14093 17255 14151 17261
rect 14093 17221 14105 17255
rect 14139 17252 14151 17255
rect 15562 17252 15568 17264
rect 14139 17224 15568 17252
rect 14139 17221 14151 17224
rect 14093 17215 14151 17221
rect 15562 17212 15568 17224
rect 15620 17212 15626 17264
rect 19702 17212 19708 17264
rect 19760 17252 19766 17264
rect 20548 17252 20576 17280
rect 19760 17224 20576 17252
rect 19760 17212 19766 17224
rect 10117 17187 10175 17193
rect 10117 17184 10129 17187
rect 10060 17156 10129 17184
rect 10117 17153 10129 17156
rect 10163 17184 10175 17187
rect 11974 17184 11980 17196
rect 10163 17156 11980 17184
rect 10163 17153 10175 17156
rect 10117 17147 10175 17153
rect 11974 17144 11980 17156
rect 12032 17144 12038 17196
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17184 12219 17187
rect 13630 17184 13636 17196
rect 12207 17156 13636 17184
rect 12207 17153 12219 17156
rect 12161 17147 12219 17153
rect 5994 17116 6000 17128
rect 5955 17088 6000 17116
rect 5994 17076 6000 17088
rect 6052 17076 6058 17128
rect 7098 17116 7104 17128
rect 6564 17088 7104 17116
rect 4890 17008 4896 17060
rect 4948 17048 4954 17060
rect 4948 17020 5212 17048
rect 4948 17008 4954 17020
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 1854 16940 1860 16992
rect 1912 16980 1918 16992
rect 4798 16980 4804 16992
rect 1912 16952 4804 16980
rect 1912 16940 1918 16952
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 4985 16983 5043 16989
rect 4985 16949 4997 16983
rect 5031 16980 5043 16983
rect 5074 16980 5080 16992
rect 5031 16952 5080 16980
rect 5031 16949 5043 16952
rect 4985 16943 5043 16949
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 5184 16980 5212 17020
rect 5258 17008 5264 17060
rect 5316 17048 5322 17060
rect 6564 17048 6592 17088
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 7469 17119 7527 17125
rect 7469 17085 7481 17119
rect 7515 17116 7527 17119
rect 7650 17116 7656 17128
rect 7515 17088 7656 17116
rect 7515 17085 7527 17088
rect 7469 17079 7527 17085
rect 5316 17020 6592 17048
rect 6641 17051 6699 17057
rect 5316 17008 5322 17020
rect 6641 17017 6653 17051
rect 6687 17048 6699 17051
rect 6730 17048 6736 17060
rect 6687 17020 6736 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 6730 17008 6736 17020
rect 6788 17048 6794 17060
rect 7484 17048 7512 17079
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 7929 17119 7987 17125
rect 7929 17085 7941 17119
rect 7975 17116 7987 17119
rect 8680 17116 8708 17144
rect 7975 17088 8708 17116
rect 8849 17119 8907 17125
rect 7975 17085 7987 17088
rect 7929 17079 7987 17085
rect 8849 17085 8861 17119
rect 8895 17085 8907 17119
rect 8849 17079 8907 17085
rect 9585 17119 9643 17125
rect 9585 17085 9597 17119
rect 9631 17116 9643 17119
rect 9674 17116 9680 17128
rect 9631 17088 9680 17116
rect 9631 17085 9643 17088
rect 9585 17079 9643 17085
rect 8294 17048 8300 17060
rect 6788 17020 7512 17048
rect 7576 17020 8300 17048
rect 6788 17008 6794 17020
rect 7576 16980 7604 17020
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 8864 17048 8892 17079
rect 9600 17048 9628 17079
rect 9674 17076 9680 17088
rect 9732 17076 9738 17128
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 9861 17119 9919 17125
rect 9861 17116 9873 17119
rect 9824 17088 9873 17116
rect 9824 17076 9830 17088
rect 9861 17085 9873 17088
rect 9907 17085 9919 17119
rect 11609 17119 11667 17125
rect 11609 17116 11621 17119
rect 9861 17079 9919 17085
rect 10888 17088 11621 17116
rect 8864 17020 9628 17048
rect 5184 16952 7604 16980
rect 7834 16940 7840 16992
rect 7892 16980 7898 16992
rect 8021 16983 8079 16989
rect 8021 16980 8033 16983
rect 7892 16952 8033 16980
rect 7892 16940 7898 16952
rect 8021 16949 8033 16952
rect 8067 16949 8079 16983
rect 8021 16943 8079 16949
rect 10594 16940 10600 16992
rect 10652 16980 10658 16992
rect 10888 16980 10916 17088
rect 11609 17085 11621 17088
rect 11655 17116 11667 17119
rect 12176 17116 12204 17147
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 13725 17187 13783 17193
rect 13725 17153 13737 17187
rect 13771 17184 13783 17187
rect 14182 17184 14188 17196
rect 13771 17156 14188 17184
rect 13771 17153 13783 17156
rect 13725 17147 13783 17153
rect 14182 17144 14188 17156
rect 14240 17184 14246 17196
rect 14458 17184 14464 17196
rect 14240 17156 14464 17184
rect 14240 17144 14246 17156
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17184 15071 17187
rect 15838 17184 15844 17196
rect 15059 17156 15700 17184
rect 15799 17156 15844 17184
rect 15059 17153 15071 17156
rect 15013 17147 15071 17153
rect 11655 17088 12204 17116
rect 12253 17119 12311 17125
rect 11655 17085 11667 17088
rect 11609 17079 11667 17085
rect 12253 17085 12265 17119
rect 12299 17085 12311 17119
rect 12253 17079 12311 17085
rect 11238 17048 11244 17060
rect 11199 17020 11244 17048
rect 11238 17008 11244 17020
rect 11296 17048 11302 17060
rect 11698 17048 11704 17060
rect 11296 17020 11704 17048
rect 11296 17008 11302 17020
rect 11698 17008 11704 17020
rect 11756 17048 11762 17060
rect 12268 17048 12296 17079
rect 12526 17076 12532 17128
rect 12584 17116 12590 17128
rect 13081 17119 13139 17125
rect 13081 17116 13093 17119
rect 12584 17088 13093 17116
rect 12584 17076 12590 17088
rect 13081 17085 13093 17088
rect 13127 17085 13139 17119
rect 13081 17079 13139 17085
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13872 17088 13921 17116
rect 13872 17076 13878 17088
rect 13909 17085 13921 17088
rect 13955 17085 13967 17119
rect 15102 17116 15108 17128
rect 15063 17088 15108 17116
rect 13909 17079 13967 17085
rect 15102 17076 15108 17088
rect 15160 17076 15166 17128
rect 15194 17076 15200 17128
rect 15252 17116 15258 17128
rect 15565 17119 15623 17125
rect 15252 17088 15297 17116
rect 15252 17076 15258 17088
rect 15565 17085 15577 17119
rect 15611 17085 15623 17119
rect 15672 17116 15700 17156
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 19794 17184 19800 17196
rect 19755 17156 19800 17184
rect 19794 17144 19800 17156
rect 19852 17144 19858 17196
rect 20530 17184 20536 17196
rect 20491 17156 20536 17184
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 20806 17184 20812 17196
rect 20767 17156 20812 17184
rect 20806 17144 20812 17156
rect 20864 17144 20870 17196
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17153 21327 17187
rect 21269 17147 21327 17153
rect 16942 17116 16948 17128
rect 15672 17088 16948 17116
rect 15565 17079 15623 17085
rect 11756 17020 12296 17048
rect 11756 17008 11762 17020
rect 14366 17008 14372 17060
rect 14424 17048 14430 17060
rect 14553 17051 14611 17057
rect 14553 17048 14565 17051
rect 14424 17020 14565 17048
rect 14424 17008 14430 17020
rect 14553 17017 14565 17020
rect 14599 17017 14611 17051
rect 14553 17011 14611 17017
rect 15286 17008 15292 17060
rect 15344 17048 15350 17060
rect 15580 17048 15608 17079
rect 16942 17076 16948 17088
rect 17000 17076 17006 17128
rect 20438 17076 20444 17128
rect 20496 17116 20502 17128
rect 21284 17116 21312 17147
rect 20496 17088 21312 17116
rect 20496 17076 20502 17088
rect 20622 17048 20628 17060
rect 15344 17020 15608 17048
rect 15672 17020 20628 17048
rect 15344 17008 15350 17020
rect 10652 16952 10916 16980
rect 10652 16940 10658 16952
rect 11974 16940 11980 16992
rect 12032 16980 12038 16992
rect 12158 16980 12164 16992
rect 12032 16952 12164 16980
rect 12032 16940 12038 16952
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 12529 16983 12587 16989
rect 12529 16949 12541 16983
rect 12575 16980 12587 16983
rect 12618 16980 12624 16992
rect 12575 16952 12624 16980
rect 12575 16949 12587 16952
rect 12529 16943 12587 16949
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 13354 16940 13360 16992
rect 13412 16980 13418 16992
rect 13541 16983 13599 16989
rect 13541 16980 13553 16983
rect 13412 16952 13553 16980
rect 13412 16940 13418 16952
rect 13541 16949 13553 16952
rect 13587 16949 13599 16983
rect 13541 16943 13599 16949
rect 13722 16940 13728 16992
rect 13780 16980 13786 16992
rect 15672 16980 15700 17020
rect 20622 17008 20628 17020
rect 20680 17008 20686 17060
rect 20806 17008 20812 17060
rect 20864 17048 20870 17060
rect 21177 17051 21235 17057
rect 21177 17048 21189 17051
rect 20864 17020 21189 17048
rect 20864 17008 20870 17020
rect 21177 17017 21189 17020
rect 21223 17048 21235 17051
rect 22830 17048 22836 17060
rect 21223 17020 22836 17048
rect 21223 17017 21235 17020
rect 21177 17011 21235 17017
rect 22830 17008 22836 17020
rect 22888 17008 22894 17060
rect 13780 16952 15700 16980
rect 13780 16940 13786 16952
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 16209 16983 16267 16989
rect 16209 16980 16221 16983
rect 16080 16952 16221 16980
rect 16080 16940 16086 16952
rect 16209 16949 16221 16952
rect 16255 16949 16267 16983
rect 16209 16943 16267 16949
rect 19886 16940 19892 16992
rect 19944 16980 19950 16992
rect 20349 16983 20407 16989
rect 20349 16980 20361 16983
rect 19944 16952 20361 16980
rect 19944 16940 19950 16952
rect 20349 16949 20361 16952
rect 20395 16980 20407 16983
rect 20530 16980 20536 16992
rect 20395 16952 20536 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 21450 16980 21456 16992
rect 21411 16952 21456 16980
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 2133 16779 2191 16785
rect 2133 16776 2145 16779
rect 1728 16748 2145 16776
rect 1728 16736 1734 16748
rect 2133 16745 2145 16748
rect 2179 16745 2191 16779
rect 2133 16739 2191 16745
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 4522 16776 4528 16788
rect 2832 16748 2877 16776
rect 4172 16748 4528 16776
rect 2832 16736 2838 16748
rect 2498 16668 2504 16720
rect 2556 16708 2562 16720
rect 4172 16708 4200 16748
rect 4522 16736 4528 16748
rect 4580 16736 4586 16788
rect 4798 16736 4804 16788
rect 4856 16776 4862 16788
rect 5629 16779 5687 16785
rect 5629 16776 5641 16779
rect 4856 16748 5641 16776
rect 4856 16736 4862 16748
rect 5629 16745 5641 16748
rect 5675 16745 5687 16779
rect 6638 16776 6644 16788
rect 6599 16748 6644 16776
rect 5629 16739 5687 16745
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 7248 16748 7665 16776
rect 7248 16736 7254 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 7653 16739 7711 16745
rect 7742 16736 7748 16788
rect 7800 16776 7806 16788
rect 7837 16779 7895 16785
rect 7837 16776 7849 16779
rect 7800 16748 7849 16776
rect 7800 16736 7806 16748
rect 7837 16745 7849 16748
rect 7883 16745 7895 16779
rect 7837 16739 7895 16745
rect 8386 16736 8392 16788
rect 8444 16776 8450 16788
rect 8757 16779 8815 16785
rect 8757 16776 8769 16779
rect 8444 16748 8769 16776
rect 8444 16736 8450 16748
rect 8757 16745 8769 16748
rect 8803 16745 8815 16779
rect 8757 16739 8815 16745
rect 9674 16736 9680 16788
rect 9732 16736 9738 16788
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 12342 16776 12348 16788
rect 11112 16748 12348 16776
rect 11112 16736 11118 16748
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 14458 16776 14464 16788
rect 14108 16748 14464 16776
rect 2556 16680 4200 16708
rect 5537 16711 5595 16717
rect 2556 16668 2562 16680
rect 5537 16677 5549 16711
rect 5583 16677 5595 16711
rect 9692 16708 9720 16736
rect 5537 16671 5595 16677
rect 7116 16680 7604 16708
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2924 16612 2973 16640
rect 2924 16600 2930 16612
rect 2961 16609 2973 16612
rect 3007 16609 3019 16643
rect 2961 16603 3019 16609
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16640 3203 16643
rect 5552 16640 5580 16671
rect 5626 16640 5632 16652
rect 3191 16612 4108 16640
rect 5539 16612 5632 16640
rect 3191 16609 3203 16612
rect 3145 16603 3203 16609
rect 1670 16572 1676 16584
rect 1631 16544 1676 16572
rect 1670 16532 1676 16544
rect 1728 16532 1734 16584
rect 2041 16575 2099 16581
rect 2041 16541 2053 16575
rect 2087 16572 2099 16575
rect 2222 16572 2228 16584
rect 2087 16544 2228 16572
rect 2087 16541 2099 16544
rect 2041 16535 2099 16541
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 2317 16575 2375 16581
rect 2317 16541 2329 16575
rect 2363 16572 2375 16575
rect 2363 16544 2544 16572
rect 2363 16541 2375 16544
rect 2317 16535 2375 16541
rect 2516 16516 2544 16544
rect 2590 16532 2596 16584
rect 2648 16572 2654 16584
rect 3970 16572 3976 16584
rect 2648 16544 2693 16572
rect 2976 16544 3976 16572
rect 2648 16532 2654 16544
rect 2976 16516 3004 16544
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 1394 16464 1400 16516
rect 1452 16504 1458 16516
rect 1452 16476 2452 16504
rect 1452 16464 1458 16476
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 1854 16436 1860 16448
rect 1815 16408 1860 16436
rect 1854 16396 1860 16408
rect 1912 16396 1918 16448
rect 2424 16445 2452 16476
rect 2498 16464 2504 16516
rect 2556 16464 2562 16516
rect 2958 16464 2964 16516
rect 3016 16464 3022 16516
rect 3237 16507 3295 16513
rect 3237 16473 3249 16507
rect 3283 16504 3295 16507
rect 3789 16507 3847 16513
rect 3789 16504 3801 16507
rect 3283 16476 3801 16504
rect 3283 16473 3295 16476
rect 3237 16467 3295 16473
rect 3789 16473 3801 16476
rect 3835 16473 3847 16507
rect 4080 16504 4108 16612
rect 5626 16600 5632 16612
rect 5684 16640 5690 16652
rect 6457 16643 6515 16649
rect 6457 16640 6469 16643
rect 5684 16612 6469 16640
rect 5684 16600 5690 16612
rect 6457 16609 6469 16612
rect 6503 16640 6515 16643
rect 6546 16640 6552 16652
rect 6503 16612 6552 16640
rect 6503 16609 6515 16612
rect 6457 16603 6515 16609
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 7116 16649 7144 16680
rect 7576 16652 7604 16680
rect 8128 16680 9720 16708
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16609 7159 16643
rect 7101 16603 7159 16609
rect 7285 16643 7343 16649
rect 7285 16609 7297 16643
rect 7331 16609 7343 16643
rect 7558 16640 7564 16652
rect 7519 16612 7564 16640
rect 7285 16603 7343 16609
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16572 4215 16575
rect 4246 16572 4252 16584
rect 4203 16544 4252 16572
rect 4203 16541 4215 16544
rect 4157 16535 4215 16541
rect 4246 16532 4252 16544
rect 4304 16532 4310 16584
rect 4430 16581 4436 16584
rect 4424 16572 4436 16581
rect 4391 16544 4436 16572
rect 4424 16535 4436 16544
rect 4430 16532 4436 16535
rect 4488 16532 4494 16584
rect 4706 16532 4712 16584
rect 4764 16572 4770 16584
rect 4764 16544 6132 16572
rect 4764 16532 4770 16544
rect 4264 16504 4292 16532
rect 4982 16504 4988 16516
rect 4080 16476 4200 16504
rect 4264 16476 4988 16504
rect 3789 16467 3847 16473
rect 2409 16439 2467 16445
rect 2409 16405 2421 16439
rect 2455 16405 2467 16439
rect 2409 16399 2467 16405
rect 3326 16396 3332 16448
rect 3384 16436 3390 16448
rect 3605 16439 3663 16445
rect 3605 16436 3617 16439
rect 3384 16408 3617 16436
rect 3384 16396 3390 16408
rect 3605 16405 3617 16408
rect 3651 16405 3663 16439
rect 4172 16436 4200 16476
rect 4982 16464 4988 16476
rect 5040 16464 5046 16516
rect 6104 16504 6132 16544
rect 6178 16532 6184 16584
rect 6236 16572 6242 16584
rect 7300 16572 7328 16603
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 8128 16649 8156 16680
rect 10410 16668 10416 16720
rect 10468 16708 10474 16720
rect 12434 16708 12440 16720
rect 10468 16680 12440 16708
rect 10468 16668 10474 16680
rect 12434 16668 12440 16680
rect 12492 16668 12498 16720
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16609 8171 16643
rect 8113 16603 8171 16609
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 9030 16640 9036 16652
rect 8628 16612 9036 16640
rect 8628 16600 8634 16612
rect 9030 16600 9036 16612
rect 9088 16640 9094 16652
rect 9309 16643 9367 16649
rect 9309 16640 9321 16643
rect 9088 16612 9321 16640
rect 9088 16600 9094 16612
rect 9309 16609 9321 16612
rect 9355 16640 9367 16643
rect 9398 16640 9404 16652
rect 9355 16612 9404 16640
rect 9355 16609 9367 16612
rect 9309 16603 9367 16609
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 10870 16640 10876 16652
rect 10831 16612 10876 16640
rect 10870 16600 10876 16612
rect 10928 16600 10934 16652
rect 11698 16640 11704 16652
rect 11659 16612 11704 16640
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 14108 16649 14136 16748
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 15562 16776 15568 16788
rect 15523 16748 15568 16776
rect 15562 16736 15568 16748
rect 15620 16736 15626 16788
rect 15838 16736 15844 16788
rect 15896 16776 15902 16788
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 15896 16748 16405 16776
rect 15896 16736 15902 16748
rect 16393 16745 16405 16748
rect 16439 16745 16451 16779
rect 16393 16739 16451 16745
rect 16482 16736 16488 16788
rect 16540 16776 16546 16788
rect 18417 16779 18475 16785
rect 18417 16776 18429 16779
rect 16540 16748 18429 16776
rect 16540 16736 16546 16748
rect 18417 16745 18429 16748
rect 18463 16776 18475 16779
rect 18782 16776 18788 16788
rect 18463 16748 18788 16776
rect 18463 16745 18475 16748
rect 18417 16739 18475 16745
rect 18782 16736 18788 16748
rect 18840 16736 18846 16788
rect 19429 16779 19487 16785
rect 19429 16745 19441 16779
rect 19475 16776 19487 16779
rect 19794 16776 19800 16788
rect 19475 16748 19800 16776
rect 19475 16745 19487 16748
rect 19429 16739 19487 16745
rect 19794 16736 19800 16748
rect 19852 16736 19858 16788
rect 20809 16779 20867 16785
rect 20809 16745 20821 16779
rect 20855 16776 20867 16779
rect 21266 16776 21272 16788
rect 20855 16748 21272 16776
rect 20855 16745 20867 16748
rect 20809 16739 20867 16745
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 18230 16708 18236 16720
rect 17052 16680 18236 16708
rect 13909 16643 13967 16649
rect 13909 16640 13921 16643
rect 13832 16612 13921 16640
rect 7650 16572 7656 16584
rect 6236 16544 6281 16572
rect 7300 16544 7656 16572
rect 6236 16532 6242 16544
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 10042 16572 10048 16584
rect 8312 16544 10048 16572
rect 8312 16504 8340 16544
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 13354 16532 13360 16584
rect 13412 16572 13418 16584
rect 13832 16572 13860 16612
rect 13909 16609 13921 16612
rect 13955 16609 13967 16643
rect 13909 16603 13967 16609
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16609 14151 16643
rect 16022 16640 16028 16652
rect 15983 16612 16028 16640
rect 14093 16603 14151 16609
rect 16022 16600 16028 16612
rect 16080 16600 16086 16652
rect 16117 16643 16175 16649
rect 16117 16609 16129 16643
rect 16163 16609 16175 16643
rect 16117 16603 16175 16609
rect 13412 16544 13860 16572
rect 13412 16532 13418 16544
rect 6104 16476 8340 16504
rect 8389 16507 8447 16513
rect 8389 16473 8401 16507
rect 8435 16504 8447 16507
rect 8941 16507 8999 16513
rect 8941 16504 8953 16507
rect 8435 16476 8953 16504
rect 8435 16473 8447 16476
rect 8389 16467 8447 16473
rect 8941 16473 8953 16476
rect 8987 16473 8999 16507
rect 10781 16507 10839 16513
rect 10781 16504 10793 16507
rect 8941 16467 8999 16473
rect 10244 16476 10793 16504
rect 4430 16436 4436 16448
rect 4172 16408 4436 16436
rect 3605 16399 3663 16405
rect 4430 16396 4436 16408
rect 4488 16396 4494 16448
rect 5810 16436 5816 16448
rect 5771 16408 5816 16436
rect 5810 16396 5816 16408
rect 5868 16396 5874 16448
rect 6273 16439 6331 16445
rect 6273 16405 6285 16439
rect 6319 16436 6331 16439
rect 6822 16436 6828 16448
rect 6319 16408 6828 16436
rect 6319 16405 6331 16408
rect 6273 16399 6331 16405
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 7006 16436 7012 16448
rect 6967 16408 7012 16436
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 7190 16396 7196 16448
rect 7248 16436 7254 16448
rect 7374 16436 7380 16448
rect 7248 16408 7380 16436
rect 7248 16396 7254 16408
rect 7374 16396 7380 16408
rect 7432 16396 7438 16448
rect 8294 16436 8300 16448
rect 8255 16408 8300 16436
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 8570 16396 8576 16448
rect 8628 16436 8634 16448
rect 9306 16436 9312 16448
rect 8628 16408 9312 16436
rect 8628 16396 8634 16408
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 9582 16396 9588 16448
rect 9640 16436 9646 16448
rect 9769 16439 9827 16445
rect 9769 16436 9781 16439
rect 9640 16408 9781 16436
rect 9640 16396 9646 16408
rect 9769 16405 9781 16408
rect 9815 16405 9827 16439
rect 9769 16399 9827 16405
rect 9858 16396 9864 16448
rect 9916 16436 9922 16448
rect 10244 16445 10272 16476
rect 10781 16473 10793 16476
rect 10827 16473 10839 16507
rect 10781 16467 10839 16473
rect 11238 16464 11244 16516
rect 11296 16504 11302 16516
rect 11609 16507 11667 16513
rect 11609 16504 11621 16507
rect 11296 16476 11621 16504
rect 11296 16464 11302 16476
rect 11609 16473 11621 16476
rect 11655 16473 11667 16507
rect 11609 16467 11667 16473
rect 13664 16507 13722 16513
rect 13664 16473 13676 16507
rect 13710 16504 13722 16507
rect 14360 16507 14418 16513
rect 13710 16476 14320 16504
rect 13710 16473 13722 16476
rect 13664 16467 13722 16473
rect 10229 16439 10287 16445
rect 9916 16408 9961 16436
rect 9916 16396 9922 16408
rect 10229 16405 10241 16439
rect 10275 16405 10287 16439
rect 10229 16399 10287 16405
rect 10318 16396 10324 16448
rect 10376 16436 10382 16448
rect 10686 16436 10692 16448
rect 10376 16408 10421 16436
rect 10647 16408 10692 16436
rect 10376 16396 10382 16408
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 11149 16439 11207 16445
rect 11149 16436 11161 16439
rect 11020 16408 11161 16436
rect 11020 16396 11026 16408
rect 11149 16405 11161 16408
rect 11195 16405 11207 16439
rect 11149 16399 11207 16405
rect 11517 16439 11575 16445
rect 11517 16405 11529 16439
rect 11563 16436 11575 16439
rect 12069 16439 12127 16445
rect 12069 16436 12081 16439
rect 11563 16408 12081 16436
rect 11563 16405 11575 16408
rect 11517 16399 11575 16405
rect 12069 16405 12081 16408
rect 12115 16436 12127 16439
rect 12342 16436 12348 16448
rect 12115 16408 12348 16436
rect 12115 16405 12127 16408
rect 12069 16399 12127 16405
rect 12342 16396 12348 16408
rect 12400 16396 12406 16448
rect 12529 16439 12587 16445
rect 12529 16405 12541 16439
rect 12575 16436 12587 16439
rect 13814 16436 13820 16448
rect 12575 16408 13820 16436
rect 12575 16405 12587 16408
rect 12529 16399 12587 16405
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 14292 16436 14320 16476
rect 14360 16473 14372 16507
rect 14406 16504 14418 16507
rect 15286 16504 15292 16516
rect 14406 16476 15292 16504
rect 14406 16473 14418 16476
rect 14360 16467 14418 16473
rect 15286 16464 15292 16476
rect 15344 16464 15350 16516
rect 16132 16504 16160 16603
rect 16298 16600 16304 16652
rect 16356 16640 16362 16652
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 16356 16612 16957 16640
rect 16356 16600 16362 16612
rect 16945 16609 16957 16612
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 17052 16572 17080 16680
rect 18230 16668 18236 16680
rect 18288 16668 18294 16720
rect 17310 16640 17316 16652
rect 17271 16612 17316 16640
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 17494 16640 17500 16652
rect 17455 16612 17500 16640
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 18049 16643 18107 16649
rect 18049 16609 18061 16643
rect 18095 16640 18107 16643
rect 20162 16640 20168 16652
rect 18095 16612 20168 16640
rect 18095 16609 18107 16612
rect 18049 16603 18107 16609
rect 18064 16572 18092 16603
rect 20162 16600 20168 16612
rect 20220 16600 20226 16652
rect 16899 16544 17080 16572
rect 17144 16544 18092 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 15488 16476 16160 16504
rect 15194 16436 15200 16448
rect 14292 16408 15200 16436
rect 15194 16396 15200 16408
rect 15252 16436 15258 16448
rect 15488 16445 15516 16476
rect 16390 16464 16396 16516
rect 16448 16504 16454 16516
rect 16761 16507 16819 16513
rect 16761 16504 16773 16507
rect 16448 16476 16773 16504
rect 16448 16464 16454 16476
rect 16761 16473 16773 16476
rect 16807 16504 16819 16507
rect 17144 16504 17172 16544
rect 18138 16532 18144 16584
rect 18196 16572 18202 16584
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 18196 16544 19257 16572
rect 18196 16532 18202 16544
rect 19245 16541 19257 16544
rect 19291 16541 19303 16575
rect 20625 16575 20683 16581
rect 20625 16572 20637 16575
rect 19245 16535 19303 16541
rect 20456 16544 20637 16572
rect 20070 16504 20076 16516
rect 16807 16476 17172 16504
rect 17972 16476 20076 16504
rect 16807 16473 16819 16476
rect 16761 16467 16819 16473
rect 15473 16439 15531 16445
rect 15473 16436 15485 16439
rect 15252 16408 15485 16436
rect 15252 16396 15258 16408
rect 15473 16405 15485 16408
rect 15519 16405 15531 16439
rect 15473 16399 15531 16405
rect 15838 16396 15844 16448
rect 15896 16436 15902 16448
rect 15933 16439 15991 16445
rect 15933 16436 15945 16439
rect 15896 16408 15945 16436
rect 15896 16396 15902 16408
rect 15933 16405 15945 16408
rect 15979 16405 15991 16439
rect 15933 16399 15991 16405
rect 17586 16396 17592 16448
rect 17644 16436 17650 16448
rect 17972 16445 18000 16476
rect 20070 16464 20076 16476
rect 20128 16464 20134 16516
rect 17957 16439 18015 16445
rect 17644 16408 17689 16436
rect 17644 16396 17650 16408
rect 17957 16405 17969 16439
rect 18003 16405 18015 16439
rect 17957 16399 18015 16405
rect 18506 16396 18512 16448
rect 18564 16436 18570 16448
rect 18601 16439 18659 16445
rect 18601 16436 18613 16439
rect 18564 16408 18613 16436
rect 18564 16396 18570 16408
rect 18601 16405 18613 16408
rect 18647 16405 18659 16439
rect 18601 16399 18659 16405
rect 19978 16396 19984 16448
rect 20036 16436 20042 16448
rect 20456 16445 20484 16544
rect 20625 16541 20637 16544
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 20901 16575 20959 16581
rect 20901 16541 20913 16575
rect 20947 16572 20959 16575
rect 20990 16572 20996 16584
rect 20947 16544 20996 16572
rect 20947 16541 20959 16544
rect 20901 16535 20959 16541
rect 20990 16532 20996 16544
rect 21048 16532 21054 16584
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16541 21327 16575
rect 21269 16535 21327 16541
rect 20714 16464 20720 16516
rect 20772 16504 20778 16516
rect 21284 16504 21312 16535
rect 20772 16476 21312 16504
rect 20772 16464 20778 16476
rect 20441 16439 20499 16445
rect 20441 16436 20453 16439
rect 20036 16408 20453 16436
rect 20036 16396 20042 16408
rect 20441 16405 20453 16408
rect 20487 16405 20499 16439
rect 21082 16436 21088 16448
rect 21043 16408 21088 16436
rect 20441 16399 20499 16405
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 21450 16436 21456 16448
rect 21411 16408 21456 16436
rect 21450 16396 21456 16408
rect 21508 16396 21514 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 1670 16192 1676 16244
rect 1728 16232 1734 16244
rect 1857 16235 1915 16241
rect 1857 16232 1869 16235
rect 1728 16204 1869 16232
rect 1728 16192 1734 16204
rect 1857 16201 1869 16204
rect 1903 16201 1915 16235
rect 2314 16232 2320 16244
rect 2275 16204 2320 16232
rect 1857 16195 1915 16201
rect 2314 16192 2320 16204
rect 2372 16192 2378 16244
rect 2406 16192 2412 16244
rect 2464 16232 2470 16244
rect 2685 16235 2743 16241
rect 2685 16232 2697 16235
rect 2464 16204 2697 16232
rect 2464 16192 2470 16204
rect 2685 16201 2697 16204
rect 2731 16201 2743 16235
rect 3326 16232 3332 16244
rect 3287 16204 3332 16232
rect 2685 16195 2743 16201
rect 3326 16192 3332 16204
rect 3384 16192 3390 16244
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 3878 16232 3884 16244
rect 3743 16204 3884 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 3878 16192 3884 16204
rect 3936 16192 3942 16244
rect 4157 16235 4215 16241
rect 4157 16201 4169 16235
rect 4203 16232 4215 16235
rect 4617 16235 4675 16241
rect 4617 16232 4629 16235
rect 4203 16204 4629 16232
rect 4203 16201 4215 16204
rect 4157 16195 4215 16201
rect 4617 16201 4629 16204
rect 4663 16201 4675 16235
rect 4617 16195 4675 16201
rect 5902 16192 5908 16244
rect 5960 16232 5966 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 5960 16204 6193 16232
rect 5960 16192 5966 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 6181 16195 6239 16201
rect 6822 16192 6828 16244
rect 6880 16232 6886 16244
rect 7101 16235 7159 16241
rect 7101 16232 7113 16235
rect 6880 16204 7113 16232
rect 6880 16192 6886 16204
rect 7101 16201 7113 16204
rect 7147 16201 7159 16235
rect 7101 16195 7159 16201
rect 8018 16192 8024 16244
rect 8076 16232 8082 16244
rect 8665 16235 8723 16241
rect 8665 16232 8677 16235
rect 8076 16204 8677 16232
rect 8076 16192 8082 16204
rect 8665 16201 8677 16204
rect 8711 16201 8723 16235
rect 8665 16195 8723 16201
rect 8941 16235 8999 16241
rect 8941 16201 8953 16235
rect 8987 16232 8999 16235
rect 9122 16232 9128 16244
rect 8987 16204 9128 16232
rect 8987 16201 8999 16204
rect 8941 16195 8999 16201
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 9306 16192 9312 16244
rect 9364 16232 9370 16244
rect 10226 16232 10232 16244
rect 9364 16204 10232 16232
rect 9364 16192 9370 16204
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 10781 16235 10839 16241
rect 10781 16201 10793 16235
rect 10827 16232 10839 16235
rect 10870 16232 10876 16244
rect 10827 16204 10876 16232
rect 10827 16201 10839 16204
rect 10781 16195 10839 16201
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 11790 16192 11796 16244
rect 11848 16232 11854 16244
rect 13449 16235 13507 16241
rect 13449 16232 13461 16235
rect 11848 16204 13461 16232
rect 11848 16192 11854 16204
rect 13449 16201 13461 16204
rect 13495 16201 13507 16235
rect 13449 16195 13507 16201
rect 13814 16192 13820 16244
rect 13872 16192 13878 16244
rect 15013 16235 15071 16241
rect 15013 16201 15025 16235
rect 15059 16232 15071 16235
rect 15102 16232 15108 16244
rect 15059 16204 15108 16232
rect 15059 16201 15071 16204
rect 15013 16195 15071 16201
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 15381 16235 15439 16241
rect 15381 16201 15393 16235
rect 15427 16232 15439 16235
rect 15654 16232 15660 16244
rect 15427 16204 15660 16232
rect 15427 16201 15439 16204
rect 15381 16195 15439 16201
rect 15654 16192 15660 16204
rect 15712 16192 15718 16244
rect 15838 16232 15844 16244
rect 15799 16204 15844 16232
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 16298 16192 16304 16244
rect 16356 16232 16362 16244
rect 16393 16235 16451 16241
rect 16393 16232 16405 16235
rect 16356 16204 16405 16232
rect 16356 16192 16362 16204
rect 16393 16201 16405 16204
rect 16439 16201 16451 16235
rect 16393 16195 16451 16201
rect 16669 16235 16727 16241
rect 16669 16201 16681 16235
rect 16715 16232 16727 16235
rect 16942 16232 16948 16244
rect 16715 16204 16948 16232
rect 16715 16201 16727 16204
rect 16669 16195 16727 16201
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 17497 16235 17555 16241
rect 17497 16201 17509 16235
rect 17543 16232 17555 16235
rect 17586 16232 17592 16244
rect 17543 16204 17592 16232
rect 17543 16201 17555 16204
rect 17497 16195 17555 16201
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 17957 16235 18015 16241
rect 17957 16201 17969 16235
rect 18003 16232 18015 16235
rect 18325 16235 18383 16241
rect 18325 16232 18337 16235
rect 18003 16204 18337 16232
rect 18003 16201 18015 16204
rect 17957 16195 18015 16201
rect 18325 16201 18337 16204
rect 18371 16201 18383 16235
rect 18782 16232 18788 16244
rect 18743 16204 18788 16232
rect 18325 16195 18383 16201
rect 18782 16192 18788 16204
rect 18840 16192 18846 16244
rect 20438 16232 20444 16244
rect 20399 16204 20444 16232
rect 20438 16192 20444 16204
rect 20496 16192 20502 16244
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 20990 16232 20996 16244
rect 20951 16204 20996 16232
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 106 16124 112 16176
rect 164 16164 170 16176
rect 164 16136 2912 16164
rect 164 16124 170 16136
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 1946 16096 1952 16108
rect 1719 16068 1952 16096
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 1946 16056 1952 16068
rect 2004 16056 2010 16108
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16065 2191 16099
rect 2133 16059 2191 16065
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16096 2559 16099
rect 2682 16096 2688 16108
rect 2547 16068 2688 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 1854 15988 1860 16040
rect 1912 16028 1918 16040
rect 2056 16028 2084 16059
rect 1912 16000 2084 16028
rect 1912 15988 1918 16000
rect 2038 15920 2044 15972
rect 2096 15960 2102 15972
rect 2148 15960 2176 16059
rect 2682 16056 2688 16068
rect 2740 16056 2746 16108
rect 2096 15932 2176 15960
rect 2096 15920 2102 15932
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 2148 15892 2176 15932
rect 2774 15892 2780 15904
rect 2148 15864 2780 15892
rect 2774 15852 2780 15864
rect 2832 15852 2838 15904
rect 2884 15901 2912 16136
rect 3970 16124 3976 16176
rect 4028 16164 4034 16176
rect 5721 16167 5779 16173
rect 5721 16164 5733 16167
rect 4028 16136 5733 16164
rect 4028 16124 4034 16136
rect 5721 16133 5733 16136
rect 5767 16133 5779 16167
rect 5721 16127 5779 16133
rect 5994 16124 6000 16176
rect 6052 16164 6058 16176
rect 6641 16167 6699 16173
rect 6641 16164 6653 16167
rect 6052 16136 6653 16164
rect 6052 16124 6058 16136
rect 6641 16133 6653 16136
rect 6687 16164 6699 16167
rect 7006 16164 7012 16176
rect 6687 16136 7012 16164
rect 6687 16133 6699 16136
rect 6641 16127 6699 16133
rect 7006 16124 7012 16136
rect 7064 16124 7070 16176
rect 9030 16164 9036 16176
rect 7116 16136 8708 16164
rect 8991 16136 9036 16164
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16096 4307 16099
rect 4706 16096 4712 16108
rect 4295 16068 4712 16096
rect 4295 16065 4307 16068
rect 4249 16059 4307 16065
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 4985 16099 5043 16105
rect 4985 16065 4997 16099
rect 5031 16096 5043 16099
rect 5350 16096 5356 16108
rect 5031 16068 5356 16096
rect 5031 16065 5043 16068
rect 4985 16059 5043 16065
rect 5350 16056 5356 16068
rect 5408 16096 5414 16108
rect 5813 16099 5871 16105
rect 5408 16068 5764 16096
rect 5408 16056 5414 16068
rect 3050 16028 3056 16040
rect 3011 16000 3056 16028
rect 3050 15988 3056 16000
rect 3108 15988 3114 16040
rect 3234 16028 3240 16040
rect 3195 16000 3240 16028
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 4062 15988 4068 16040
rect 4120 16028 4126 16040
rect 4341 16031 4399 16037
rect 4341 16028 4353 16031
rect 4120 16000 4353 16028
rect 4120 15988 4126 16000
rect 4341 15997 4353 16000
rect 4387 15997 4399 16031
rect 5074 16028 5080 16040
rect 5035 16000 5080 16028
rect 4341 15991 4399 15997
rect 5074 15988 5080 16000
rect 5132 15988 5138 16040
rect 5261 16031 5319 16037
rect 5261 15997 5273 16031
rect 5307 16028 5319 16031
rect 5442 16028 5448 16040
rect 5307 16000 5448 16028
rect 5307 15997 5319 16000
rect 5261 15991 5319 15997
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 5626 16028 5632 16040
rect 5587 16000 5632 16028
rect 5626 15988 5632 16000
rect 5684 15988 5690 16040
rect 5736 16028 5764 16068
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6365 16099 6423 16105
rect 6365 16096 6377 16099
rect 5859 16068 6377 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 6365 16065 6377 16068
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 7116 16028 7144 16136
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16096 7527 16099
rect 8113 16099 8171 16105
rect 8113 16096 8125 16099
rect 7515 16068 8125 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 8113 16065 8125 16068
rect 8159 16065 8171 16099
rect 8113 16059 8171 16065
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16065 8631 16099
rect 8680 16096 8708 16136
rect 9030 16124 9036 16136
rect 9088 16124 9094 16176
rect 11422 16164 11428 16176
rect 9140 16136 11428 16164
rect 9140 16096 9168 16136
rect 11422 16124 11428 16136
rect 11480 16164 11486 16176
rect 11882 16164 11888 16176
rect 11480 16136 11888 16164
rect 11480 16124 11486 16136
rect 11882 16124 11888 16136
rect 11940 16124 11946 16176
rect 13112 16167 13170 16173
rect 13112 16133 13124 16167
rect 13158 16164 13170 16167
rect 13832 16164 13860 16192
rect 13158 16136 13860 16164
rect 13158 16133 13170 16136
rect 13112 16127 13170 16133
rect 14366 16124 14372 16176
rect 14424 16164 14430 16176
rect 14645 16167 14703 16173
rect 14645 16164 14657 16167
rect 14424 16136 14657 16164
rect 14424 16124 14430 16136
rect 14645 16133 14657 16136
rect 14691 16133 14703 16167
rect 14645 16127 14703 16133
rect 18506 16124 18512 16176
rect 18564 16164 18570 16176
rect 18693 16167 18751 16173
rect 18693 16164 18705 16167
rect 18564 16136 18705 16164
rect 18564 16124 18570 16136
rect 18693 16133 18705 16136
rect 18739 16133 18751 16167
rect 21085 16167 21143 16173
rect 21085 16164 21097 16167
rect 18693 16127 18751 16133
rect 20548 16136 21097 16164
rect 20548 16108 20576 16136
rect 21085 16133 21097 16136
rect 21131 16133 21143 16167
rect 21085 16127 21143 16133
rect 8680 16068 9168 16096
rect 8573 16059 8631 16065
rect 5736 16000 7144 16028
rect 3142 15920 3148 15972
rect 3200 15960 3206 15972
rect 3789 15963 3847 15969
rect 3789 15960 3801 15963
rect 3200 15932 3801 15960
rect 3200 15920 3206 15932
rect 3789 15929 3801 15932
rect 3835 15929 3847 15963
rect 3789 15923 3847 15929
rect 3878 15920 3884 15972
rect 3936 15960 3942 15972
rect 7484 15960 7512 16059
rect 7561 16031 7619 16037
rect 7561 15997 7573 16031
rect 7607 15997 7619 16031
rect 7561 15991 7619 15997
rect 3936 15932 7512 15960
rect 7576 15960 7604 15991
rect 7650 15988 7656 16040
rect 7708 16028 7714 16040
rect 8588 16028 8616 16059
rect 9306 16056 9312 16108
rect 9364 16096 9370 16108
rect 9674 16105 9680 16108
rect 9657 16099 9680 16105
rect 9657 16096 9669 16099
rect 9364 16068 9669 16096
rect 9364 16056 9370 16068
rect 9657 16065 9669 16068
rect 9732 16096 9738 16108
rect 9732 16068 9805 16096
rect 9657 16059 9680 16065
rect 9674 16056 9680 16059
rect 9732 16056 9738 16068
rect 10502 16056 10508 16108
rect 10560 16096 10566 16108
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 10560 16068 11069 16096
rect 10560 16056 10566 16068
rect 11057 16065 11069 16068
rect 11103 16096 11115 16099
rect 13354 16096 13360 16108
rect 11103 16068 13360 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 13354 16056 13360 16068
rect 13412 16056 13418 16108
rect 13817 16099 13875 16105
rect 13817 16065 13829 16099
rect 13863 16096 13875 16099
rect 13863 16068 14228 16096
rect 13863 16065 13875 16068
rect 13817 16059 13875 16065
rect 9401 16031 9459 16037
rect 9401 16028 9413 16031
rect 7708 16000 7753 16028
rect 8588 16000 9413 16028
rect 7708 15988 7714 16000
rect 9401 15997 9413 16000
rect 9447 15997 9459 16031
rect 9401 15991 9459 15997
rect 8018 15960 8024 15972
rect 7576 15932 8024 15960
rect 3936 15920 3942 15932
rect 8018 15920 8024 15932
rect 8076 15920 8082 15972
rect 2869 15895 2927 15901
rect 2869 15861 2881 15895
rect 2915 15892 2927 15895
rect 3050 15892 3056 15904
rect 2915 15864 3056 15892
rect 2915 15861 2927 15864
rect 2869 15855 2927 15861
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 6822 15852 6828 15904
rect 6880 15892 6886 15904
rect 6917 15895 6975 15901
rect 6917 15892 6929 15895
rect 6880 15864 6929 15892
rect 6880 15852 6886 15864
rect 6917 15861 6929 15864
rect 6963 15892 6975 15895
rect 7742 15892 7748 15904
rect 6963 15864 7748 15892
rect 6963 15861 6975 15864
rect 6917 15855 6975 15861
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 8202 15852 8208 15904
rect 8260 15892 8266 15904
rect 8389 15895 8447 15901
rect 8389 15892 8401 15895
rect 8260 15864 8401 15892
rect 8260 15852 8266 15864
rect 8389 15861 8401 15864
rect 8435 15861 8447 15895
rect 9416 15892 9444 15991
rect 13722 15988 13728 16040
rect 13780 16028 13786 16040
rect 13909 16031 13967 16037
rect 13909 16028 13921 16031
rect 13780 16000 13921 16028
rect 13780 15988 13786 16000
rect 13909 15997 13921 16000
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 15997 14059 16031
rect 14001 15991 14059 15997
rect 14016 15960 14044 15991
rect 13372 15932 14044 15960
rect 14200 15960 14228 16068
rect 14274 16056 14280 16108
rect 14332 16096 14338 16108
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 14332 16068 14565 16096
rect 14332 16056 14338 16068
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 15102 16056 15108 16108
rect 15160 16096 15166 16108
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 15160 16068 15485 16096
rect 15160 16056 15166 16068
rect 15473 16065 15485 16068
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 16163 16068 17049 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 17037 16065 17049 16068
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16096 17923 16099
rect 18598 16096 18604 16108
rect 17911 16068 18604 16096
rect 17911 16065 17923 16068
rect 17865 16059 17923 16065
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 20254 16096 20260 16108
rect 20215 16068 20260 16096
rect 20254 16056 20260 16068
rect 20312 16056 20318 16108
rect 20530 16096 20536 16108
rect 20443 16068 20536 16096
rect 20530 16056 20536 16068
rect 20588 16056 20594 16108
rect 20809 16099 20867 16105
rect 20809 16065 20821 16099
rect 20855 16065 20867 16099
rect 21266 16096 21272 16108
rect 21227 16068 21272 16096
rect 20809 16059 20867 16065
rect 14461 16031 14519 16037
rect 14461 15997 14473 16031
rect 14507 16028 14519 16031
rect 15286 16028 15292 16040
rect 14507 16000 15292 16028
rect 14507 15997 14519 16000
rect 14461 15991 14519 15997
rect 15286 15988 15292 16000
rect 15344 15988 15350 16040
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 17126 16028 17132 16040
rect 16356 16000 17132 16028
rect 16356 15988 16362 16000
rect 17126 15988 17132 16000
rect 17184 15988 17190 16040
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 15997 17279 16031
rect 17221 15991 17279 15997
rect 14550 15960 14556 15972
rect 14200 15932 14556 15960
rect 9674 15892 9680 15904
rect 9416 15864 9680 15892
rect 8389 15855 8447 15861
rect 9674 15852 9680 15864
rect 9732 15892 9738 15904
rect 10873 15895 10931 15901
rect 10873 15892 10885 15895
rect 9732 15864 10885 15892
rect 9732 15852 9738 15864
rect 10873 15861 10885 15864
rect 10919 15861 10931 15895
rect 11238 15892 11244 15904
rect 11199 15864 11244 15892
rect 10873 15855 10931 15861
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 11974 15892 11980 15904
rect 11935 15864 11980 15892
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 12066 15852 12072 15904
rect 12124 15892 12130 15904
rect 13372 15892 13400 15932
rect 14550 15920 14556 15932
rect 14608 15920 14614 15972
rect 15304 15960 15332 15988
rect 17236 15960 17264 15991
rect 17770 15988 17776 16040
rect 17828 16028 17834 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17828 16000 18061 16028
rect 17828 15988 17834 16000
rect 18049 15997 18061 16000
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 16028 19027 16031
rect 19058 16028 19064 16040
rect 19015 16000 19064 16028
rect 19015 15997 19027 16000
rect 18969 15991 19027 15997
rect 19058 15988 19064 16000
rect 19116 15988 19122 16040
rect 20165 16031 20223 16037
rect 20165 15997 20177 16031
rect 20211 16028 20223 16031
rect 20824 16028 20852 16059
rect 21266 16056 21272 16068
rect 21324 16056 21330 16108
rect 20211 16000 20852 16028
rect 20211 15997 20223 16000
rect 20165 15991 20223 15997
rect 15304 15932 17264 15960
rect 12124 15864 13400 15892
rect 12124 15852 12130 15864
rect 13814 15852 13820 15904
rect 13872 15892 13878 15904
rect 15286 15892 15292 15904
rect 13872 15864 15292 15892
rect 13872 15852 13878 15864
rect 15286 15852 15292 15864
rect 15344 15892 15350 15904
rect 20180 15892 20208 15991
rect 21450 15892 21456 15904
rect 15344 15864 20208 15892
rect 21411 15864 21456 15892
rect 15344 15852 15350 15864
rect 21450 15852 21456 15864
rect 21508 15852 21514 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1762 15648 1768 15700
rect 1820 15688 1826 15700
rect 1857 15691 1915 15697
rect 1857 15688 1869 15691
rect 1820 15660 1869 15688
rect 1820 15648 1826 15660
rect 1857 15657 1869 15660
rect 1903 15657 1915 15691
rect 1857 15651 1915 15657
rect 1946 15648 1952 15700
rect 2004 15688 2010 15700
rect 2133 15691 2191 15697
rect 2133 15688 2145 15691
rect 2004 15660 2145 15688
rect 2004 15648 2010 15660
rect 2133 15657 2145 15660
rect 2179 15657 2191 15691
rect 2133 15651 2191 15657
rect 2222 15648 2228 15700
rect 2280 15688 2286 15700
rect 2409 15691 2467 15697
rect 2409 15688 2421 15691
rect 2280 15660 2421 15688
rect 2280 15648 2286 15660
rect 2409 15657 2421 15660
rect 2455 15657 2467 15691
rect 2409 15651 2467 15657
rect 2958 15648 2964 15700
rect 3016 15688 3022 15700
rect 3145 15691 3203 15697
rect 3145 15688 3157 15691
rect 3016 15660 3157 15688
rect 3016 15648 3022 15660
rect 3145 15657 3157 15660
rect 3191 15657 3203 15691
rect 3145 15651 3203 15657
rect 3234 15648 3240 15700
rect 3292 15688 3298 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 3292 15660 3801 15688
rect 3292 15648 3298 15660
rect 3789 15657 3801 15660
rect 3835 15657 3847 15691
rect 3789 15651 3847 15657
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 4617 15691 4675 15697
rect 4617 15688 4629 15691
rect 4212 15660 4629 15688
rect 4212 15648 4218 15660
rect 4617 15657 4629 15660
rect 4663 15657 4675 15691
rect 4982 15688 4988 15700
rect 4943 15660 4988 15688
rect 4617 15651 4675 15657
rect 4982 15648 4988 15660
rect 5040 15648 5046 15700
rect 5350 15648 5356 15700
rect 5408 15688 5414 15700
rect 5629 15691 5687 15697
rect 5629 15688 5641 15691
rect 5408 15660 5641 15688
rect 5408 15648 5414 15660
rect 5629 15657 5641 15660
rect 5675 15657 5687 15691
rect 5629 15651 5687 15657
rect 5718 15648 5724 15700
rect 5776 15688 5782 15700
rect 6365 15691 6423 15697
rect 6365 15688 6377 15691
rect 5776 15660 6377 15688
rect 5776 15648 5782 15660
rect 6365 15657 6377 15660
rect 6411 15657 6423 15691
rect 6365 15651 6423 15657
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7742 15688 7748 15700
rect 6972 15660 7748 15688
rect 6972 15648 6978 15660
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 8662 15648 8668 15700
rect 8720 15688 8726 15700
rect 10778 15688 10784 15700
rect 8720 15660 10784 15688
rect 8720 15648 8726 15660
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 11885 15691 11943 15697
rect 11885 15657 11897 15691
rect 11931 15688 11943 15691
rect 12066 15688 12072 15700
rect 11931 15660 12072 15688
rect 11931 15657 11943 15660
rect 11885 15651 11943 15657
rect 12066 15648 12072 15660
rect 12124 15648 12130 15700
rect 12250 15648 12256 15700
rect 12308 15688 12314 15700
rect 13170 15688 13176 15700
rect 12308 15660 13176 15688
rect 12308 15648 12314 15660
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 13357 15691 13415 15697
rect 13357 15657 13369 15691
rect 13403 15688 13415 15691
rect 13814 15688 13820 15700
rect 13403 15660 13820 15688
rect 13403 15657 13415 15660
rect 13357 15651 13415 15657
rect 13814 15648 13820 15660
rect 13872 15648 13878 15700
rect 14366 15648 14372 15700
rect 14424 15688 14430 15700
rect 17037 15691 17095 15697
rect 14424 15660 16988 15688
rect 14424 15648 14430 15660
rect 2774 15580 2780 15632
rect 2832 15620 2838 15632
rect 6181 15623 6239 15629
rect 6181 15620 6193 15623
rect 2832 15592 6193 15620
rect 2832 15580 2838 15592
rect 6181 15589 6193 15592
rect 6227 15589 6239 15623
rect 12710 15620 12716 15632
rect 6181 15583 6239 15589
rect 12452 15592 12716 15620
rect 198 15512 204 15564
rect 256 15552 262 15564
rect 256 15524 2728 15552
rect 256 15512 262 15524
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15484 2099 15487
rect 2222 15484 2228 15496
rect 2087 15456 2228 15484
rect 2087 15453 2099 15456
rect 2041 15447 2099 15453
rect 290 15376 296 15428
rect 348 15416 354 15428
rect 1688 15416 1716 15447
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 2314 15444 2320 15496
rect 2372 15484 2378 15496
rect 2590 15484 2596 15496
rect 2372 15456 2417 15484
rect 2551 15456 2596 15484
rect 2372 15444 2378 15456
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 2700 15493 2728 15524
rect 2866 15512 2872 15564
rect 2924 15552 2930 15564
rect 4062 15552 4068 15564
rect 2924 15524 4068 15552
rect 2924 15512 2930 15524
rect 4062 15512 4068 15524
rect 4120 15552 4126 15564
rect 4341 15555 4399 15561
rect 4341 15552 4353 15555
rect 4120 15524 4353 15552
rect 4120 15512 4126 15524
rect 4341 15521 4353 15524
rect 4387 15521 4399 15555
rect 4341 15515 4399 15521
rect 4614 15512 4620 15564
rect 4672 15552 4678 15564
rect 5074 15552 5080 15564
rect 4672 15524 5080 15552
rect 4672 15512 4678 15524
rect 5074 15512 5080 15524
rect 5132 15552 5138 15564
rect 5445 15555 5503 15561
rect 5445 15552 5457 15555
rect 5132 15524 5457 15552
rect 5132 15512 5138 15524
rect 5445 15521 5457 15524
rect 5491 15521 5503 15555
rect 5994 15552 6000 15564
rect 5955 15524 6000 15552
rect 5445 15515 5503 15521
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 7098 15552 7104 15564
rect 7059 15524 7104 15552
rect 7098 15512 7104 15524
rect 7156 15512 7162 15564
rect 10502 15552 10508 15564
rect 10463 15524 10508 15552
rect 10502 15512 10508 15524
rect 10560 15512 10566 15564
rect 12452 15561 12480 15592
rect 12710 15580 12716 15592
rect 12768 15580 12774 15632
rect 12802 15580 12808 15632
rect 12860 15620 12866 15632
rect 13722 15620 13728 15632
rect 12860 15592 13728 15620
rect 12860 15580 12866 15592
rect 13722 15580 13728 15592
rect 13780 15620 13786 15632
rect 14645 15623 14703 15629
rect 14645 15620 14657 15623
rect 13780 15592 14657 15620
rect 13780 15580 13786 15592
rect 14645 15589 14657 15592
rect 14691 15589 14703 15623
rect 16960 15620 16988 15660
rect 17037 15657 17049 15691
rect 17083 15688 17095 15691
rect 17310 15688 17316 15700
rect 17083 15660 17316 15688
rect 17083 15657 17095 15660
rect 17037 15651 17095 15657
rect 17310 15648 17316 15660
rect 17368 15648 17374 15700
rect 17420 15660 18460 15688
rect 17420 15620 17448 15660
rect 16960 15592 17448 15620
rect 14645 15583 14703 15589
rect 12437 15555 12495 15561
rect 12437 15521 12449 15555
rect 12483 15521 12495 15555
rect 12437 15515 12495 15521
rect 12618 15512 12624 15564
rect 12676 15552 12682 15564
rect 12676 15524 12721 15552
rect 12676 15512 12682 15524
rect 13170 15512 13176 15564
rect 13228 15552 13234 15564
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 13228 15524 14105 15552
rect 13228 15512 13234 15524
rect 14093 15521 14105 15524
rect 14139 15552 14151 15555
rect 14366 15552 14372 15564
rect 14139 15524 14372 15552
rect 14139 15521 14151 15524
rect 14093 15515 14151 15521
rect 14366 15512 14372 15524
rect 14424 15512 14430 15564
rect 18432 15552 18460 15660
rect 18598 15648 18604 15700
rect 18656 15688 18662 15700
rect 19245 15691 19303 15697
rect 19245 15688 19257 15691
rect 18656 15660 19257 15688
rect 18656 15648 18662 15660
rect 19245 15657 19257 15660
rect 19291 15657 19303 15691
rect 19245 15651 19303 15657
rect 19426 15648 19432 15700
rect 19484 15688 19490 15700
rect 20530 15688 20536 15700
rect 19484 15660 20536 15688
rect 19484 15648 19490 15660
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 20717 15691 20775 15697
rect 20717 15657 20729 15691
rect 20763 15688 20775 15691
rect 21266 15688 21272 15700
rect 20763 15660 21272 15688
rect 20763 15657 20775 15660
rect 20717 15651 20775 15657
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 18506 15580 18512 15632
rect 18564 15620 18570 15632
rect 20349 15623 20407 15629
rect 20349 15620 20361 15623
rect 18564 15592 20361 15620
rect 18564 15580 18570 15592
rect 20349 15589 20361 15592
rect 20395 15589 20407 15623
rect 20349 15583 20407 15589
rect 18432 15524 19104 15552
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15484 2743 15487
rect 2774 15484 2780 15496
rect 2731 15456 2780 15484
rect 2731 15453 2743 15456
rect 2685 15447 2743 15453
rect 2774 15444 2780 15456
rect 2832 15444 2838 15496
rect 2958 15484 2964 15496
rect 2919 15456 2964 15484
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 3050 15444 3056 15496
rect 3108 15484 3114 15496
rect 3237 15487 3295 15493
rect 3237 15484 3249 15487
rect 3108 15456 3249 15484
rect 3108 15444 3114 15456
rect 3237 15453 3249 15456
rect 3283 15453 3295 15487
rect 3237 15447 3295 15453
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15453 4859 15487
rect 4801 15447 4859 15453
rect 2406 15416 2412 15428
rect 348 15388 1624 15416
rect 1688 15388 2412 15416
rect 348 15376 354 15388
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 1596 15348 1624 15388
rect 2406 15376 2412 15388
rect 2464 15376 2470 15428
rect 2976 15416 3004 15444
rect 2746 15388 3004 15416
rect 4816 15416 4844 15447
rect 4982 15444 4988 15496
rect 5040 15484 5046 15496
rect 5169 15487 5227 15493
rect 5169 15484 5181 15487
rect 5040 15456 5181 15484
rect 5040 15444 5046 15456
rect 5169 15453 5181 15456
rect 5215 15453 5227 15487
rect 5169 15447 5227 15453
rect 5350 15416 5356 15428
rect 4816 15388 5356 15416
rect 2746 15348 2774 15388
rect 5350 15376 5356 15388
rect 5408 15376 5414 15428
rect 6012 15416 6040 15512
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15484 7435 15487
rect 7926 15484 7932 15496
rect 7423 15456 7932 15484
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 7926 15444 7932 15456
rect 7984 15484 7990 15496
rect 8202 15484 8208 15496
rect 7984 15456 8208 15484
rect 7984 15444 7990 15456
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15484 8999 15487
rect 9674 15484 9680 15496
rect 8987 15456 9680 15484
rect 8987 15453 8999 15456
rect 8941 15447 8999 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 11698 15484 11704 15496
rect 10284 15456 11704 15484
rect 10284 15444 10290 15456
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 11974 15444 11980 15496
rect 12032 15484 12038 15496
rect 12526 15484 12532 15496
rect 12032 15456 12532 15484
rect 12032 15444 12038 15456
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 13817 15487 13875 15493
rect 13817 15453 13829 15487
rect 13863 15484 13875 15487
rect 14274 15484 14280 15496
rect 13863 15456 14280 15484
rect 13863 15453 13875 15456
rect 13817 15447 13875 15453
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 15013 15487 15071 15493
rect 15013 15453 15025 15487
rect 15059 15484 15071 15487
rect 15102 15484 15108 15496
rect 15059 15456 15108 15484
rect 15059 15453 15071 15456
rect 15013 15447 15071 15453
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 15473 15487 15531 15493
rect 15473 15453 15485 15487
rect 15519 15484 15531 15487
rect 15565 15487 15623 15493
rect 15565 15484 15577 15487
rect 15519 15456 15577 15484
rect 15519 15453 15531 15456
rect 15473 15447 15531 15453
rect 15565 15453 15577 15456
rect 15611 15484 15623 15487
rect 15832 15487 15890 15493
rect 15832 15484 15844 15487
rect 15611 15456 15700 15484
rect 15611 15453 15623 15456
rect 15565 15447 15623 15453
rect 7644 15419 7702 15425
rect 6012 15388 7604 15416
rect 1596 15320 2774 15348
rect 2869 15351 2927 15357
rect 2869 15317 2881 15351
rect 2915 15348 2927 15351
rect 3050 15348 3056 15360
rect 2915 15320 3056 15348
rect 2915 15317 2927 15320
rect 2869 15311 2927 15317
rect 3050 15308 3056 15320
rect 3108 15308 3114 15360
rect 3326 15308 3332 15360
rect 3384 15348 3390 15360
rect 3421 15351 3479 15357
rect 3421 15348 3433 15351
rect 3384 15320 3433 15348
rect 3384 15308 3390 15320
rect 3421 15317 3433 15320
rect 3467 15317 3479 15351
rect 3421 15311 3479 15317
rect 3605 15351 3663 15357
rect 3605 15317 3617 15351
rect 3651 15348 3663 15351
rect 4154 15348 4160 15360
rect 3651 15320 4160 15348
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 4154 15308 4160 15320
rect 4212 15308 4218 15360
rect 4249 15351 4307 15357
rect 4249 15317 4261 15351
rect 4295 15348 4307 15351
rect 4890 15348 4896 15360
rect 4295 15320 4896 15348
rect 4295 15317 4307 15320
rect 4249 15311 4307 15317
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 5905 15351 5963 15357
rect 5905 15317 5917 15351
rect 5951 15348 5963 15351
rect 5994 15348 6000 15360
rect 5951 15320 6000 15348
rect 5951 15317 5963 15320
rect 5905 15311 5963 15317
rect 5994 15308 6000 15320
rect 6052 15308 6058 15360
rect 6546 15348 6552 15360
rect 6507 15320 6552 15348
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 6914 15348 6920 15360
rect 6875 15320 6920 15348
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 7576 15348 7604 15388
rect 7644 15385 7656 15419
rect 7690 15416 7702 15419
rect 8662 15416 8668 15428
rect 7690 15388 8668 15416
rect 7690 15385 7702 15388
rect 7644 15379 7702 15385
rect 8662 15376 8668 15388
rect 8720 15376 8726 15428
rect 9214 15425 9220 15428
rect 9208 15416 9220 15425
rect 8772 15388 9220 15416
rect 8110 15348 8116 15360
rect 7064 15320 7109 15348
rect 7576 15320 8116 15348
rect 7064 15308 7070 15320
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 8772 15357 8800 15388
rect 9208 15379 9220 15388
rect 9214 15376 9220 15379
rect 9272 15376 9278 15428
rect 10772 15419 10830 15425
rect 10772 15385 10784 15419
rect 10818 15416 10830 15419
rect 10870 15416 10876 15428
rect 10818 15388 10876 15416
rect 10818 15385 10830 15388
rect 10772 15379 10830 15385
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 11422 15376 11428 15428
rect 11480 15416 11486 15428
rect 12066 15416 12072 15428
rect 11480 15388 12072 15416
rect 11480 15376 11486 15388
rect 12066 15376 12072 15388
rect 12124 15376 12130 15428
rect 12713 15419 12771 15425
rect 12713 15385 12725 15419
rect 12759 15416 12771 15419
rect 13446 15416 13452 15428
rect 12759 15388 13452 15416
rect 12759 15385 12771 15388
rect 12713 15379 12771 15385
rect 13446 15376 13452 15388
rect 13504 15376 13510 15428
rect 8757 15351 8815 15357
rect 8757 15317 8769 15351
rect 8803 15317 8815 15351
rect 8757 15311 8815 15317
rect 9398 15308 9404 15360
rect 9456 15348 9462 15360
rect 10321 15351 10379 15357
rect 10321 15348 10333 15351
rect 9456 15320 10333 15348
rect 9456 15308 9462 15320
rect 10321 15317 10333 15320
rect 10367 15317 10379 15351
rect 10321 15311 10379 15317
rect 12986 15308 12992 15360
rect 13044 15348 13050 15360
rect 13081 15351 13139 15357
rect 13081 15348 13093 15351
rect 13044 15320 13093 15348
rect 13044 15308 13050 15320
rect 13081 15317 13093 15320
rect 13127 15317 13139 15351
rect 13630 15348 13636 15360
rect 13591 15320 13636 15348
rect 13081 15311 13139 15317
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 14182 15308 14188 15360
rect 14240 15348 14246 15360
rect 14277 15351 14335 15357
rect 14277 15348 14289 15351
rect 14240 15320 14289 15348
rect 14240 15308 14246 15320
rect 14277 15317 14289 15320
rect 14323 15317 14335 15351
rect 14550 15348 14556 15360
rect 14511 15320 14556 15348
rect 14277 15311 14335 15317
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 15010 15308 15016 15360
rect 15068 15348 15074 15360
rect 15289 15351 15347 15357
rect 15289 15348 15301 15351
rect 15068 15320 15301 15348
rect 15068 15308 15074 15320
rect 15289 15317 15301 15320
rect 15335 15317 15347 15351
rect 15672 15348 15700 15456
rect 15764 15456 15844 15484
rect 15764 15428 15792 15456
rect 15832 15453 15844 15456
rect 15878 15453 15890 15487
rect 15832 15447 15890 15453
rect 16942 15444 16948 15496
rect 17000 15484 17006 15496
rect 18417 15487 18475 15493
rect 18417 15484 18429 15487
rect 17000 15456 18429 15484
rect 17000 15444 17006 15456
rect 18417 15453 18429 15456
rect 18463 15484 18475 15487
rect 18969 15487 19027 15493
rect 18969 15484 18981 15487
rect 18463 15456 18981 15484
rect 18463 15453 18475 15456
rect 18417 15447 18475 15453
rect 18969 15453 18981 15456
rect 19015 15453 19027 15487
rect 19076 15484 19104 15524
rect 19242 15512 19248 15564
rect 19300 15552 19306 15564
rect 19797 15555 19855 15561
rect 19797 15552 19809 15555
rect 19300 15524 19809 15552
rect 19300 15512 19306 15524
rect 19797 15521 19809 15524
rect 19843 15521 19855 15555
rect 19797 15515 19855 15521
rect 19426 15484 19432 15496
rect 19076 15456 19432 15484
rect 18969 15447 19027 15453
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 19518 15444 19524 15496
rect 19576 15484 19582 15496
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19576 15456 19717 15484
rect 19576 15444 19582 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 20070 15484 20076 15496
rect 20031 15456 20076 15484
rect 19705 15447 19763 15453
rect 20070 15444 20076 15456
rect 20128 15444 20134 15496
rect 20364 15484 20392 15583
rect 20533 15487 20591 15493
rect 20533 15484 20545 15487
rect 20364 15456 20545 15484
rect 20533 15453 20545 15456
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 20809 15487 20867 15493
rect 20809 15453 20821 15487
rect 20855 15453 20867 15487
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 20809 15447 20867 15453
rect 21008 15456 21281 15484
rect 15746 15376 15752 15428
rect 15804 15376 15810 15428
rect 16960 15416 16988 15444
rect 17770 15416 17776 15428
rect 15948 15388 16988 15416
rect 17144 15388 17776 15416
rect 15948 15348 15976 15388
rect 17144 15360 17172 15388
rect 17770 15376 17776 15388
rect 17828 15416 17834 15428
rect 18150 15419 18208 15425
rect 18150 15416 18162 15419
rect 17828 15388 18162 15416
rect 17828 15376 17834 15388
rect 18150 15385 18162 15388
rect 18196 15385 18208 15419
rect 18150 15379 18208 15385
rect 18693 15419 18751 15425
rect 18693 15385 18705 15419
rect 18739 15416 18751 15419
rect 19613 15419 19671 15425
rect 19613 15416 19625 15419
rect 18739 15388 19625 15416
rect 18739 15385 18751 15388
rect 18693 15379 18751 15385
rect 19613 15385 19625 15388
rect 19659 15385 19671 15419
rect 20824 15416 20852 15447
rect 19613 15379 19671 15385
rect 20272 15388 20852 15416
rect 15672 15320 15976 15348
rect 16945 15351 17003 15357
rect 15289 15311 15347 15317
rect 16945 15317 16957 15351
rect 16991 15348 17003 15351
rect 17126 15348 17132 15360
rect 16991 15320 17132 15348
rect 16991 15317 17003 15320
rect 16945 15311 17003 15317
rect 17126 15308 17132 15320
rect 17184 15308 17190 15360
rect 18782 15348 18788 15360
rect 18743 15320 18788 15348
rect 18782 15308 18788 15320
rect 18840 15308 18846 15360
rect 20272 15357 20300 15388
rect 21008 15357 21036 15456
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 20257 15351 20315 15357
rect 20257 15317 20269 15351
rect 20303 15317 20315 15351
rect 20257 15311 20315 15317
rect 20993 15351 21051 15357
rect 20993 15317 21005 15351
rect 21039 15317 21051 15351
rect 21174 15348 21180 15360
rect 21135 15320 21180 15348
rect 20993 15311 21051 15317
rect 21174 15308 21180 15320
rect 21232 15308 21238 15360
rect 21450 15348 21456 15360
rect 21411 15320 21456 15348
rect 21450 15308 21456 15320
rect 21508 15308 21514 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 2317 15147 2375 15153
rect 2317 15113 2329 15147
rect 2363 15113 2375 15147
rect 2317 15107 2375 15113
rect 1670 15008 1676 15020
rect 1631 14980 1676 15008
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 2038 15008 2044 15020
rect 1999 14980 2044 15008
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 14977 2191 15011
rect 2332 15008 2360 15107
rect 2406 15104 2412 15156
rect 2464 15144 2470 15156
rect 4617 15147 4675 15153
rect 4617 15144 4629 15147
rect 2464 15116 2509 15144
rect 2746 15116 4629 15144
rect 2464 15104 2470 15116
rect 2593 15011 2651 15017
rect 2593 15008 2605 15011
rect 2332 14980 2605 15008
rect 2133 14971 2191 14977
rect 2593 14977 2605 14980
rect 2639 14977 2651 15011
rect 2593 14971 2651 14977
rect 2148 14940 2176 14971
rect 2746 14940 2774 15116
rect 4617 15113 4629 15116
rect 4663 15113 4675 15147
rect 4617 15107 4675 15113
rect 5077 15147 5135 15153
rect 5077 15113 5089 15147
rect 5123 15144 5135 15147
rect 5445 15147 5503 15153
rect 5445 15144 5457 15147
rect 5123 15116 5457 15144
rect 5123 15113 5135 15116
rect 5077 15107 5135 15113
rect 5445 15113 5457 15116
rect 5491 15113 5503 15147
rect 5445 15107 5503 15113
rect 5905 15147 5963 15153
rect 5905 15113 5917 15147
rect 5951 15144 5963 15147
rect 6546 15144 6552 15156
rect 5951 15116 6552 15144
rect 5951 15113 5963 15116
rect 5905 15107 5963 15113
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 6917 15147 6975 15153
rect 6917 15113 6929 15147
rect 6963 15144 6975 15147
rect 7006 15144 7012 15156
rect 6963 15116 7012 15144
rect 6963 15113 6975 15116
rect 6917 15107 6975 15113
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 7374 15104 7380 15156
rect 7432 15144 7438 15156
rect 7432 15116 7477 15144
rect 7432 15104 7438 15116
rect 7742 15104 7748 15156
rect 7800 15144 7806 15156
rect 8021 15147 8079 15153
rect 8021 15144 8033 15147
rect 7800 15116 8033 15144
rect 7800 15104 7806 15116
rect 8021 15113 8033 15116
rect 8067 15144 8079 15147
rect 8294 15144 8300 15156
rect 8067 15116 8300 15144
rect 8067 15113 8079 15116
rect 8021 15107 8079 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 8478 15144 8484 15156
rect 8439 15116 8484 15144
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 8570 15104 8576 15156
rect 8628 15144 8634 15156
rect 8941 15147 8999 15153
rect 8628 15116 8673 15144
rect 8628 15104 8634 15116
rect 8941 15113 8953 15147
rect 8987 15144 8999 15147
rect 9582 15144 9588 15156
rect 8987 15116 9588 15144
rect 8987 15113 8999 15116
rect 8941 15107 8999 15113
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 9769 15147 9827 15153
rect 9769 15113 9781 15147
rect 9815 15144 9827 15147
rect 9858 15144 9864 15156
rect 9815 15116 9864 15144
rect 9815 15113 9827 15116
rect 9769 15107 9827 15113
rect 9858 15104 9864 15116
rect 9916 15104 9922 15156
rect 12989 15147 13047 15153
rect 10069 15116 12388 15144
rect 3912 15079 3970 15085
rect 3912 15045 3924 15079
rect 3958 15076 3970 15079
rect 4062 15076 4068 15088
rect 3958 15048 4068 15076
rect 3958 15045 3970 15048
rect 3912 15039 3970 15045
rect 4062 15036 4068 15048
rect 4120 15076 4126 15088
rect 5534 15076 5540 15088
rect 4120 15048 5540 15076
rect 4120 15036 4126 15048
rect 5534 15036 5540 15048
rect 5592 15036 5598 15088
rect 6748 15048 6914 15076
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 15008 4215 15011
rect 4246 15008 4252 15020
rect 4203 14980 4252 15008
rect 4203 14977 4215 14980
rect 4157 14971 4215 14977
rect 4246 14968 4252 14980
rect 4304 14968 4310 15020
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 15008 4399 15011
rect 4522 15008 4528 15020
rect 4387 14980 4528 15008
rect 4387 14977 4399 14980
rect 4341 14971 4399 14977
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 4798 14968 4804 15020
rect 4856 15008 4862 15020
rect 4985 15011 5043 15017
rect 4985 15008 4997 15011
rect 4856 14980 4997 15008
rect 4856 14968 4862 14980
rect 4985 14977 4997 14980
rect 5031 14977 5043 15011
rect 5810 15008 5816 15020
rect 5771 14980 5816 15008
rect 4985 14971 5043 14977
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 5902 14968 5908 15020
rect 5960 15008 5966 15020
rect 6748 15017 6776 15048
rect 6733 15011 6791 15017
rect 6733 15008 6745 15011
rect 5960 14980 6745 15008
rect 5960 14968 5966 14980
rect 6733 14977 6745 14980
rect 6779 14977 6791 15011
rect 6886 15008 6914 15048
rect 9122 15036 9128 15088
rect 9180 15076 9186 15088
rect 9401 15079 9459 15085
rect 9401 15076 9413 15079
rect 9180 15048 9413 15076
rect 9180 15036 9186 15048
rect 9401 15045 9413 15048
rect 9447 15045 9459 15079
rect 9401 15039 9459 15045
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 6886 14980 7297 15008
rect 6733 14971 6791 14977
rect 7285 14977 7297 14980
rect 7331 15008 7343 15011
rect 8202 15008 8208 15020
rect 7331 14980 8208 15008
rect 7331 14977 7343 14980
rect 7285 14971 7343 14977
rect 8202 14968 8208 14980
rect 8260 15008 8266 15020
rect 10069 15008 10097 15116
rect 10410 15076 10416 15088
rect 8260 14980 10097 15008
rect 10152 15048 10416 15076
rect 8260 14968 8266 14980
rect 5258 14940 5264 14952
rect 2148 14912 2774 14940
rect 5219 14912 5264 14940
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 5997 14943 6055 14949
rect 5997 14940 6009 14943
rect 5684 14912 6009 14940
rect 5684 14900 5690 14912
rect 5997 14909 6009 14912
rect 6043 14909 6055 14943
rect 5997 14903 6055 14909
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 7190 14940 7196 14952
rect 6687 14912 7196 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 7558 14940 7564 14952
rect 7519 14912 7564 14940
rect 7558 14900 7564 14912
rect 7616 14900 7622 14952
rect 8389 14943 8447 14949
rect 8389 14909 8401 14943
rect 8435 14940 8447 14943
rect 9214 14940 9220 14952
rect 8435 14912 9220 14940
rect 8435 14909 8447 14912
rect 8389 14903 8447 14909
rect 9214 14900 9220 14912
rect 9272 14900 9278 14952
rect 9309 14943 9367 14949
rect 9309 14909 9321 14943
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 1854 14872 1860 14884
rect 1815 14844 1860 14872
rect 1854 14832 1860 14844
rect 1912 14832 1918 14884
rect 2777 14875 2835 14881
rect 2777 14841 2789 14875
rect 2823 14872 2835 14875
rect 2866 14872 2872 14884
rect 2823 14844 2872 14872
rect 2823 14841 2835 14844
rect 2777 14835 2835 14841
rect 2866 14832 2872 14844
rect 2924 14832 2930 14884
rect 4522 14872 4528 14884
rect 4483 14844 4528 14872
rect 4522 14832 4528 14844
rect 4580 14832 4586 14884
rect 6454 14872 6460 14884
rect 6415 14844 6460 14872
rect 6454 14832 6460 14844
rect 6512 14832 6518 14884
rect 6546 14832 6552 14884
rect 6604 14872 6610 14884
rect 6822 14872 6828 14884
rect 6604 14844 6828 14872
rect 6604 14832 6610 14844
rect 6822 14832 6828 14844
rect 6880 14832 6886 14884
rect 7006 14832 7012 14884
rect 7064 14872 7070 14884
rect 9122 14872 9128 14884
rect 7064 14844 9128 14872
rect 7064 14832 7070 14844
rect 9122 14832 9128 14844
rect 9180 14832 9186 14884
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 4338 14764 4344 14816
rect 4396 14804 4402 14816
rect 5350 14804 5356 14816
rect 4396 14776 5356 14804
rect 4396 14764 4402 14776
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 5994 14764 6000 14816
rect 6052 14804 6058 14816
rect 7834 14804 7840 14816
rect 6052 14776 7840 14804
rect 6052 14764 6058 14776
rect 7834 14764 7840 14776
rect 7892 14764 7898 14816
rect 9232 14804 9260 14900
rect 9324 14872 9352 14903
rect 9674 14900 9680 14952
rect 9732 14940 9738 14952
rect 10152 14940 10180 15048
rect 10410 15036 10416 15048
rect 10468 15036 10474 15088
rect 11333 15079 11391 15085
rect 11333 15045 11345 15079
rect 11379 15076 11391 15079
rect 11885 15079 11943 15085
rect 11885 15076 11897 15079
rect 11379 15048 11897 15076
rect 11379 15045 11391 15048
rect 11333 15039 11391 15045
rect 11885 15045 11897 15048
rect 11931 15076 11943 15079
rect 12250 15076 12256 15088
rect 11931 15048 12256 15076
rect 11931 15045 11943 15048
rect 11885 15039 11943 15045
rect 12250 15036 12256 15048
rect 12308 15036 12314 15088
rect 12360 15076 12388 15116
rect 12989 15113 13001 15147
rect 13035 15144 13047 15147
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 13035 15116 13461 15144
rect 13035 15113 13047 15116
rect 12989 15107 13047 15113
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 13909 15147 13967 15153
rect 13909 15144 13921 15147
rect 13872 15116 13921 15144
rect 13872 15104 13878 15116
rect 13909 15113 13921 15116
rect 13955 15113 13967 15147
rect 14458 15144 14464 15156
rect 14419 15116 14464 15144
rect 13909 15107 13967 15113
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 16942 15144 16948 15156
rect 16903 15116 16948 15144
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 19153 15147 19211 15153
rect 17236 15116 19104 15144
rect 12360 15048 13032 15076
rect 10229 15011 10287 15017
rect 10229 14977 10241 15011
rect 10275 15008 10287 15011
rect 10689 15011 10747 15017
rect 10689 15008 10701 15011
rect 10275 14980 10701 15008
rect 10275 14977 10287 14980
rect 10229 14971 10287 14977
rect 10689 14977 10701 14980
rect 10735 14977 10747 15011
rect 10689 14971 10747 14977
rect 11698 14968 11704 15020
rect 11756 15008 11762 15020
rect 11977 15011 12035 15017
rect 11977 15008 11989 15011
rect 11756 14980 11989 15008
rect 11756 14968 11762 14980
rect 11977 14977 11989 14980
rect 12023 15008 12035 15011
rect 12023 14980 12480 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 10318 14940 10324 14952
rect 9732 14912 10180 14940
rect 10279 14912 10324 14940
rect 9732 14900 9738 14912
rect 10318 14900 10324 14912
rect 10376 14900 10382 14952
rect 10410 14900 10416 14952
rect 10468 14940 10474 14952
rect 10468 14912 10513 14940
rect 10468 14900 10474 14912
rect 10778 14900 10784 14952
rect 10836 14940 10842 14952
rect 12069 14943 12127 14949
rect 12069 14940 12081 14943
rect 10836 14912 12081 14940
rect 10836 14900 10842 14912
rect 12069 14909 12081 14912
rect 12115 14909 12127 14943
rect 12069 14903 12127 14909
rect 11517 14875 11575 14881
rect 11517 14872 11529 14875
rect 9324 14844 11529 14872
rect 11517 14841 11529 14844
rect 11563 14841 11575 14875
rect 11517 14835 11575 14841
rect 9398 14804 9404 14816
rect 9232 14776 9404 14804
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 9490 14764 9496 14816
rect 9548 14804 9554 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9548 14776 9873 14804
rect 9548 14764 9554 14776
rect 9861 14773 9873 14776
rect 9907 14773 9919 14807
rect 10962 14804 10968 14816
rect 10923 14776 10968 14804
rect 9861 14767 9919 14773
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 12452 14813 12480 14980
rect 12710 14940 12716 14952
rect 12671 14912 12716 14940
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 12897 14943 12955 14949
rect 12897 14909 12909 14943
rect 12943 14909 12955 14943
rect 13004 14940 13032 15048
rect 13630 15036 13636 15088
rect 13688 15076 13694 15088
rect 13688 15048 14320 15076
rect 13688 15036 13694 15048
rect 13814 15008 13820 15020
rect 13775 14980 13820 15008
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14292 15017 14320 15048
rect 14826 15036 14832 15088
rect 14884 15076 14890 15088
rect 17236 15076 17264 15116
rect 14884 15048 17264 15076
rect 14884 15036 14890 15048
rect 17310 15036 17316 15088
rect 17368 15076 17374 15088
rect 17466 15079 17524 15085
rect 17466 15076 17478 15079
rect 17368 15048 17478 15076
rect 17368 15036 17374 15048
rect 17466 15045 17478 15048
rect 17512 15045 17524 15079
rect 19076 15076 19104 15116
rect 19153 15113 19165 15147
rect 19199 15144 19211 15147
rect 19518 15144 19524 15156
rect 19199 15116 19524 15144
rect 19199 15113 19211 15116
rect 19153 15107 19211 15113
rect 19518 15104 19524 15116
rect 19576 15104 19582 15156
rect 19889 15147 19947 15153
rect 19889 15113 19901 15147
rect 19935 15144 19947 15147
rect 20254 15144 20260 15156
rect 19935 15116 20260 15144
rect 19935 15113 19947 15116
rect 19889 15107 19947 15113
rect 20254 15104 20260 15116
rect 20312 15104 20318 15156
rect 22646 15144 22652 15156
rect 20548 15116 22652 15144
rect 19978 15076 19984 15088
rect 19076 15048 19984 15076
rect 17466 15039 17524 15045
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 20073 15079 20131 15085
rect 20073 15045 20085 15079
rect 20119 15076 20131 15079
rect 20548 15076 20576 15116
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 20119 15048 20576 15076
rect 20625 15079 20683 15085
rect 20119 15045 20131 15048
rect 20073 15039 20131 15045
rect 20625 15045 20637 15079
rect 20671 15076 20683 15079
rect 22186 15076 22192 15088
rect 20671 15048 22192 15076
rect 20671 15045 20683 15048
rect 20625 15039 20683 15045
rect 22186 15036 22192 15048
rect 22244 15036 22250 15088
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 15010 15008 15016 15020
rect 14424 14980 15016 15008
rect 14424 14968 14430 14980
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 16022 15008 16028 15020
rect 15983 14980 16028 15008
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 15008 17187 15011
rect 17221 15011 17279 15017
rect 17221 15008 17233 15011
rect 17175 14980 17233 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 17221 14977 17233 14980
rect 17267 15008 17279 15011
rect 18046 15008 18052 15020
rect 17267 14980 18052 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 18046 14968 18052 14980
rect 18104 14968 18110 15020
rect 19702 15008 19708 15020
rect 19663 14980 19708 15008
rect 19702 14968 19708 14980
rect 19760 14968 19766 15020
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 20901 15011 20959 15017
rect 20901 15008 20913 15011
rect 20772 14980 20913 15008
rect 20772 14968 20778 14980
rect 20901 14977 20913 14980
rect 20947 14977 20959 15011
rect 20901 14971 20959 14977
rect 20990 14968 20996 15020
rect 21048 15008 21054 15020
rect 21269 15011 21327 15017
rect 21269 15008 21281 15011
rect 21048 14980 21281 15008
rect 21048 14968 21054 14980
rect 21269 14977 21281 14980
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 13722 14940 13728 14952
rect 13004 14912 13728 14940
rect 12897 14903 12955 14909
rect 12912 14816 12940 14903
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 13998 14940 14004 14952
rect 13959 14912 14004 14940
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 15746 14940 15752 14952
rect 15707 14912 15752 14940
rect 15746 14900 15752 14912
rect 15804 14900 15810 14952
rect 15930 14940 15936 14952
rect 15891 14912 15936 14940
rect 15930 14900 15936 14912
rect 15988 14900 15994 14952
rect 18598 14900 18604 14952
rect 18656 14940 18662 14952
rect 20165 14943 20223 14949
rect 20165 14940 20177 14943
rect 18656 14912 20177 14940
rect 18656 14900 18662 14912
rect 20165 14909 20177 14912
rect 20211 14909 20223 14943
rect 20165 14903 20223 14909
rect 20809 14943 20867 14949
rect 20809 14909 20821 14943
rect 20855 14940 20867 14943
rect 21358 14940 21364 14952
rect 20855 14912 21364 14940
rect 20855 14909 20867 14912
rect 20809 14903 20867 14909
rect 21358 14900 21364 14912
rect 21416 14900 21422 14952
rect 21082 14872 21088 14884
rect 21043 14844 21088 14872
rect 21082 14832 21088 14844
rect 21140 14832 21146 14884
rect 22278 14872 22284 14884
rect 21284 14844 22284 14872
rect 12437 14807 12495 14813
rect 12437 14773 12449 14807
rect 12483 14804 12495 14807
rect 12618 14804 12624 14816
rect 12483 14776 12624 14804
rect 12483 14773 12495 14776
rect 12437 14767 12495 14773
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 12894 14764 12900 14816
rect 12952 14764 12958 14816
rect 13354 14804 13360 14816
rect 13315 14776 13360 14804
rect 13354 14764 13360 14776
rect 13412 14764 13418 14816
rect 15194 14804 15200 14816
rect 15155 14776 15200 14804
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 16393 14807 16451 14813
rect 16393 14773 16405 14807
rect 16439 14804 16451 14807
rect 16850 14804 16856 14816
rect 16439 14776 16856 14804
rect 16439 14773 16451 14776
rect 16393 14767 16451 14773
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18601 14807 18659 14813
rect 18601 14804 18613 14807
rect 18012 14776 18613 14804
rect 18012 14764 18018 14776
rect 18601 14773 18613 14776
rect 18647 14773 18659 14807
rect 18601 14767 18659 14773
rect 20441 14807 20499 14813
rect 20441 14773 20453 14807
rect 20487 14804 20499 14807
rect 21284 14804 21312 14844
rect 22278 14832 22284 14844
rect 22336 14832 22342 14884
rect 21450 14804 21456 14816
rect 20487 14776 21312 14804
rect 21411 14776 21456 14804
rect 20487 14773 20499 14776
rect 20441 14767 20499 14773
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 1670 14560 1676 14612
rect 1728 14600 1734 14612
rect 2133 14603 2191 14609
rect 2133 14600 2145 14603
rect 1728 14572 2145 14600
rect 1728 14560 1734 14572
rect 2133 14569 2145 14572
rect 2179 14569 2191 14603
rect 2133 14563 2191 14569
rect 2222 14560 2228 14612
rect 2280 14600 2286 14612
rect 2409 14603 2467 14609
rect 2409 14600 2421 14603
rect 2280 14572 2421 14600
rect 2280 14560 2286 14572
rect 2409 14569 2421 14572
rect 2455 14569 2467 14603
rect 2409 14563 2467 14569
rect 2958 14560 2964 14612
rect 3016 14600 3022 14612
rect 3513 14603 3571 14609
rect 3513 14600 3525 14603
rect 3016 14572 3525 14600
rect 3016 14560 3022 14572
rect 3513 14569 3525 14572
rect 3559 14569 3571 14603
rect 4798 14600 4804 14612
rect 4759 14572 4804 14600
rect 3513 14563 3571 14569
rect 4798 14560 4804 14572
rect 4856 14560 4862 14612
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 6273 14603 6331 14609
rect 6273 14600 6285 14603
rect 5316 14572 6285 14600
rect 5316 14560 5322 14572
rect 6273 14569 6285 14572
rect 6319 14600 6331 14603
rect 6822 14600 6828 14612
rect 6319 14572 6828 14600
rect 6319 14569 6331 14572
rect 6273 14563 6331 14569
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 6972 14572 7941 14600
rect 6972 14560 6978 14572
rect 7929 14569 7941 14572
rect 7975 14569 7987 14603
rect 7929 14563 7987 14569
rect 8570 14560 8576 14612
rect 8628 14600 8634 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 8628 14572 9965 14600
rect 8628 14560 8634 14572
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 9953 14563 10011 14569
rect 10502 14560 10508 14612
rect 10560 14600 10566 14612
rect 10560 14572 15139 14600
rect 10560 14560 10566 14572
rect 1857 14535 1915 14541
rect 1857 14501 1869 14535
rect 1903 14501 1915 14535
rect 1857 14495 1915 14501
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1872 14396 1900 14495
rect 2038 14492 2044 14544
rect 2096 14532 2102 14544
rect 2685 14535 2743 14541
rect 2685 14532 2697 14535
rect 2096 14504 2697 14532
rect 2096 14492 2102 14504
rect 2685 14501 2697 14504
rect 2731 14501 2743 14535
rect 2685 14495 2743 14501
rect 2774 14492 2780 14544
rect 2832 14532 2838 14544
rect 3789 14535 3847 14541
rect 3789 14532 3801 14535
rect 2832 14504 3801 14532
rect 2832 14492 2838 14504
rect 3789 14501 3801 14504
rect 3835 14501 3847 14535
rect 3789 14495 3847 14501
rect 9861 14535 9919 14541
rect 9861 14501 9873 14535
rect 9907 14532 9919 14535
rect 10686 14532 10692 14544
rect 9907 14504 10692 14532
rect 9907 14501 9919 14504
rect 9861 14495 9919 14501
rect 10686 14492 10692 14504
rect 10744 14492 10750 14544
rect 3234 14464 3240 14476
rect 2332 14436 3240 14464
rect 2038 14396 2044 14408
rect 1719 14368 1900 14396
rect 1999 14368 2044 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 2332 14405 2360 14436
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 4249 14467 4307 14473
rect 4249 14433 4261 14467
rect 4295 14464 4307 14467
rect 8478 14464 8484 14476
rect 4295 14436 5028 14464
rect 4295 14433 4307 14436
rect 4249 14427 4307 14433
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14365 2375 14399
rect 2317 14359 2375 14365
rect 2406 14356 2412 14408
rect 2464 14396 2470 14408
rect 2593 14399 2651 14405
rect 2593 14396 2605 14399
rect 2464 14368 2605 14396
rect 2464 14356 2470 14368
rect 2593 14365 2605 14368
rect 2639 14365 2651 14399
rect 2593 14359 2651 14365
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14396 2927 14399
rect 2961 14399 3019 14405
rect 2961 14396 2973 14399
rect 2915 14368 2973 14396
rect 2915 14365 2927 14368
rect 2869 14359 2927 14365
rect 2961 14365 2973 14368
rect 3007 14396 3019 14399
rect 4893 14399 4951 14405
rect 3007 14368 4844 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 2056 14328 2084 14356
rect 3329 14331 3387 14337
rect 3329 14328 3341 14331
rect 2056 14300 3341 14328
rect 3329 14297 3341 14300
rect 3375 14328 3387 14331
rect 3878 14328 3884 14340
rect 3375 14300 3884 14328
rect 3375 14297 3387 14300
rect 3329 14291 3387 14297
rect 3878 14288 3884 14300
rect 3936 14288 3942 14340
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 4338 14260 4344 14272
rect 4299 14232 4344 14260
rect 4338 14220 4344 14232
rect 4396 14220 4402 14272
rect 4430 14220 4436 14272
rect 4488 14260 4494 14272
rect 4816 14260 4844 14368
rect 4893 14365 4905 14399
rect 4939 14365 4951 14399
rect 5000 14396 5028 14436
rect 7760 14436 8484 14464
rect 5160 14399 5218 14405
rect 5160 14396 5172 14399
rect 5000 14368 5172 14396
rect 4893 14359 4951 14365
rect 5160 14365 5172 14368
rect 5206 14396 5218 14399
rect 5626 14396 5632 14408
rect 5206 14368 5632 14396
rect 5206 14365 5218 14368
rect 5160 14359 5218 14365
rect 4908 14328 4936 14359
rect 5626 14356 5632 14368
rect 5684 14356 5690 14408
rect 6454 14356 6460 14408
rect 6512 14396 6518 14408
rect 7282 14396 7288 14408
rect 6512 14368 7288 14396
rect 6512 14356 6518 14368
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7558 14396 7564 14408
rect 7616 14405 7622 14408
rect 7616 14399 7639 14405
rect 7491 14368 7564 14396
rect 7558 14356 7564 14368
rect 7627 14396 7639 14399
rect 7760 14396 7788 14436
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 8938 14424 8944 14476
rect 8996 14464 9002 14476
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 8996 14436 9229 14464
rect 8996 14424 9002 14436
rect 9217 14433 9229 14436
rect 9263 14433 9275 14467
rect 10318 14464 10324 14476
rect 9217 14427 9275 14433
rect 9324 14436 10324 14464
rect 7627 14368 7788 14396
rect 7837 14399 7895 14405
rect 7627 14365 7639 14368
rect 7616 14359 7639 14365
rect 7837 14365 7849 14399
rect 7883 14396 7895 14399
rect 7926 14396 7932 14408
rect 7883 14368 7932 14396
rect 7883 14365 7895 14368
rect 7837 14359 7895 14365
rect 7616 14356 7622 14359
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 8389 14399 8447 14405
rect 8389 14396 8401 14399
rect 8352 14368 8401 14396
rect 8352 14356 8358 14368
rect 8389 14365 8401 14368
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 9033 14399 9091 14405
rect 9033 14365 9045 14399
rect 9079 14396 9091 14399
rect 9324 14396 9352 14436
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14464 10655 14467
rect 10778 14464 10784 14476
rect 10643 14436 10784 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 10778 14424 10784 14436
rect 10836 14424 10842 14476
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 13909 14467 13967 14473
rect 13909 14464 13921 14467
rect 13872 14436 13921 14464
rect 13872 14424 13878 14436
rect 13909 14433 13921 14436
rect 13955 14433 13967 14467
rect 15111 14464 15139 14572
rect 15746 14560 15752 14612
rect 15804 14600 15810 14612
rect 16945 14603 17003 14609
rect 16945 14600 16957 14603
rect 15804 14572 16957 14600
rect 15804 14560 15810 14572
rect 16945 14569 16957 14572
rect 16991 14600 17003 14603
rect 16991 14572 17448 14600
rect 16991 14569 17003 14572
rect 16945 14563 17003 14569
rect 16850 14492 16856 14544
rect 16908 14532 16914 14544
rect 17420 14532 17448 14572
rect 17494 14560 17500 14612
rect 17552 14600 17558 14612
rect 17773 14603 17831 14609
rect 17773 14600 17785 14603
rect 17552 14572 17785 14600
rect 17552 14560 17558 14572
rect 17773 14569 17785 14572
rect 17819 14569 17831 14603
rect 17773 14563 17831 14569
rect 19337 14603 19395 14609
rect 19337 14569 19349 14603
rect 19383 14600 19395 14603
rect 19518 14600 19524 14612
rect 19383 14572 19524 14600
rect 19383 14569 19395 14572
rect 19337 14563 19395 14569
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 20714 14600 20720 14612
rect 20675 14572 20720 14600
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 20990 14600 20996 14612
rect 20951 14572 20996 14600
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 19058 14532 19064 14544
rect 16908 14504 17356 14532
rect 17420 14504 19064 14532
rect 16908 14492 16914 14504
rect 17126 14464 17132 14476
rect 15111 14436 15700 14464
rect 17087 14436 17132 14464
rect 13909 14427 13967 14433
rect 9490 14396 9496 14408
rect 9079 14368 9352 14396
rect 9451 14368 9496 14396
rect 9079 14365 9091 14368
rect 9033 14359 9091 14365
rect 9490 14356 9496 14368
rect 9548 14356 9554 14408
rect 10336 14396 10364 14424
rect 10686 14396 10692 14408
rect 10336 14368 10692 14396
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 11882 14356 11888 14408
rect 11940 14405 11946 14408
rect 11940 14396 11952 14405
rect 12161 14399 12219 14405
rect 11940 14368 11985 14396
rect 11940 14359 11952 14368
rect 12161 14365 12173 14399
rect 12207 14396 12219 14399
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 12207 14368 12265 14396
rect 12207 14365 12219 14368
rect 12161 14359 12219 14365
rect 12253 14365 12265 14368
rect 12299 14396 12311 14399
rect 13630 14396 13636 14408
rect 12299 14368 13636 14396
rect 12299 14365 12311 14368
rect 12253 14359 12311 14365
rect 11940 14356 11946 14359
rect 4982 14328 4988 14340
rect 4908 14300 4988 14328
rect 4982 14288 4988 14300
rect 5040 14288 5046 14340
rect 10413 14331 10471 14337
rect 10413 14328 10425 14331
rect 5368 14300 10425 14328
rect 5368 14260 5396 14300
rect 10413 14297 10425 14300
rect 10459 14328 10471 14331
rect 10870 14328 10876 14340
rect 10459 14300 10876 14328
rect 10459 14297 10471 14300
rect 10413 14291 10471 14297
rect 10870 14288 10876 14300
rect 10928 14288 10934 14340
rect 11698 14288 11704 14340
rect 11756 14328 11762 14340
rect 12176 14328 12204 14359
rect 13630 14356 13636 14368
rect 13688 14356 13694 14408
rect 14093 14399 14151 14405
rect 14093 14365 14105 14399
rect 14139 14396 14151 14399
rect 14182 14396 14188 14408
rect 14139 14368 14188 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14182 14356 14188 14368
rect 14240 14396 14246 14408
rect 15565 14399 15623 14405
rect 15565 14396 15577 14399
rect 14240 14368 15577 14396
rect 14240 14356 14246 14368
rect 15565 14365 15577 14368
rect 15611 14365 15623 14399
rect 15672 14396 15700 14436
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 17328 14473 17356 14504
rect 19058 14492 19064 14504
rect 19116 14492 19122 14544
rect 17313 14467 17371 14473
rect 17313 14433 17325 14467
rect 17359 14433 17371 14467
rect 17313 14427 17371 14433
rect 17770 14424 17776 14476
rect 17828 14464 17834 14476
rect 21085 14467 21143 14473
rect 21085 14464 21097 14467
rect 17828 14436 21097 14464
rect 17828 14424 17834 14436
rect 20824 14405 20852 14436
rect 21085 14433 21097 14436
rect 21131 14433 21143 14467
rect 21085 14427 21143 14433
rect 20349 14399 20407 14405
rect 20349 14396 20361 14399
rect 15672 14368 20361 14396
rect 15565 14359 15623 14365
rect 17144 14340 17172 14368
rect 20349 14365 20361 14368
rect 20395 14396 20407 14399
rect 20533 14399 20591 14405
rect 20533 14396 20545 14399
rect 20395 14368 20545 14396
rect 20395 14365 20407 14368
rect 20349 14359 20407 14365
rect 20533 14365 20545 14368
rect 20579 14365 20591 14399
rect 20533 14359 20591 14365
rect 20809 14399 20867 14405
rect 20809 14365 20821 14399
rect 20855 14365 20867 14399
rect 20809 14359 20867 14365
rect 20990 14356 20996 14408
rect 21048 14396 21054 14408
rect 21269 14399 21327 14405
rect 21269 14396 21281 14399
rect 21048 14368 21281 14396
rect 21048 14356 21054 14368
rect 21269 14365 21281 14368
rect 21315 14365 21327 14399
rect 21269 14359 21327 14365
rect 11756 14300 12204 14328
rect 12498 14331 12556 14337
rect 11756 14288 11762 14300
rect 12498 14297 12510 14331
rect 12544 14328 12556 14331
rect 12710 14328 12716 14340
rect 12544 14300 12716 14328
rect 12544 14297 12556 14300
rect 12498 14291 12556 14297
rect 4488 14232 4533 14260
rect 4816 14232 5396 14260
rect 4488 14220 4494 14232
rect 5442 14220 5448 14272
rect 5500 14260 5506 14272
rect 6457 14263 6515 14269
rect 6457 14260 6469 14263
rect 5500 14232 6469 14260
rect 5500 14220 5506 14232
rect 6457 14229 6469 14232
rect 6503 14260 6515 14263
rect 7098 14260 7104 14272
rect 6503 14232 7104 14260
rect 6503 14229 6515 14232
rect 6457 14223 6515 14229
rect 7098 14220 7104 14232
rect 7156 14220 7162 14272
rect 7834 14220 7840 14272
rect 7892 14260 7898 14272
rect 8297 14263 8355 14269
rect 8297 14260 8309 14263
rect 7892 14232 8309 14260
rect 7892 14220 7898 14232
rect 8297 14229 8309 14232
rect 8343 14260 8355 14263
rect 9306 14260 9312 14272
rect 8343 14232 9312 14260
rect 8343 14229 8355 14232
rect 8297 14223 8355 14229
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 9401 14263 9459 14269
rect 9401 14229 9413 14263
rect 9447 14260 9459 14263
rect 9858 14260 9864 14272
rect 9447 14232 9864 14260
rect 9447 14229 9459 14232
rect 9401 14223 9459 14229
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 10318 14260 10324 14272
rect 10279 14232 10324 14260
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 10781 14263 10839 14269
rect 10781 14229 10793 14263
rect 10827 14260 10839 14263
rect 12513 14260 12541 14291
rect 12710 14288 12716 14300
rect 12768 14288 12774 14340
rect 14338 14331 14396 14337
rect 14338 14328 14350 14331
rect 13648 14300 14350 14328
rect 10827 14232 12541 14260
rect 10827 14229 10839 14232
rect 10781 14223 10839 14229
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 13648 14269 13676 14300
rect 14338 14297 14350 14300
rect 14384 14297 14396 14331
rect 14338 14291 14396 14297
rect 14826 14288 14832 14340
rect 14884 14328 14890 14340
rect 15102 14328 15108 14340
rect 14884 14300 15108 14328
rect 14884 14288 14890 14300
rect 15102 14288 15108 14300
rect 15160 14328 15166 14340
rect 15838 14337 15844 14340
rect 15832 14328 15844 14337
rect 15160 14300 15700 14328
rect 15799 14300 15844 14328
rect 15160 14288 15166 14300
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 12860 14232 13645 14260
rect 12860 14220 12866 14232
rect 13633 14229 13645 14232
rect 13679 14229 13691 14263
rect 13633 14223 13691 14229
rect 15473 14263 15531 14269
rect 15473 14229 15485 14263
rect 15519 14260 15531 14263
rect 15562 14260 15568 14272
rect 15519 14232 15568 14260
rect 15519 14229 15531 14232
rect 15473 14223 15531 14229
rect 15562 14220 15568 14232
rect 15620 14220 15626 14272
rect 15672 14260 15700 14300
rect 15832 14291 15844 14300
rect 15838 14288 15844 14291
rect 15896 14288 15902 14340
rect 17126 14288 17132 14340
rect 17184 14288 17190 14340
rect 17236 14300 17601 14328
rect 17236 14260 17264 14300
rect 15672 14232 17264 14260
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 17573 14260 17601 14300
rect 18506 14288 18512 14340
rect 18564 14328 18570 14340
rect 19429 14331 19487 14337
rect 19429 14328 19441 14331
rect 18564 14300 19441 14328
rect 18564 14288 18570 14300
rect 19429 14297 19441 14300
rect 19475 14297 19487 14331
rect 19429 14291 19487 14297
rect 19889 14331 19947 14337
rect 19889 14297 19901 14331
rect 19935 14328 19947 14331
rect 20070 14328 20076 14340
rect 19935 14300 20076 14328
rect 19935 14297 19947 14300
rect 19889 14291 19947 14297
rect 20070 14288 20076 14300
rect 20128 14288 20134 14340
rect 20257 14331 20315 14337
rect 20257 14297 20269 14331
rect 20303 14328 20315 14331
rect 22922 14328 22928 14340
rect 20303 14300 22928 14328
rect 20303 14297 20315 14300
rect 20257 14291 20315 14297
rect 22922 14288 22928 14300
rect 22980 14288 22986 14340
rect 18322 14260 18328 14272
rect 17460 14232 17505 14260
rect 17573 14232 18328 14260
rect 17460 14220 17466 14232
rect 18322 14220 18328 14232
rect 18380 14260 18386 14272
rect 18874 14260 18880 14272
rect 18380 14232 18880 14260
rect 18380 14220 18386 14232
rect 18874 14220 18880 14232
rect 18932 14220 18938 14272
rect 19610 14260 19616 14272
rect 19571 14232 19616 14260
rect 19610 14220 19616 14232
rect 19668 14220 19674 14272
rect 19978 14260 19984 14272
rect 19939 14232 19984 14260
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 21450 14260 21456 14272
rect 21411 14232 21456 14260
rect 21450 14220 21456 14232
rect 21508 14220 21514 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 1857 14059 1915 14065
rect 1857 14025 1869 14059
rect 1903 14025 1915 14059
rect 1857 14019 1915 14025
rect 2225 14059 2283 14065
rect 2225 14025 2237 14059
rect 2271 14056 2283 14059
rect 2406 14056 2412 14068
rect 2271 14028 2412 14056
rect 2271 14025 2283 14028
rect 2225 14019 2283 14025
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 1872 13920 1900 14019
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 2593 14059 2651 14065
rect 2593 14025 2605 14059
rect 2639 14056 2651 14059
rect 3053 14059 3111 14065
rect 3053 14056 3065 14059
rect 2639 14028 3065 14056
rect 2639 14025 2651 14028
rect 2593 14019 2651 14025
rect 3053 14025 3065 14028
rect 3099 14025 3111 14059
rect 3053 14019 3111 14025
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 3476 14028 4936 14056
rect 3476 14016 3482 14028
rect 3234 13988 3240 14000
rect 2056 13960 3240 13988
rect 2056 13929 2084 13960
rect 3234 13948 3240 13960
rect 3292 13948 3298 14000
rect 4516 13991 4574 13997
rect 4516 13957 4528 13991
rect 4562 13988 4574 13991
rect 4798 13988 4804 14000
rect 4562 13960 4804 13988
rect 4562 13957 4574 13960
rect 4516 13951 4574 13957
rect 4798 13948 4804 13960
rect 4856 13948 4862 14000
rect 1719 13892 1900 13920
rect 2041 13923 2099 13929
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 2041 13889 2053 13923
rect 2087 13889 2099 13923
rect 2041 13883 2099 13889
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 3418 13920 3424 13932
rect 2731 13892 3280 13920
rect 3379 13892 3424 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13821 2835 13855
rect 3252 13852 3280 13892
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13920 3571 13923
rect 3878 13920 3884 13932
rect 3559 13892 3884 13920
rect 3559 13889 3571 13892
rect 3513 13883 3571 13889
rect 3878 13880 3884 13892
rect 3936 13880 3942 13932
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13920 4031 13923
rect 4062 13920 4068 13932
rect 4019 13892 4068 13920
rect 4019 13889 4031 13892
rect 3973 13883 4031 13889
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4246 13920 4252 13932
rect 4207 13892 4252 13920
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 4908 13920 4936 14028
rect 4982 14016 4988 14068
rect 5040 14056 5046 14068
rect 5626 14056 5632 14068
rect 5040 14028 5488 14056
rect 5587 14028 5632 14056
rect 5040 14016 5046 14028
rect 5460 13988 5488 14028
rect 5626 14016 5632 14028
rect 5684 14016 5690 14068
rect 6457 14059 6515 14065
rect 6457 14056 6469 14059
rect 5828 14028 6469 14056
rect 5828 13988 5856 14028
rect 6457 14025 6469 14028
rect 6503 14025 6515 14059
rect 7834 14056 7840 14068
rect 6457 14019 6515 14025
rect 6748 14028 7840 14056
rect 5902 13988 5908 14000
rect 5460 13960 5908 13988
rect 5902 13948 5908 13960
rect 5960 13948 5966 14000
rect 6748 13988 6776 14028
rect 7834 14016 7840 14028
rect 7892 14016 7898 14068
rect 8481 14059 8539 14065
rect 8481 14025 8493 14059
rect 8527 14025 8539 14059
rect 8481 14019 8539 14025
rect 8665 14059 8723 14065
rect 8665 14025 8677 14059
rect 8711 14056 8723 14059
rect 9398 14056 9404 14068
rect 8711 14028 9404 14056
rect 8711 14025 8723 14028
rect 8665 14019 8723 14025
rect 6012 13960 6776 13988
rect 6012 13929 6040 13960
rect 6822 13948 6828 14000
rect 6880 13988 6886 14000
rect 7346 13991 7404 13997
rect 7346 13988 7358 13991
rect 6880 13960 7358 13988
rect 6880 13948 6886 13960
rect 7346 13957 7358 13960
rect 7392 13957 7404 13991
rect 8496 13988 8524 14019
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 9858 14056 9864 14068
rect 9548 14028 9720 14056
rect 9819 14028 9864 14056
rect 9548 14016 9554 14028
rect 9508 13988 9536 14016
rect 8496 13960 9536 13988
rect 7346 13951 7404 13957
rect 5997 13923 6055 13929
rect 5997 13920 6009 13923
rect 4908 13892 6009 13920
rect 5997 13889 6009 13892
rect 6043 13889 6055 13923
rect 5997 13883 6055 13889
rect 6641 13923 6699 13929
rect 6641 13889 6653 13923
rect 6687 13920 6699 13923
rect 7101 13923 7159 13929
rect 7101 13920 7113 13923
rect 6687 13892 7113 13920
rect 6687 13889 6699 13892
rect 6641 13883 6699 13889
rect 7101 13889 7113 13892
rect 7147 13920 7159 13923
rect 7926 13920 7932 13932
rect 7147 13892 7932 13920
rect 7147 13889 7159 13892
rect 7101 13883 7159 13889
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 8110 13880 8116 13932
rect 8168 13920 8174 13932
rect 9030 13920 9036 13932
rect 8168 13892 9036 13920
rect 8168 13880 8174 13892
rect 9030 13880 9036 13892
rect 9088 13920 9094 13932
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 9088 13892 9505 13920
rect 9088 13880 9094 13892
rect 9493 13889 9505 13892
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 3326 13852 3332 13864
rect 3252 13824 3332 13852
rect 2777 13815 2835 13821
rect 2498 13744 2504 13796
rect 2556 13784 2562 13796
rect 2792 13784 2820 13815
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13821 3755 13855
rect 4154 13852 4160 13864
rect 4115 13824 4160 13852
rect 3697 13815 3755 13821
rect 2556 13756 2820 13784
rect 3712 13784 3740 13815
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 5258 13812 5264 13864
rect 5316 13852 5322 13864
rect 5721 13855 5779 13861
rect 5721 13852 5733 13855
rect 5316 13824 5733 13852
rect 5316 13812 5322 13824
rect 5721 13821 5733 13824
rect 5767 13821 5779 13855
rect 6733 13855 6791 13861
rect 6733 13852 6745 13855
rect 5721 13815 5779 13821
rect 5828 13824 6745 13852
rect 4246 13784 4252 13796
rect 3712 13756 4252 13784
rect 2556 13744 2562 13756
rect 4246 13744 4252 13756
rect 4304 13744 4310 13796
rect 5350 13744 5356 13796
rect 5408 13784 5414 13796
rect 5828 13784 5856 13824
rect 6733 13821 6745 13824
rect 6779 13821 6791 13855
rect 6914 13852 6920 13864
rect 6875 13824 6920 13852
rect 6733 13815 6791 13821
rect 6914 13812 6920 13824
rect 6972 13812 6978 13864
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 9692 13861 9720 14028
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10321 14059 10379 14065
rect 10321 14025 10333 14059
rect 10367 14056 10379 14059
rect 10502 14056 10508 14068
rect 10367 14028 10508 14056
rect 10367 14025 10379 14028
rect 10321 14019 10379 14025
rect 10502 14016 10508 14028
rect 10560 14016 10566 14068
rect 11054 14056 11060 14068
rect 11015 14028 11060 14056
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 11241 14059 11299 14065
rect 11241 14025 11253 14059
rect 11287 14056 11299 14059
rect 11790 14056 11796 14068
rect 11287 14028 11796 14056
rect 11287 14025 11299 14028
rect 11241 14019 11299 14025
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 12158 14056 12164 14068
rect 12119 14028 12164 14056
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 12250 14016 12256 14068
rect 12308 14056 12314 14068
rect 12710 14056 12716 14068
rect 12308 14028 12716 14056
rect 12308 14016 12314 14028
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 12894 14016 12900 14068
rect 12952 14056 12958 14068
rect 13357 14059 13415 14065
rect 13357 14056 13369 14059
rect 12952 14028 13369 14056
rect 12952 14016 12958 14028
rect 13357 14025 13369 14028
rect 13403 14025 13415 14059
rect 13357 14019 13415 14025
rect 13446 14016 13452 14068
rect 13504 14056 13510 14068
rect 13504 14028 13549 14056
rect 13504 14016 13510 14028
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 15657 14059 15715 14065
rect 13780 14028 15332 14056
rect 13780 14016 13786 14028
rect 9766 13948 9772 14000
rect 9824 13988 9830 14000
rect 11514 13988 11520 14000
rect 9824 13960 11376 13988
rect 11475 13960 11520 13988
rect 9824 13948 9830 13960
rect 10226 13920 10232 13932
rect 10187 13892 10232 13920
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 11348 13920 11376 13960
rect 11514 13948 11520 13960
rect 11572 13948 11578 14000
rect 15197 13991 15255 13997
rect 15197 13988 15209 13991
rect 11716 13960 15209 13988
rect 11716 13920 11744 13960
rect 15197 13957 15209 13960
rect 15243 13957 15255 13991
rect 15197 13951 15255 13957
rect 11348 13892 11744 13920
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12529 13923 12587 13929
rect 12032 13892 12434 13920
rect 12032 13880 12038 13892
rect 9677 13855 9735 13861
rect 8444 13824 9628 13852
rect 8444 13812 8450 13824
rect 6086 13784 6092 13796
rect 5408 13756 5856 13784
rect 5920 13756 6092 13784
rect 5408 13744 5414 13756
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 2314 13676 2320 13728
rect 2372 13716 2378 13728
rect 3970 13716 3976 13728
rect 2372 13688 3976 13716
rect 2372 13676 2378 13688
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 4982 13716 4988 13728
rect 4580 13688 4988 13716
rect 4580 13676 4586 13688
rect 4982 13676 4988 13688
rect 5040 13676 5046 13728
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 5920 13716 5948 13756
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 6178 13744 6184 13796
rect 6236 13784 6242 13796
rect 6638 13784 6644 13796
rect 6236 13756 6644 13784
rect 6236 13744 6242 13756
rect 6638 13744 6644 13756
rect 6696 13744 6702 13796
rect 8938 13784 8944 13796
rect 8899 13756 8944 13784
rect 8938 13744 8944 13756
rect 8996 13744 9002 13796
rect 9600 13784 9628 13824
rect 9677 13821 9689 13855
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 10410 13812 10416 13864
rect 10468 13852 10474 13864
rect 10870 13852 10876 13864
rect 10468 13824 10513 13852
rect 10831 13824 10876 13852
rect 10468 13812 10474 13824
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 11330 13812 11336 13864
rect 11388 13852 11394 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11388 13824 11713 13852
rect 11388 13812 11394 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 11790 13812 11796 13864
rect 11848 13852 11854 13864
rect 11885 13855 11943 13861
rect 11885 13852 11897 13855
rect 11848 13824 11897 13852
rect 11848 13812 11854 13824
rect 11885 13821 11897 13824
rect 11931 13821 11943 13855
rect 12250 13852 12256 13864
rect 12211 13824 12256 13852
rect 11885 13815 11943 13821
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 12406 13852 12434 13892
rect 12529 13889 12541 13923
rect 12575 13920 12587 13923
rect 12989 13923 13047 13929
rect 12575 13892 12940 13920
rect 12575 13889 12587 13892
rect 12529 13883 12587 13889
rect 12912 13861 12940 13892
rect 12989 13889 13001 13923
rect 13035 13920 13047 13923
rect 13446 13920 13452 13932
rect 13035 13892 13452 13920
rect 13035 13889 13047 13892
rect 12989 13883 13047 13889
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 13814 13920 13820 13932
rect 13775 13892 13820 13920
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 13909 13923 13967 13929
rect 13909 13889 13921 13923
rect 13955 13920 13967 13923
rect 14274 13920 14280 13932
rect 13955 13892 14280 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 14366 13880 14372 13932
rect 14424 13920 14430 13932
rect 15304 13929 15332 14028
rect 15657 14025 15669 14059
rect 15703 14056 15715 14059
rect 15930 14056 15936 14068
rect 15703 14028 15936 14056
rect 15703 14025 15715 14028
rect 15657 14019 15715 14025
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16485 14059 16543 14065
rect 16485 14025 16497 14059
rect 16531 14056 16543 14059
rect 17402 14056 17408 14068
rect 16531 14028 17408 14056
rect 16531 14025 16543 14028
rect 16485 14019 16543 14025
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 20990 14056 20996 14068
rect 20951 14028 20996 14056
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 15746 13948 15752 14000
rect 15804 13948 15810 14000
rect 18782 13988 18788 14000
rect 17696 13960 18788 13988
rect 14829 13923 14887 13929
rect 14424 13892 14469 13920
rect 14424 13880 14430 13892
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15289 13923 15347 13929
rect 15289 13920 15301 13923
rect 14875 13892 15301 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 15289 13889 15301 13892
rect 15335 13889 15347 13923
rect 15764 13920 15792 13948
rect 15764 13892 15884 13920
rect 15289 13883 15347 13889
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12406 13824 12817 13852
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 13998 13852 14004 13864
rect 12943 13824 14004 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 11606 13784 11612 13796
rect 9600 13756 11612 13784
rect 11606 13744 11612 13756
rect 11664 13744 11670 13796
rect 12820 13784 12848 13815
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 14093 13855 14151 13861
rect 14093 13821 14105 13855
rect 14139 13821 14151 13855
rect 14093 13815 14151 13821
rect 14108 13784 14136 13815
rect 14182 13812 14188 13864
rect 14240 13852 14246 13864
rect 15010 13852 15016 13864
rect 14240 13824 15016 13852
rect 14240 13812 14246 13824
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 15105 13855 15163 13861
rect 15105 13821 15117 13855
rect 15151 13852 15163 13855
rect 15746 13852 15752 13864
rect 15151 13824 15752 13852
rect 15151 13821 15163 13824
rect 15105 13815 15163 13821
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 15856 13861 15884 13892
rect 15930 13880 15936 13932
rect 15988 13920 15994 13932
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 15988 13892 16129 13920
rect 15988 13880 15994 13892
rect 16117 13889 16129 13892
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 17586 13880 17592 13932
rect 17644 13920 17650 13932
rect 17696 13929 17724 13960
rect 18782 13948 18788 13960
rect 18840 13948 18846 14000
rect 17954 13929 17960 13932
rect 17681 13923 17739 13929
rect 17681 13920 17693 13923
rect 17644 13892 17693 13920
rect 17644 13880 17650 13892
rect 17681 13889 17693 13892
rect 17727 13889 17739 13923
rect 17948 13920 17960 13929
rect 17915 13892 17960 13920
rect 17681 13883 17739 13889
rect 17948 13883 17960 13892
rect 17954 13880 17960 13883
rect 18012 13880 18018 13932
rect 19058 13880 19064 13932
rect 19116 13920 19122 13932
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19116 13892 19441 13920
rect 19116 13880 19122 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 19518 13880 19524 13932
rect 19576 13920 19582 13932
rect 20533 13923 20591 13929
rect 19576 13892 19621 13920
rect 19576 13880 19582 13892
rect 20533 13889 20545 13923
rect 20579 13889 20591 13923
rect 20533 13883 20591 13889
rect 15841 13855 15899 13861
rect 15841 13821 15853 13855
rect 15887 13821 15899 13855
rect 15841 13815 15899 13821
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13852 16083 13855
rect 16390 13852 16396 13864
rect 16071 13824 16396 13852
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13821 19303 13855
rect 20162 13852 20168 13864
rect 20123 13824 20168 13852
rect 19245 13815 19303 13821
rect 12820 13756 14136 13784
rect 16206 13744 16212 13796
rect 16264 13784 16270 13796
rect 17402 13784 17408 13796
rect 16264 13756 17408 13784
rect 16264 13744 16270 13756
rect 17402 13744 17408 13756
rect 17460 13744 17466 13796
rect 18966 13744 18972 13796
rect 19024 13784 19030 13796
rect 19260 13784 19288 13815
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20346 13852 20352 13864
rect 20307 13824 20352 13852
rect 20346 13812 20352 13824
rect 20404 13852 20410 13864
rect 20548 13852 20576 13883
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 20809 13923 20867 13929
rect 20809 13920 20821 13923
rect 20772 13892 20821 13920
rect 20772 13880 20778 13892
rect 20809 13889 20821 13892
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 20404 13824 20576 13852
rect 20824 13852 20852 13883
rect 20990 13880 20996 13932
rect 21048 13920 21054 13932
rect 21269 13923 21327 13929
rect 21269 13920 21281 13923
rect 21048 13892 21281 13920
rect 21048 13880 21054 13892
rect 21269 13889 21281 13892
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 21085 13855 21143 13861
rect 21085 13852 21097 13855
rect 20824 13824 21097 13852
rect 20404 13812 20410 13824
rect 21085 13821 21097 13824
rect 21131 13821 21143 13855
rect 21085 13815 21143 13821
rect 19024 13756 19288 13784
rect 20717 13787 20775 13793
rect 19024 13744 19030 13756
rect 20717 13753 20729 13787
rect 20763 13784 20775 13787
rect 21266 13784 21272 13796
rect 20763 13756 21272 13784
rect 20763 13753 20775 13756
rect 20717 13747 20775 13753
rect 21266 13744 21272 13756
rect 21324 13744 21330 13796
rect 5868 13688 5948 13716
rect 5868 13676 5874 13688
rect 7834 13676 7840 13728
rect 7892 13716 7898 13728
rect 8662 13716 8668 13728
rect 7892 13688 8668 13716
rect 7892 13676 7898 13688
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 9033 13719 9091 13725
rect 9033 13685 9045 13719
rect 9079 13716 9091 13719
rect 9122 13716 9128 13728
rect 9079 13688 9128 13716
rect 9079 13685 9091 13688
rect 9033 13679 9091 13685
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 9306 13676 9312 13728
rect 9364 13716 9370 13728
rect 9950 13716 9956 13728
rect 9364 13688 9956 13716
rect 9364 13676 9370 13688
rect 9950 13676 9956 13688
rect 10008 13716 10014 13728
rect 13814 13716 13820 13728
rect 10008 13688 13820 13716
rect 10008 13676 10014 13688
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 14366 13676 14372 13728
rect 14424 13716 14430 13728
rect 15746 13716 15752 13728
rect 14424 13688 15752 13716
rect 14424 13676 14430 13688
rect 15746 13676 15752 13688
rect 15804 13676 15810 13728
rect 17494 13676 17500 13728
rect 17552 13716 17558 13728
rect 18874 13716 18880 13728
rect 17552 13688 18880 13716
rect 17552 13676 17558 13688
rect 18874 13676 18880 13688
rect 18932 13716 18938 13728
rect 19061 13719 19119 13725
rect 19061 13716 19073 13719
rect 18932 13688 19073 13716
rect 18932 13676 18938 13688
rect 19061 13685 19073 13688
rect 19107 13685 19119 13719
rect 19886 13716 19892 13728
rect 19847 13688 19892 13716
rect 19061 13679 19119 13685
rect 19886 13676 19892 13688
rect 19944 13676 19950 13728
rect 21450 13716 21456 13728
rect 21411 13688 21456 13716
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 4157 13515 4215 13521
rect 4157 13481 4169 13515
rect 4203 13512 4215 13515
rect 4430 13512 4436 13524
rect 4203 13484 4436 13512
rect 4203 13481 4215 13484
rect 4157 13475 4215 13481
rect 4430 13472 4436 13484
rect 4488 13472 4494 13524
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 4580 13484 5856 13512
rect 4580 13472 4586 13484
rect 4338 13404 4344 13456
rect 4396 13444 4402 13456
rect 4985 13447 5043 13453
rect 4985 13444 4997 13447
rect 4396 13416 4997 13444
rect 4396 13404 4402 13416
rect 4985 13413 4997 13416
rect 5031 13413 5043 13447
rect 4985 13407 5043 13413
rect 4522 13376 4528 13388
rect 3528 13348 4528 13376
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 2038 13308 2044 13320
rect 1999 13280 2044 13308
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 3349 13311 3407 13317
rect 3349 13277 3361 13311
rect 3395 13308 3407 13311
rect 3528 13308 3556 13348
rect 4522 13336 4528 13348
rect 4580 13336 4586 13388
rect 4798 13336 4804 13388
rect 4856 13376 4862 13388
rect 5442 13376 5448 13388
rect 4856 13348 5448 13376
rect 4856 13336 4862 13348
rect 5442 13336 5448 13348
rect 5500 13376 5506 13388
rect 5537 13379 5595 13385
rect 5537 13376 5549 13379
rect 5500 13348 5549 13376
rect 5500 13336 5506 13348
rect 5537 13345 5549 13348
rect 5583 13345 5595 13379
rect 5828 13376 5856 13484
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 6917 13515 6975 13521
rect 6917 13512 6929 13515
rect 6144 13484 6929 13512
rect 6144 13472 6150 13484
rect 6917 13481 6929 13484
rect 6963 13481 6975 13515
rect 6917 13475 6975 13481
rect 8570 13472 8576 13524
rect 8628 13512 8634 13524
rect 11793 13515 11851 13521
rect 11793 13512 11805 13515
rect 8628 13484 11805 13512
rect 8628 13472 8634 13484
rect 11793 13481 11805 13484
rect 11839 13481 11851 13515
rect 11793 13475 11851 13481
rect 12066 13472 12072 13524
rect 12124 13472 12130 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12492 13484 12537 13512
rect 12492 13472 12498 13484
rect 13078 13472 13084 13524
rect 13136 13512 13142 13524
rect 13538 13512 13544 13524
rect 13136 13484 13544 13512
rect 13136 13472 13142 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 15841 13515 15899 13521
rect 15841 13512 15853 13515
rect 13872 13484 15853 13512
rect 13872 13472 13878 13484
rect 15841 13481 15853 13484
rect 15887 13512 15899 13515
rect 15930 13512 15936 13524
rect 15887 13484 15936 13512
rect 15887 13481 15899 13484
rect 15841 13475 15899 13481
rect 15930 13472 15936 13484
rect 15988 13472 15994 13524
rect 16022 13472 16028 13524
rect 16080 13512 16086 13524
rect 16209 13515 16267 13521
rect 16209 13512 16221 13515
rect 16080 13484 16221 13512
rect 16080 13472 16086 13484
rect 16209 13481 16221 13484
rect 16255 13481 16267 13515
rect 18966 13512 18972 13524
rect 18927 13484 18972 13512
rect 16209 13475 16267 13481
rect 18966 13472 18972 13484
rect 19024 13472 19030 13524
rect 19058 13472 19064 13524
rect 19116 13512 19122 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 19116 13484 19257 13512
rect 19116 13472 19122 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 19702 13472 19708 13524
rect 19760 13512 19766 13524
rect 20073 13515 20131 13521
rect 20073 13512 20085 13515
rect 19760 13484 20085 13512
rect 19760 13472 19766 13484
rect 20073 13481 20085 13484
rect 20119 13481 20131 13515
rect 20073 13475 20131 13481
rect 7006 13404 7012 13456
rect 7064 13444 7070 13456
rect 8021 13447 8079 13453
rect 8021 13444 8033 13447
rect 7064 13416 8033 13444
rect 7064 13404 7070 13416
rect 8021 13413 8033 13416
rect 8067 13413 8079 13447
rect 8941 13447 8999 13453
rect 8941 13444 8953 13447
rect 8021 13407 8079 13413
rect 8588 13416 8953 13444
rect 5828 13348 7052 13376
rect 5537 13339 5595 13345
rect 3395 13280 3556 13308
rect 3605 13311 3663 13317
rect 3395 13277 3407 13280
rect 3349 13271 3407 13277
rect 3605 13277 3617 13311
rect 3651 13308 3663 13311
rect 3970 13308 3976 13320
rect 3651 13280 3976 13308
rect 3651 13277 3663 13280
rect 3605 13271 3663 13277
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 5353 13311 5411 13317
rect 5353 13308 5365 13311
rect 4120 13280 5365 13308
rect 4120 13268 4126 13280
rect 5353 13277 5365 13280
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 5626 13268 5632 13320
rect 5684 13308 5690 13320
rect 5684 13280 6500 13308
rect 5684 13268 5690 13280
rect 842 13200 848 13252
rect 900 13240 906 13252
rect 4338 13240 4344 13252
rect 900 13212 4344 13240
rect 900 13200 906 13212
rect 4338 13200 4344 13212
rect 4396 13200 4402 13252
rect 4430 13200 4436 13252
rect 4488 13240 4494 13252
rect 4617 13243 4675 13249
rect 4617 13240 4629 13243
rect 4488 13212 4629 13240
rect 4488 13200 4494 13212
rect 4617 13209 4629 13212
rect 4663 13209 4675 13243
rect 4617 13203 4675 13209
rect 5534 13200 5540 13252
rect 5592 13240 5598 13252
rect 5813 13243 5871 13249
rect 5813 13240 5825 13243
rect 5592 13212 5825 13240
rect 5592 13200 5598 13212
rect 5813 13209 5825 13212
rect 5859 13209 5871 13243
rect 5994 13240 6000 13252
rect 5955 13212 6000 13240
rect 5813 13203 5871 13209
rect 5994 13200 6000 13212
rect 6052 13200 6058 13252
rect 6472 13249 6500 13280
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 6733 13311 6791 13317
rect 6733 13308 6745 13311
rect 6604 13280 6745 13308
rect 6604 13268 6610 13280
rect 6733 13277 6745 13280
rect 6779 13277 6791 13311
rect 7024 13308 7052 13348
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 8588 13385 8616 13416
rect 8941 13413 8953 13416
rect 8987 13444 8999 13447
rect 9214 13444 9220 13456
rect 8987 13416 9220 13444
rect 8987 13413 8999 13416
rect 8941 13407 8999 13413
rect 9214 13404 9220 13416
rect 9272 13404 9278 13456
rect 10594 13404 10600 13456
rect 10652 13444 10658 13456
rect 11333 13447 11391 13453
rect 10652 13416 11284 13444
rect 10652 13404 10658 13416
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 7156 13348 7481 13376
rect 7156 13336 7162 13348
rect 7469 13345 7481 13348
rect 7515 13345 7527 13379
rect 8573 13379 8631 13385
rect 8573 13376 8585 13379
rect 7469 13339 7527 13345
rect 7567 13348 8585 13376
rect 7567 13308 7595 13348
rect 8573 13345 8585 13348
rect 8619 13345 8631 13379
rect 10965 13379 11023 13385
rect 10965 13376 10977 13379
rect 8573 13339 8631 13345
rect 10612 13348 10977 13376
rect 7024 13280 7595 13308
rect 8389 13311 8447 13317
rect 6733 13271 6791 13277
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 9490 13308 9496 13320
rect 8435 13280 9496 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 10321 13311 10379 13317
rect 10321 13308 10333 13311
rect 9824 13280 10333 13308
rect 9824 13268 9830 13280
rect 10321 13277 10333 13280
rect 10367 13277 10379 13311
rect 10321 13271 10379 13277
rect 6457 13243 6515 13249
rect 6457 13209 6469 13243
rect 6503 13240 6515 13243
rect 6638 13240 6644 13252
rect 6503 13212 6644 13240
rect 6503 13209 6515 13212
rect 6457 13203 6515 13209
rect 6638 13200 6644 13212
rect 6696 13200 6702 13252
rect 7285 13243 7343 13249
rect 7285 13209 7297 13243
rect 7331 13240 7343 13243
rect 8481 13243 8539 13249
rect 7331 13212 7880 13240
rect 7331 13209 7343 13212
rect 7285 13203 7343 13209
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 1854 13172 1860 13184
rect 1815 13144 1860 13172
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 2222 13172 2228 13184
rect 2183 13144 2228 13172
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 2774 13132 2780 13184
rect 2832 13172 2838 13184
rect 3789 13175 3847 13181
rect 3789 13172 3801 13175
rect 2832 13144 3801 13172
rect 2832 13132 2838 13144
rect 3789 13141 3801 13144
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 3878 13132 3884 13184
rect 3936 13172 3942 13184
rect 3973 13175 4031 13181
rect 3973 13172 3985 13175
rect 3936 13144 3985 13172
rect 3936 13132 3942 13144
rect 3973 13141 3985 13144
rect 4019 13141 4031 13175
rect 3973 13135 4031 13141
rect 4525 13175 4583 13181
rect 4525 13141 4537 13175
rect 4571 13172 4583 13175
rect 5258 13172 5264 13184
rect 4571 13144 5264 13172
rect 4571 13141 4583 13144
rect 4525 13135 4583 13141
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 5442 13172 5448 13184
rect 5403 13144 5448 13172
rect 5442 13132 5448 13144
rect 5500 13172 5506 13184
rect 6178 13172 6184 13184
rect 5500 13144 6184 13172
rect 5500 13132 5506 13144
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 6546 13172 6552 13184
rect 6507 13144 6552 13172
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 7374 13132 7380 13184
rect 7432 13172 7438 13184
rect 7852 13181 7880 13212
rect 8481 13209 8493 13243
rect 8527 13240 8539 13243
rect 8527 13212 9444 13240
rect 8527 13209 8539 13212
rect 8481 13203 8539 13209
rect 7837 13175 7895 13181
rect 7432 13144 7477 13172
rect 7432 13132 7438 13144
rect 7837 13141 7849 13175
rect 7883 13172 7895 13175
rect 8110 13172 8116 13184
rect 7883 13144 8116 13172
rect 7883 13141 7895 13144
rect 7837 13135 7895 13141
rect 8110 13132 8116 13144
rect 8168 13172 8174 13184
rect 9306 13172 9312 13184
rect 8168 13144 9312 13172
rect 8168 13132 8174 13144
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 9416 13172 9444 13212
rect 9582 13200 9588 13252
rect 9640 13240 9646 13252
rect 10042 13240 10048 13252
rect 10100 13249 10106 13252
rect 9640 13212 10048 13240
rect 9640 13200 9646 13212
rect 10042 13200 10048 13212
rect 10100 13240 10112 13249
rect 10612 13240 10640 13348
rect 10965 13345 10977 13348
rect 11011 13345 11023 13379
rect 11256 13376 11284 13416
rect 11333 13413 11345 13447
rect 11379 13444 11391 13447
rect 12084 13444 12112 13472
rect 12250 13444 12256 13456
rect 11379 13416 12256 13444
rect 11379 13413 11391 13416
rect 11333 13407 11391 13413
rect 12250 13404 12256 13416
rect 12308 13404 12314 13456
rect 12526 13444 12532 13456
rect 12487 13416 12532 13444
rect 12526 13404 12532 13416
rect 12584 13404 12590 13456
rect 13449 13447 13507 13453
rect 13449 13413 13461 13447
rect 13495 13444 13507 13447
rect 14366 13444 14372 13456
rect 13495 13416 14372 13444
rect 13495 13413 13507 13416
rect 13449 13407 13507 13413
rect 14366 13404 14372 13416
rect 14424 13404 14430 13456
rect 15749 13447 15807 13453
rect 15749 13413 15761 13447
rect 15795 13413 15807 13447
rect 15749 13407 15807 13413
rect 12069 13379 12127 13385
rect 11256 13348 11928 13376
rect 10965 13339 11023 13345
rect 10778 13308 10784 13320
rect 10739 13280 10784 13308
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 11701 13311 11759 13317
rect 11701 13277 11713 13311
rect 11747 13308 11759 13311
rect 11790 13308 11796 13320
rect 11747 13280 11796 13308
rect 11747 13277 11759 13280
rect 11701 13271 11759 13277
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 11900 13308 11928 13348
rect 12069 13345 12081 13379
rect 12115 13376 12127 13379
rect 12158 13376 12164 13388
rect 12115 13348 12164 13376
rect 12115 13345 12127 13348
rect 12069 13339 12127 13345
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 12802 13376 12808 13388
rect 12763 13348 12808 13376
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 12986 13376 12992 13388
rect 12947 13348 12992 13376
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 15764 13376 15792 13407
rect 15838 13376 15844 13388
rect 15751 13348 15844 13376
rect 15838 13336 15844 13348
rect 15896 13376 15902 13388
rect 16853 13379 16911 13385
rect 16853 13376 16865 13379
rect 15896 13348 16865 13376
rect 15896 13336 15902 13348
rect 16853 13345 16865 13348
rect 16899 13376 16911 13379
rect 16942 13376 16948 13388
rect 16899 13348 16948 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 17586 13376 17592 13388
rect 17328 13348 17592 13376
rect 13081 13311 13139 13317
rect 11900 13280 12572 13308
rect 10100 13212 10640 13240
rect 10100 13203 10112 13212
rect 10100 13200 10106 13203
rect 10686 13200 10692 13252
rect 10744 13240 10750 13252
rect 10744 13212 11560 13240
rect 10744 13200 10750 13212
rect 10413 13175 10471 13181
rect 10413 13172 10425 13175
rect 9416 13144 10425 13172
rect 10413 13141 10425 13144
rect 10459 13141 10471 13175
rect 10413 13135 10471 13141
rect 10594 13132 10600 13184
rect 10652 13172 10658 13184
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10652 13144 10885 13172
rect 10652 13132 10658 13144
rect 10873 13141 10885 13144
rect 10919 13141 10931 13175
rect 10873 13135 10931 13141
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 11330 13172 11336 13184
rect 11204 13144 11336 13172
rect 11204 13132 11210 13144
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 11532 13181 11560 13212
rect 11606 13200 11612 13252
rect 11664 13240 11670 13252
rect 12544 13240 12572 13280
rect 13081 13277 13093 13311
rect 13127 13308 13139 13311
rect 13354 13308 13360 13320
rect 13127 13280 13360 13308
rect 13127 13277 13139 13280
rect 13081 13271 13139 13277
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 13630 13308 13636 13320
rect 13591 13280 13636 13308
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 14369 13311 14427 13317
rect 14369 13308 14381 13311
rect 13872 13280 14381 13308
rect 13872 13268 13878 13280
rect 14369 13277 14381 13280
rect 14415 13308 14427 13311
rect 15102 13308 15108 13320
rect 14415 13280 15108 13308
rect 14415 13277 14427 13280
rect 14369 13271 14427 13277
rect 15102 13268 15108 13280
rect 15160 13308 15166 13320
rect 15378 13308 15384 13320
rect 15160 13280 15384 13308
rect 15160 13268 15166 13280
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 17328 13317 17356 13348
rect 17586 13336 17592 13348
rect 17644 13336 17650 13388
rect 18874 13336 18880 13388
rect 18932 13376 18938 13388
rect 19797 13379 19855 13385
rect 19797 13376 19809 13379
rect 18932 13348 19809 13376
rect 18932 13336 18938 13348
rect 19797 13345 19809 13348
rect 19843 13345 19855 13379
rect 19797 13339 19855 13345
rect 20530 13336 20536 13388
rect 20588 13376 20594 13388
rect 20625 13379 20683 13385
rect 20625 13376 20637 13379
rect 20588 13348 20637 13376
rect 20588 13336 20594 13348
rect 20625 13345 20637 13348
rect 20671 13345 20683 13379
rect 20625 13339 20683 13345
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13277 17371 13311
rect 17313 13271 17371 13277
rect 17494 13268 17500 13320
rect 17552 13308 17558 13320
rect 17845 13311 17903 13317
rect 17845 13308 17857 13311
rect 17552 13280 17857 13308
rect 17552 13268 17558 13280
rect 17845 13277 17857 13280
rect 17891 13277 17903 13311
rect 17845 13271 17903 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13308 19671 13311
rect 19702 13308 19708 13320
rect 19659 13280 19708 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 19886 13268 19892 13320
rect 19944 13308 19950 13320
rect 20441 13311 20499 13317
rect 20441 13308 20453 13311
rect 19944 13280 20453 13308
rect 19944 13268 19950 13280
rect 20441 13277 20453 13280
rect 20487 13277 20499 13311
rect 20901 13311 20959 13317
rect 20901 13308 20913 13311
rect 20441 13271 20499 13277
rect 20640 13280 20913 13308
rect 20640 13252 20668 13280
rect 20901 13277 20913 13280
rect 20947 13277 20959 13311
rect 21266 13308 21272 13320
rect 21227 13280 21272 13308
rect 20901 13271 20959 13277
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 14458 13240 14464 13252
rect 11664 13212 12296 13240
rect 12544 13212 14464 13240
rect 11664 13200 11670 13212
rect 11517 13175 11575 13181
rect 11517 13141 11529 13175
rect 11563 13172 11575 13175
rect 12158 13172 12164 13184
rect 11563 13144 12164 13172
rect 11563 13141 11575 13144
rect 11517 13135 11575 13141
rect 12158 13132 12164 13144
rect 12216 13132 12222 13184
rect 12268 13172 12296 13212
rect 14458 13200 14464 13212
rect 14516 13200 14522 13252
rect 14636 13243 14694 13249
rect 14636 13209 14648 13243
rect 14682 13240 14694 13243
rect 15194 13240 15200 13252
rect 14682 13212 15200 13240
rect 14682 13209 14694 13212
rect 14636 13203 14694 13209
rect 15194 13200 15200 13212
rect 15252 13200 15258 13252
rect 16577 13243 16635 13249
rect 16577 13209 16589 13243
rect 16623 13240 16635 13243
rect 17678 13240 17684 13252
rect 16623 13212 17684 13240
rect 16623 13209 16635 13212
rect 16577 13203 16635 13209
rect 17678 13200 17684 13212
rect 17736 13200 17742 13252
rect 18230 13200 18236 13252
rect 18288 13240 18294 13252
rect 20533 13243 20591 13249
rect 20533 13240 20545 13243
rect 18288 13212 20545 13240
rect 18288 13200 18294 13212
rect 20533 13209 20545 13212
rect 20579 13209 20591 13243
rect 20533 13203 20591 13209
rect 20622 13200 20628 13252
rect 20680 13200 20686 13252
rect 16025 13175 16083 13181
rect 16025 13172 16037 13175
rect 12268 13144 16037 13172
rect 16025 13141 16037 13144
rect 16071 13172 16083 13175
rect 16298 13172 16304 13184
rect 16071 13144 16304 13172
rect 16071 13141 16083 13144
rect 16025 13135 16083 13141
rect 16298 13132 16304 13144
rect 16356 13172 16362 13184
rect 16669 13175 16727 13181
rect 16669 13172 16681 13175
rect 16356 13144 16681 13172
rect 16356 13132 16362 13144
rect 16669 13141 16681 13144
rect 16715 13141 16727 13175
rect 17218 13172 17224 13184
rect 17179 13144 17224 13172
rect 16669 13135 16727 13141
rect 17218 13132 17224 13144
rect 17276 13132 17282 13184
rect 17497 13175 17555 13181
rect 17497 13141 17509 13175
rect 17543 13172 17555 13175
rect 18322 13172 18328 13184
rect 17543 13144 18328 13172
rect 17543 13141 17555 13144
rect 17497 13135 17555 13141
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 18782 13132 18788 13184
rect 18840 13172 18846 13184
rect 19705 13175 19763 13181
rect 19705 13172 19717 13175
rect 18840 13144 19717 13172
rect 18840 13132 18846 13144
rect 19705 13141 19717 13144
rect 19751 13141 19763 13175
rect 21082 13172 21088 13184
rect 21043 13144 21088 13172
rect 19705 13135 19763 13141
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 21450 13172 21456 13184
rect 21411 13144 21456 13172
rect 21450 13132 21456 13144
rect 21508 13132 21514 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 2961 12971 3019 12977
rect 2961 12968 2973 12971
rect 1728 12940 2973 12968
rect 1728 12928 1734 12940
rect 2961 12937 2973 12940
rect 3007 12937 3019 12971
rect 3234 12968 3240 12980
rect 3195 12940 3240 12968
rect 2961 12931 3019 12937
rect 3234 12928 3240 12940
rect 3292 12928 3298 12980
rect 3326 12928 3332 12980
rect 3384 12968 3390 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3384 12940 3525 12968
rect 3384 12928 3390 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 3513 12931 3571 12937
rect 3881 12971 3939 12977
rect 3881 12937 3893 12971
rect 3927 12968 3939 12971
rect 6362 12968 6368 12980
rect 3927 12940 6368 12968
rect 3927 12937 3939 12940
rect 3881 12931 3939 12937
rect 6362 12928 6368 12940
rect 6420 12928 6426 12980
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 7432 12940 7849 12968
rect 7432 12928 7438 12940
rect 7837 12937 7849 12940
rect 7883 12937 7895 12971
rect 8294 12968 8300 12980
rect 8207 12940 8300 12968
rect 7837 12931 7895 12937
rect 8294 12928 8300 12940
rect 8352 12968 8358 12980
rect 8662 12968 8668 12980
rect 8352 12940 8668 12968
rect 8352 12928 8358 12940
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 9122 12968 9128 12980
rect 9083 12940 9128 12968
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9490 12968 9496 12980
rect 9451 12940 9496 12968
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 9858 12968 9864 12980
rect 9732 12940 9864 12968
rect 9732 12928 9738 12940
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 9953 12971 10011 12977
rect 9953 12937 9965 12971
rect 9999 12968 10011 12971
rect 10781 12971 10839 12977
rect 10781 12968 10793 12971
rect 9999 12940 10793 12968
rect 9999 12937 10011 12940
rect 9953 12931 10011 12937
rect 10781 12937 10793 12940
rect 10827 12968 10839 12971
rect 10962 12968 10968 12980
rect 10827 12940 10968 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 10962 12928 10968 12940
rect 11020 12968 11026 12980
rect 11422 12968 11428 12980
rect 11020 12940 11428 12968
rect 11020 12928 11026 12940
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 11532 12940 11928 12968
rect 2222 12860 2228 12912
rect 2280 12900 2286 12912
rect 2624 12903 2682 12909
rect 2624 12900 2636 12903
rect 2280 12872 2636 12900
rect 2280 12860 2286 12872
rect 2624 12869 2636 12872
rect 2670 12900 2682 12903
rect 4246 12900 4252 12912
rect 2670 12872 4252 12900
rect 2670 12869 2682 12872
rect 2624 12863 2682 12869
rect 3145 12835 3203 12841
rect 3145 12801 3157 12835
rect 3191 12832 3203 12835
rect 3326 12832 3332 12844
rect 3191 12804 3332 12832
rect 3191 12801 3203 12804
rect 3145 12795 3203 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 2866 12764 2872 12776
rect 2827 12736 2872 12764
rect 2866 12724 2872 12736
rect 2924 12724 2930 12776
rect 3436 12696 3464 12795
rect 3896 12764 3924 12872
rect 4246 12860 4252 12872
rect 4304 12860 4310 12912
rect 5261 12903 5319 12909
rect 5261 12869 5273 12903
rect 5307 12900 5319 12903
rect 5626 12900 5632 12912
rect 5307 12872 5632 12900
rect 5307 12869 5319 12872
rect 5261 12863 5319 12869
rect 5626 12860 5632 12872
rect 5684 12860 5690 12912
rect 6178 12860 6184 12912
rect 6236 12900 6242 12912
rect 6236 12872 6767 12900
rect 6236 12860 6242 12872
rect 3973 12835 4031 12841
rect 3973 12801 3985 12835
rect 4019 12832 4031 12835
rect 4614 12832 4620 12844
rect 4019 12804 4620 12832
rect 4019 12801 4031 12804
rect 3973 12795 4031 12801
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12832 5227 12835
rect 5350 12832 5356 12844
rect 5215 12804 5356 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 5718 12832 5724 12844
rect 5592 12804 5724 12832
rect 5592 12792 5598 12804
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 5902 12792 5908 12844
rect 5960 12832 5966 12844
rect 6638 12841 6644 12844
rect 6089 12835 6147 12841
rect 6089 12832 6101 12835
rect 5960 12804 6101 12832
rect 5960 12792 5966 12804
rect 6089 12801 6101 12804
rect 6135 12832 6147 12835
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 6135 12804 6377 12832
rect 6135 12801 6147 12804
rect 6089 12795 6147 12801
rect 6365 12801 6377 12804
rect 6411 12801 6423 12835
rect 6632 12832 6644 12841
rect 6599 12804 6644 12832
rect 6365 12795 6423 12801
rect 6632 12795 6644 12804
rect 6638 12792 6644 12795
rect 6696 12792 6702 12844
rect 6739 12832 6767 12872
rect 7190 12860 7196 12912
rect 7248 12900 7254 12912
rect 7650 12900 7656 12912
rect 7248 12872 7656 12900
rect 7248 12860 7254 12872
rect 7650 12860 7656 12872
rect 7708 12860 7714 12912
rect 8018 12860 8024 12912
rect 8076 12900 8082 12912
rect 8205 12903 8263 12909
rect 8205 12900 8217 12903
rect 8076 12872 8217 12900
rect 8076 12860 8082 12872
rect 8205 12869 8217 12872
rect 8251 12869 8263 12903
rect 8570 12900 8576 12912
rect 8205 12863 8263 12869
rect 8292 12872 8576 12900
rect 6739 12804 7420 12832
rect 4065 12767 4123 12773
rect 4065 12764 4077 12767
rect 3896 12736 4077 12764
rect 4065 12733 4077 12736
rect 4111 12733 4123 12767
rect 4338 12764 4344 12776
rect 4299 12736 4344 12764
rect 4065 12727 4123 12733
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 5445 12767 5503 12773
rect 5445 12733 5457 12767
rect 5491 12764 5503 12767
rect 5626 12764 5632 12776
rect 5491 12736 5632 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 5626 12724 5632 12736
rect 5684 12764 5690 12776
rect 5994 12764 6000 12776
rect 5684 12736 6000 12764
rect 5684 12724 5690 12736
rect 5994 12724 6000 12736
rect 6052 12724 6058 12776
rect 7392 12764 7420 12804
rect 8292 12764 8320 12872
rect 8570 12860 8576 12872
rect 8628 12860 8634 12912
rect 9033 12903 9091 12909
rect 9033 12869 9045 12903
rect 9079 12900 9091 12903
rect 11054 12900 11060 12912
rect 9079 12872 11060 12900
rect 9079 12869 9091 12872
rect 9033 12863 9091 12869
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 11532 12900 11560 12940
rect 11164 12872 11560 12900
rect 11900 12900 11928 12940
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 12897 12971 12955 12977
rect 12897 12968 12909 12971
rect 12216 12940 12909 12968
rect 12216 12928 12222 12940
rect 12897 12937 12909 12940
rect 12943 12937 12955 12971
rect 13354 12968 13360 12980
rect 13315 12940 13360 12968
rect 12897 12931 12955 12937
rect 13354 12928 13360 12940
rect 13412 12928 13418 12980
rect 15194 12968 15200 12980
rect 15155 12940 15200 12968
rect 15194 12928 15200 12940
rect 15252 12928 15258 12980
rect 18230 12968 18236 12980
rect 18191 12940 18236 12968
rect 18230 12928 18236 12940
rect 18288 12928 18294 12980
rect 19518 12928 19524 12980
rect 19576 12968 19582 12980
rect 19797 12971 19855 12977
rect 19797 12968 19809 12971
rect 19576 12940 19809 12968
rect 19576 12928 19582 12940
rect 19797 12937 19809 12940
rect 19843 12937 19855 12971
rect 20162 12968 20168 12980
rect 20123 12940 20168 12968
rect 19797 12931 19855 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20257 12971 20315 12977
rect 20257 12937 20269 12971
rect 20303 12968 20315 12971
rect 20438 12968 20444 12980
rect 20303 12940 20444 12968
rect 20303 12937 20315 12940
rect 20257 12931 20315 12937
rect 20438 12928 20444 12940
rect 20496 12968 20502 12980
rect 20625 12971 20683 12977
rect 20625 12968 20637 12971
rect 20496 12940 20637 12968
rect 20496 12928 20502 12940
rect 20625 12937 20637 12940
rect 20671 12937 20683 12971
rect 20625 12931 20683 12937
rect 20806 12928 20812 12980
rect 20864 12928 20870 12980
rect 20990 12968 20996 12980
rect 20951 12940 20996 12968
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 12986 12900 12992 12912
rect 11900 12872 12992 12900
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 10873 12835 10931 12841
rect 10873 12832 10885 12835
rect 9916 12804 10885 12832
rect 9916 12792 9922 12804
rect 10873 12801 10885 12804
rect 10919 12832 10931 12835
rect 11164 12832 11192 12872
rect 12986 12860 12992 12872
rect 13044 12860 13050 12912
rect 14084 12903 14142 12909
rect 14084 12869 14096 12903
rect 14130 12900 14142 12903
rect 14274 12900 14280 12912
rect 14130 12872 14280 12900
rect 14130 12869 14142 12872
rect 14084 12863 14142 12869
rect 14274 12860 14280 12872
rect 14332 12860 14338 12912
rect 10919 12804 11192 12832
rect 11333 12835 11391 12841
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 11333 12801 11345 12835
rect 11379 12832 11391 12835
rect 11514 12832 11520 12844
rect 11379 12804 11520 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 11784 12835 11842 12841
rect 11784 12801 11796 12835
rect 11830 12832 11842 12835
rect 11830 12804 12572 12832
rect 11830 12801 11842 12804
rect 11784 12795 11842 12801
rect 12544 12776 12572 12804
rect 13170 12792 13176 12844
rect 13228 12792 13234 12844
rect 13725 12835 13783 12841
rect 13725 12801 13737 12835
rect 13771 12832 13783 12835
rect 13814 12832 13820 12844
rect 13771 12804 13820 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 7392 12736 8320 12764
rect 8478 12724 8484 12776
rect 8536 12764 8542 12776
rect 9214 12764 9220 12776
rect 8536 12736 8629 12764
rect 9175 12736 9220 12764
rect 8536 12724 8542 12736
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 10042 12764 10048 12776
rect 10003 12736 10048 12764
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10318 12764 10324 12776
rect 10279 12736 10324 12764
rect 10318 12724 10324 12736
rect 10376 12724 10382 12776
rect 10597 12767 10655 12773
rect 10597 12733 10609 12767
rect 10643 12764 10655 12767
rect 10778 12764 10784 12776
rect 10643 12736 10784 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 12526 12724 12532 12776
rect 12584 12724 12590 12776
rect 12802 12724 12808 12776
rect 12860 12764 12866 12776
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12860 12736 13001 12764
rect 12860 12724 12866 12736
rect 12989 12733 13001 12736
rect 13035 12764 13047 12767
rect 13188 12764 13216 12792
rect 13035 12736 13216 12764
rect 15212 12764 15240 12928
rect 15470 12860 15476 12912
rect 15528 12900 15534 12912
rect 16393 12903 16451 12909
rect 16393 12900 16405 12903
rect 15528 12872 16405 12900
rect 15528 12860 15534 12872
rect 16393 12869 16405 12872
rect 16439 12869 16451 12903
rect 18592 12903 18650 12909
rect 18592 12900 18604 12903
rect 16393 12863 16451 12869
rect 17788 12872 18604 12900
rect 15654 12832 15660 12844
rect 15615 12804 15660 12832
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 16206 12792 16212 12844
rect 16264 12832 16270 12844
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16264 12804 16865 12832
rect 16264 12792 16270 12804
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 17788 12832 17816 12872
rect 18592 12869 18604 12872
rect 18638 12900 18650 12903
rect 18966 12900 18972 12912
rect 18638 12872 18972 12900
rect 18638 12869 18650 12872
rect 18592 12863 18650 12869
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 20824 12900 20852 12928
rect 20824 12872 21036 12900
rect 21008 12844 21036 12872
rect 16853 12795 16911 12801
rect 17696 12804 17816 12832
rect 17865 12835 17923 12841
rect 17696 12773 17724 12804
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 18230 12832 18236 12844
rect 17911 12804 18236 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 18230 12792 18236 12804
rect 18288 12792 18294 12844
rect 18322 12792 18328 12844
rect 18380 12832 18386 12844
rect 18380 12804 18425 12832
rect 18380 12792 18386 12804
rect 18874 12792 18880 12844
rect 18932 12832 18938 12844
rect 20806 12832 20812 12844
rect 18932 12804 20392 12832
rect 20767 12804 20812 12832
rect 18932 12792 18938 12804
rect 15381 12767 15439 12773
rect 15381 12764 15393 12767
rect 15212 12736 15393 12764
rect 13035 12733 13047 12736
rect 12989 12727 13047 12733
rect 15381 12733 15393 12736
rect 15427 12733 15439 12767
rect 15381 12727 15439 12733
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12733 15623 12767
rect 17681 12767 17739 12773
rect 15565 12727 15623 12733
rect 16040 12736 17632 12764
rect 4246 12696 4252 12708
rect 3436 12668 4252 12696
rect 4246 12656 4252 12668
rect 4304 12656 4310 12708
rect 4706 12656 4712 12708
rect 4764 12696 4770 12708
rect 4801 12699 4859 12705
rect 4801 12696 4813 12699
rect 4764 12668 4813 12696
rect 4764 12656 4770 12668
rect 4801 12665 4813 12668
rect 4847 12665 4859 12699
rect 4801 12659 4859 12665
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 5905 12699 5963 12705
rect 5905 12696 5917 12699
rect 4948 12668 5917 12696
rect 4948 12656 4954 12668
rect 5905 12665 5917 12668
rect 5951 12665 5963 12699
rect 5905 12659 5963 12665
rect 7745 12699 7803 12705
rect 7745 12665 7757 12699
rect 7791 12696 7803 12699
rect 8496 12696 8524 12724
rect 7791 12668 8524 12696
rect 7791 12665 7803 12668
rect 7745 12659 7803 12665
rect 8570 12656 8576 12708
rect 8628 12696 8634 12708
rect 13173 12699 13231 12705
rect 13173 12696 13185 12699
rect 8628 12668 11284 12696
rect 8628 12656 8634 12668
rect 1489 12631 1547 12637
rect 1489 12597 1501 12631
rect 1535 12628 1547 12631
rect 2498 12628 2504 12640
rect 1535 12600 2504 12628
rect 1535 12597 1547 12600
rect 1489 12591 1547 12597
rect 2498 12588 2504 12600
rect 2556 12588 2562 12640
rect 3786 12588 3792 12640
rect 3844 12628 3850 12640
rect 3970 12628 3976 12640
rect 3844 12600 3976 12628
rect 3844 12588 3850 12600
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 4617 12631 4675 12637
rect 4617 12597 4629 12631
rect 4663 12628 4675 12631
rect 4982 12628 4988 12640
rect 4663 12600 4988 12628
rect 4663 12597 4675 12600
rect 4617 12591 4675 12597
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 5813 12631 5871 12637
rect 5813 12628 5825 12631
rect 5408 12600 5825 12628
rect 5408 12588 5414 12600
rect 5813 12597 5825 12600
rect 5859 12628 5871 12631
rect 6270 12628 6276 12640
rect 5859 12600 6276 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 6270 12588 6276 12600
rect 6328 12588 6334 12640
rect 6362 12588 6368 12640
rect 6420 12628 6426 12640
rect 8665 12631 8723 12637
rect 8665 12628 8677 12631
rect 6420 12600 8677 12628
rect 6420 12588 6426 12600
rect 8665 12597 8677 12600
rect 8711 12597 8723 12631
rect 8665 12591 8723 12597
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 10870 12628 10876 12640
rect 9180 12600 10876 12628
rect 9180 12588 9186 12600
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 11149 12631 11207 12637
rect 11149 12628 11161 12631
rect 11112 12600 11161 12628
rect 11112 12588 11118 12600
rect 11149 12597 11161 12600
rect 11195 12597 11207 12631
rect 11256 12628 11284 12668
rect 12820 12668 13185 12696
rect 12820 12628 12848 12668
rect 13173 12665 13185 12668
rect 13219 12665 13231 12699
rect 13541 12699 13599 12705
rect 13541 12696 13553 12699
rect 13173 12659 13231 12665
rect 13280 12668 13553 12696
rect 11256 12600 12848 12628
rect 11149 12591 11207 12597
rect 13078 12588 13084 12640
rect 13136 12628 13142 12640
rect 13280 12628 13308 12668
rect 13541 12665 13553 12668
rect 13587 12665 13599 12699
rect 13541 12659 13599 12665
rect 15102 12656 15108 12708
rect 15160 12696 15166 12708
rect 15580 12696 15608 12727
rect 16040 12705 16068 12736
rect 15160 12668 15608 12696
rect 16025 12699 16083 12705
rect 15160 12656 15166 12668
rect 16025 12665 16037 12699
rect 16071 12665 16083 12699
rect 16025 12659 16083 12665
rect 16301 12699 16359 12705
rect 16301 12665 16313 12699
rect 16347 12696 16359 12699
rect 16574 12696 16580 12708
rect 16347 12668 16580 12696
rect 16347 12665 16359 12668
rect 16301 12659 16359 12665
rect 16574 12656 16580 12668
rect 16632 12656 16638 12708
rect 16758 12628 16764 12640
rect 13136 12600 13308 12628
rect 16719 12600 16764 12628
rect 13136 12588 13142 12600
rect 16758 12588 16764 12600
rect 16816 12588 16822 12640
rect 17034 12628 17040 12640
rect 16995 12600 17040 12628
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 17402 12628 17408 12640
rect 17363 12600 17408 12628
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 17604 12628 17632 12736
rect 17681 12733 17693 12767
rect 17727 12733 17739 12767
rect 17681 12727 17739 12733
rect 17773 12767 17831 12773
rect 17773 12733 17785 12767
rect 17819 12764 17831 12767
rect 18046 12764 18052 12776
rect 17819 12736 18052 12764
rect 17819 12733 17831 12736
rect 17773 12727 17831 12733
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 20364 12773 20392 12804
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 20990 12792 20996 12844
rect 21048 12792 21054 12844
rect 21266 12832 21272 12844
rect 21227 12804 21272 12832
rect 21266 12792 21272 12804
rect 21324 12792 21330 12844
rect 20349 12767 20407 12773
rect 20349 12733 20361 12767
rect 20395 12733 20407 12767
rect 20349 12727 20407 12733
rect 19518 12656 19524 12708
rect 19576 12696 19582 12708
rect 19705 12699 19763 12705
rect 19705 12696 19717 12699
rect 19576 12668 19717 12696
rect 19576 12656 19582 12668
rect 19705 12665 19717 12668
rect 19751 12696 19763 12699
rect 20530 12696 20536 12708
rect 19751 12668 20536 12696
rect 19751 12665 19763 12668
rect 19705 12659 19763 12665
rect 20530 12656 20536 12668
rect 20588 12656 20594 12708
rect 21177 12699 21235 12705
rect 21177 12665 21189 12699
rect 21223 12696 21235 12699
rect 21542 12696 21548 12708
rect 21223 12668 21548 12696
rect 21223 12665 21235 12668
rect 21177 12659 21235 12665
rect 21542 12656 21548 12668
rect 21600 12656 21606 12708
rect 20438 12628 20444 12640
rect 17604 12600 20444 12628
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 21450 12628 21456 12640
rect 21411 12600 21456 12628
rect 21450 12588 21456 12600
rect 21508 12588 21514 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 1486 12424 1492 12436
rect 1447 12396 1492 12424
rect 1486 12384 1492 12396
rect 1544 12384 1550 12436
rect 3970 12424 3976 12436
rect 3931 12396 3976 12424
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4246 12384 4252 12436
rect 4304 12424 4310 12436
rect 6273 12427 6331 12433
rect 6273 12424 6285 12427
rect 4304 12396 6285 12424
rect 4304 12384 4310 12396
rect 6273 12393 6285 12396
rect 6319 12393 6331 12427
rect 6273 12387 6331 12393
rect 6362 12384 6368 12436
rect 6420 12424 6426 12436
rect 7374 12424 7380 12436
rect 6420 12396 7380 12424
rect 6420 12384 6426 12396
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 7926 12384 7932 12436
rect 7984 12424 7990 12436
rect 8294 12424 8300 12436
rect 7984 12396 8300 12424
rect 7984 12384 7990 12396
rect 8294 12384 8300 12396
rect 8352 12424 8358 12436
rect 8665 12427 8723 12433
rect 8665 12424 8677 12427
rect 8352 12396 8677 12424
rect 8352 12384 8358 12396
rect 8665 12393 8677 12396
rect 8711 12393 8723 12427
rect 8665 12387 8723 12393
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 8812 12396 8953 12424
rect 8812 12384 8818 12396
rect 8941 12393 8953 12396
rect 8987 12393 8999 12427
rect 9490 12424 9496 12436
rect 9451 12396 9496 12424
rect 8941 12387 8999 12393
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 10594 12424 10600 12436
rect 10555 12396 10600 12424
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 10962 12384 10968 12436
rect 11020 12424 11026 12436
rect 11238 12424 11244 12436
rect 11020 12396 11244 12424
rect 11020 12384 11026 12396
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12250 12424 12256 12436
rect 12032 12396 12256 12424
rect 12032 12384 12038 12396
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 13449 12427 13507 12433
rect 13449 12393 13461 12427
rect 13495 12424 13507 12427
rect 13538 12424 13544 12436
rect 13495 12396 13544 12424
rect 13495 12393 13507 12396
rect 13449 12387 13507 12393
rect 3234 12316 3240 12368
rect 3292 12356 3298 12368
rect 4154 12356 4160 12368
rect 3292 12328 4160 12356
rect 3292 12316 3298 12328
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 6181 12359 6239 12365
rect 6181 12325 6193 12359
rect 6227 12356 6239 12359
rect 6638 12356 6644 12368
rect 6227 12328 6644 12356
rect 6227 12325 6239 12328
rect 6181 12319 6239 12325
rect 6638 12316 6644 12328
rect 6696 12356 6702 12368
rect 6696 12328 6868 12356
rect 6696 12316 6702 12328
rect 3326 12248 3332 12300
rect 3384 12288 3390 12300
rect 3694 12288 3700 12300
rect 3384 12260 3700 12288
rect 3384 12248 3390 12260
rect 3694 12248 3700 12260
rect 3752 12288 3758 12300
rect 3789 12291 3847 12297
rect 3789 12288 3801 12291
rect 3752 12260 3801 12288
rect 3752 12248 3758 12260
rect 3789 12257 3801 12260
rect 3835 12257 3847 12291
rect 3789 12251 3847 12257
rect 3878 12248 3884 12300
rect 3936 12288 3942 12300
rect 4522 12288 4528 12300
rect 3936 12260 4528 12288
rect 3936 12248 3942 12260
rect 4522 12248 4528 12260
rect 4580 12248 4586 12300
rect 6840 12297 6868 12328
rect 7282 12316 7288 12368
rect 7340 12356 7346 12368
rect 8021 12359 8079 12365
rect 8021 12356 8033 12359
rect 7340 12328 8033 12356
rect 7340 12316 7346 12328
rect 8021 12325 8033 12328
rect 8067 12325 8079 12359
rect 8021 12319 8079 12325
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 9214 12356 9220 12368
rect 8260 12328 9220 12356
rect 8260 12316 8266 12328
rect 9214 12316 9220 12328
rect 9272 12316 9278 12368
rect 9309 12359 9367 12365
rect 9309 12325 9321 12359
rect 9355 12356 9367 12359
rect 9766 12356 9772 12368
rect 9355 12328 9772 12356
rect 9355 12325 9367 12328
rect 9309 12319 9367 12325
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 9858 12316 9864 12368
rect 9916 12356 9922 12368
rect 10689 12359 10747 12365
rect 10689 12356 10701 12359
rect 9916 12328 10701 12356
rect 9916 12316 9922 12328
rect 10689 12325 10701 12328
rect 10735 12325 10747 12359
rect 10689 12319 10747 12325
rect 12526 12316 12532 12368
rect 12584 12356 12590 12368
rect 12894 12356 12900 12368
rect 12584 12328 12900 12356
rect 12584 12316 12590 12328
rect 12894 12316 12900 12328
rect 12952 12316 12958 12368
rect 12986 12316 12992 12368
rect 13044 12356 13050 12368
rect 13354 12356 13360 12368
rect 13044 12328 13360 12356
rect 13044 12316 13050 12328
rect 13354 12316 13360 12328
rect 13412 12316 13418 12368
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12257 6883 12291
rect 7098 12288 7104 12300
rect 7059 12260 7104 12288
rect 6825 12251 6883 12257
rect 7098 12248 7104 12260
rect 7156 12248 7162 12300
rect 7377 12291 7435 12297
rect 7377 12257 7389 12291
rect 7423 12288 7435 12291
rect 7742 12288 7748 12300
rect 7423 12260 7748 12288
rect 7423 12257 7435 12260
rect 7377 12251 7435 12257
rect 7742 12248 7748 12260
rect 7800 12288 7806 12300
rect 10778 12288 10784 12300
rect 7800 12260 10784 12288
rect 7800 12248 7806 12260
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11054 12288 11060 12300
rect 11015 12260 11060 12288
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 12434 12288 12440 12300
rect 12347 12260 12440 12288
rect 12434 12248 12440 12260
rect 12492 12288 12498 12300
rect 13081 12291 13139 12297
rect 13081 12288 13093 12291
rect 12492 12260 13093 12288
rect 12492 12248 12498 12260
rect 13081 12257 13093 12260
rect 13127 12288 13139 12291
rect 13170 12288 13176 12300
rect 13127 12260 13176 12288
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 1946 12220 1952 12232
rect 1719 12192 1952 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 1946 12180 1952 12192
rect 2004 12180 2010 12232
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12220 2099 12223
rect 2130 12220 2136 12232
rect 2087 12192 2136 12220
rect 2087 12189 2099 12192
rect 2041 12183 2099 12189
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 2498 12229 2504 12232
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 2492 12183 2504 12229
rect 2556 12220 2562 12232
rect 2866 12220 2872 12232
rect 2556 12192 2592 12220
rect 2746 12192 2872 12220
rect 1486 12112 1492 12164
rect 1544 12152 1550 12164
rect 2240 12152 2268 12183
rect 2498 12180 2504 12183
rect 2556 12180 2562 12192
rect 2746 12152 2774 12192
rect 2866 12180 2872 12192
rect 2924 12220 2930 12232
rect 4062 12220 4068 12232
rect 2924 12192 4068 12220
rect 2924 12180 2930 12192
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 4706 12220 4712 12232
rect 4479 12192 4712 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12220 4859 12223
rect 4890 12220 4896 12232
rect 4847 12192 4896 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 7469 12223 7527 12229
rect 7469 12220 7481 12223
rect 4991 12192 7481 12220
rect 4991 12152 5019 12192
rect 7469 12189 7481 12192
rect 7515 12189 7527 12223
rect 7469 12183 7527 12189
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 8846 12220 8852 12232
rect 7708 12192 8852 12220
rect 7708 12180 7714 12192
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12220 9183 12223
rect 9214 12220 9220 12232
rect 9171 12192 9220 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 9214 12180 9220 12192
rect 9272 12220 9278 12232
rect 11072 12220 11100 12248
rect 12342 12220 12348 12232
rect 9272 12192 11100 12220
rect 11164 12192 12348 12220
rect 9272 12180 9278 12192
rect 1544 12124 1992 12152
rect 2240 12124 2774 12152
rect 2884 12124 5019 12152
rect 5068 12155 5126 12161
rect 1544 12112 1550 12124
rect 1854 12084 1860 12096
rect 1815 12056 1860 12084
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 1964 12084 1992 12124
rect 2884 12084 2912 12124
rect 5068 12121 5080 12155
rect 5114 12152 5126 12155
rect 5114 12124 5304 12152
rect 5114 12121 5126 12124
rect 5068 12115 5126 12121
rect 1964 12056 2912 12084
rect 3605 12087 3663 12093
rect 3605 12053 3617 12087
rect 3651 12084 3663 12087
rect 4154 12084 4160 12096
rect 3651 12056 4160 12084
rect 3651 12053 3663 12056
rect 3605 12047 3663 12053
rect 4154 12044 4160 12056
rect 4212 12044 4218 12096
rect 4341 12087 4399 12093
rect 4341 12053 4353 12087
rect 4387 12084 4399 12087
rect 4890 12084 4896 12096
rect 4387 12056 4896 12084
rect 4387 12053 4399 12056
rect 4341 12047 4399 12053
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 5276 12084 5304 12124
rect 5350 12112 5356 12164
rect 5408 12152 5414 12164
rect 6641 12155 6699 12161
rect 6641 12152 6653 12155
rect 5408 12124 6653 12152
rect 5408 12112 5414 12124
rect 6641 12121 6653 12124
rect 6687 12121 6699 12155
rect 6641 12115 6699 12121
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 8294 12152 8300 12164
rect 6972 12124 8300 12152
rect 6972 12112 6978 12124
rect 8294 12112 8300 12124
rect 8352 12152 8358 12164
rect 11164 12152 11192 12192
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 11330 12161 11336 12164
rect 8352 12124 11192 12152
rect 8352 12112 8358 12124
rect 11324 12115 11336 12161
rect 11388 12152 11394 12164
rect 11388 12124 11424 12152
rect 11330 12112 11336 12115
rect 11388 12112 11394 12124
rect 11790 12112 11796 12164
rect 11848 12152 11854 12164
rect 12452 12152 12480 12248
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12220 12955 12223
rect 13464 12220 13492 12387
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 14093 12427 14151 12433
rect 14093 12393 14105 12427
rect 14139 12424 14151 12427
rect 14274 12424 14280 12436
rect 14139 12396 14280 12424
rect 14139 12393 14151 12396
rect 14093 12387 14151 12393
rect 14274 12384 14280 12396
rect 14332 12424 14338 12436
rect 15565 12427 15623 12433
rect 14332 12396 15516 12424
rect 14332 12384 14338 12396
rect 15488 12356 15516 12396
rect 15565 12393 15577 12427
rect 15611 12424 15623 12427
rect 15654 12424 15660 12436
rect 15611 12396 15660 12424
rect 15611 12393 15623 12396
rect 15565 12387 15623 12393
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 16390 12424 16396 12436
rect 16351 12396 16396 12424
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 18046 12424 18052 12436
rect 18007 12396 18052 12424
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 19429 12427 19487 12433
rect 19429 12393 19441 12427
rect 19475 12424 19487 12427
rect 20622 12424 20628 12436
rect 19475 12396 20628 12424
rect 19475 12393 19487 12396
rect 19429 12387 19487 12393
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 20717 12427 20775 12433
rect 20717 12393 20729 12427
rect 20763 12424 20775 12427
rect 20806 12424 20812 12436
rect 20763 12396 20812 12424
rect 20763 12393 20775 12396
rect 20717 12387 20775 12393
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 22278 12384 22284 12436
rect 22336 12424 22342 12436
rect 22336 12396 22600 12424
rect 22336 12384 22342 12396
rect 22572 12368 22600 12396
rect 17954 12356 17960 12368
rect 15488 12328 16160 12356
rect 16132 12297 16160 12328
rect 17420 12328 17960 12356
rect 16117 12291 16175 12297
rect 16117 12257 16129 12291
rect 16163 12257 16175 12291
rect 16942 12288 16948 12300
rect 16903 12260 16948 12288
rect 16117 12251 16175 12257
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 17420 12297 17448 12328
rect 17954 12316 17960 12328
rect 18012 12316 18018 12368
rect 20254 12316 20260 12368
rect 20312 12356 20318 12368
rect 20901 12359 20959 12365
rect 20901 12356 20913 12359
rect 20312 12328 20913 12356
rect 20312 12316 20318 12328
rect 20901 12325 20913 12328
rect 20947 12325 20959 12359
rect 20901 12319 20959 12325
rect 22554 12316 22560 12368
rect 22612 12316 22618 12368
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12257 17463 12291
rect 17405 12251 17463 12257
rect 17586 12248 17592 12300
rect 17644 12288 17650 12300
rect 18601 12291 18659 12297
rect 18601 12288 18613 12291
rect 17644 12260 18613 12288
rect 17644 12248 17650 12260
rect 18601 12257 18613 12260
rect 18647 12257 18659 12291
rect 18601 12251 18659 12257
rect 19705 12291 19763 12297
rect 19705 12257 19717 12291
rect 19751 12288 19763 12291
rect 20346 12288 20352 12300
rect 19751 12260 20352 12288
rect 19751 12257 19763 12260
rect 19705 12251 19763 12257
rect 20346 12248 20352 12260
rect 20404 12248 20410 12300
rect 22094 12248 22100 12300
rect 22152 12288 22158 12300
rect 22370 12288 22376 12300
rect 22152 12260 22376 12288
rect 22152 12248 22158 12260
rect 22370 12248 22376 12260
rect 22428 12248 22434 12300
rect 12943 12192 13492 12220
rect 12943 12189 12955 12192
rect 12897 12183 12955 12189
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14826 12220 14832 12232
rect 13872 12192 14832 12220
rect 13872 12180 13878 12192
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 15378 12180 15384 12232
rect 15436 12220 15442 12232
rect 15473 12223 15531 12229
rect 15473 12220 15485 12223
rect 15436 12192 15485 12220
rect 15436 12180 15442 12192
rect 15473 12189 15485 12192
rect 15519 12189 15531 12223
rect 15473 12183 15531 12189
rect 16206 12180 16212 12232
rect 16264 12220 16270 12232
rect 17497 12223 17555 12229
rect 17497 12220 17509 12223
rect 16264 12192 17509 12220
rect 16264 12180 16270 12192
rect 17497 12189 17509 12192
rect 17543 12189 17555 12223
rect 18874 12220 18880 12232
rect 18835 12192 18880 12220
rect 17497 12183 17555 12189
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 20530 12220 20536 12232
rect 19291 12192 20392 12220
rect 20491 12192 20536 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 11848 12124 12480 12152
rect 11848 12112 11854 12124
rect 5626 12084 5632 12096
rect 5276 12056 5632 12084
rect 5626 12044 5632 12056
rect 5684 12044 5690 12096
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 6788 12056 6833 12084
rect 6788 12044 6794 12056
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 7653 12087 7711 12093
rect 7653 12084 7665 12087
rect 7064 12056 7665 12084
rect 7064 12044 7070 12056
rect 7653 12053 7665 12056
rect 7699 12053 7711 12087
rect 7653 12047 7711 12053
rect 7929 12087 7987 12093
rect 7929 12053 7941 12087
rect 7975 12084 7987 12087
rect 8018 12084 8024 12096
rect 7975 12056 8024 12084
rect 7975 12053 7987 12056
rect 7929 12047 7987 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8202 12084 8208 12096
rect 8163 12056 8208 12084
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 8481 12087 8539 12093
rect 8481 12053 8493 12087
rect 8527 12084 8539 12087
rect 8570 12084 8576 12096
rect 8527 12056 8576 12084
rect 8527 12053 8539 12056
rect 8481 12047 8539 12053
rect 8570 12044 8576 12056
rect 8628 12044 8634 12096
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 9585 12087 9643 12093
rect 9585 12084 9597 12087
rect 8720 12056 9597 12084
rect 8720 12044 8726 12056
rect 9585 12053 9597 12056
rect 9631 12053 9643 12087
rect 9858 12084 9864 12096
rect 9819 12056 9864 12084
rect 9585 12047 9643 12053
rect 9858 12044 9864 12056
rect 9916 12044 9922 12096
rect 10042 12084 10048 12096
rect 10003 12056 10048 12084
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 10226 12084 10232 12096
rect 10187 12056 10232 12084
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 10376 12056 10421 12084
rect 10376 12044 10382 12056
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 12452 12093 12480 12124
rect 13446 12112 13452 12164
rect 13504 12152 13510 12164
rect 14642 12152 14648 12164
rect 13504 12124 14648 12152
rect 13504 12112 13510 12124
rect 14642 12112 14648 12124
rect 14700 12112 14706 12164
rect 15206 12155 15264 12161
rect 15206 12121 15218 12155
rect 15252 12121 15264 12155
rect 16114 12152 16120 12164
rect 15206 12115 15264 12121
rect 15396 12124 16120 12152
rect 10873 12087 10931 12093
rect 10873 12084 10885 12087
rect 10836 12056 10885 12084
rect 10836 12044 10842 12056
rect 10873 12053 10885 12056
rect 10919 12053 10931 12087
rect 10873 12047 10931 12053
rect 12437 12087 12495 12093
rect 12437 12053 12449 12087
rect 12483 12053 12495 12087
rect 12437 12047 12495 12053
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12584 12056 12629 12084
rect 12584 12044 12590 12056
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 12989 12087 13047 12093
rect 12989 12084 13001 12087
rect 12952 12056 13001 12084
rect 12952 12044 12958 12056
rect 12989 12053 13001 12056
rect 13035 12053 13047 12087
rect 12989 12047 13047 12053
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 13541 12087 13599 12093
rect 13541 12084 13553 12087
rect 13136 12056 13553 12084
rect 13136 12044 13142 12056
rect 13541 12053 13553 12056
rect 13587 12053 13599 12087
rect 13814 12084 13820 12096
rect 13775 12056 13820 12084
rect 13541 12047 13599 12053
rect 13814 12044 13820 12056
rect 13872 12044 13878 12096
rect 15212 12084 15240 12115
rect 15396 12096 15424 12124
rect 16114 12112 16120 12124
rect 16172 12112 16178 12164
rect 16758 12152 16764 12164
rect 16719 12124 16764 12152
rect 16758 12112 16764 12124
rect 16816 12112 16822 12164
rect 17034 12112 17040 12164
rect 17092 12152 17098 12164
rect 17589 12155 17647 12161
rect 17589 12152 17601 12155
rect 17092 12124 17601 12152
rect 17092 12112 17098 12124
rect 17589 12121 17601 12124
rect 17635 12121 17647 12155
rect 18509 12155 18567 12161
rect 18509 12152 18521 12155
rect 17589 12115 17647 12121
rect 17972 12124 18521 12152
rect 15286 12084 15292 12096
rect 15212 12056 15292 12084
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 15378 12044 15384 12096
rect 15436 12044 15442 12096
rect 15930 12084 15936 12096
rect 15891 12056 15936 12084
rect 15930 12044 15936 12056
rect 15988 12044 15994 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16853 12087 16911 12093
rect 16080 12056 16125 12084
rect 16080 12044 16086 12056
rect 16853 12053 16865 12087
rect 16899 12084 16911 12087
rect 17218 12084 17224 12096
rect 16899 12056 17224 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 17972 12093 18000 12124
rect 18509 12121 18521 12124
rect 18555 12121 18567 12155
rect 18509 12115 18567 12121
rect 19797 12155 19855 12161
rect 19797 12121 19809 12155
rect 19843 12152 19855 12155
rect 20162 12152 20168 12164
rect 19843 12124 20168 12152
rect 19843 12121 19855 12124
rect 19797 12115 19855 12121
rect 20162 12112 20168 12124
rect 20220 12112 20226 12164
rect 20364 12152 20392 12192
rect 20530 12180 20536 12192
rect 20588 12180 20594 12232
rect 21269 12223 21327 12229
rect 21269 12189 21281 12223
rect 21315 12220 21327 12223
rect 21634 12220 21640 12232
rect 21315 12192 21640 12220
rect 21315 12189 21327 12192
rect 21269 12183 21327 12189
rect 21634 12180 21640 12192
rect 21692 12180 21698 12232
rect 20438 12152 20444 12164
rect 20364 12124 20444 12152
rect 20438 12112 20444 12124
rect 20496 12112 20502 12164
rect 21082 12152 21088 12164
rect 20916 12124 21088 12152
rect 17957 12087 18015 12093
rect 17957 12053 17969 12087
rect 18003 12053 18015 12087
rect 18414 12084 18420 12096
rect 18375 12056 18420 12084
rect 17957 12047 18015 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 19061 12087 19119 12093
rect 19061 12053 19073 12087
rect 19107 12084 19119 12087
rect 19334 12084 19340 12096
rect 19107 12056 19340 12084
rect 19107 12053 19119 12056
rect 19061 12047 19119 12053
rect 19334 12044 19340 12056
rect 19392 12044 19398 12096
rect 19886 12044 19892 12096
rect 19944 12084 19950 12096
rect 20254 12084 20260 12096
rect 19944 12056 19989 12084
rect 20215 12056 20260 12084
rect 19944 12044 19950 12056
rect 20254 12044 20260 12056
rect 20312 12044 20318 12096
rect 20349 12087 20407 12093
rect 20349 12053 20361 12087
rect 20395 12084 20407 12087
rect 20916 12084 20944 12124
rect 21082 12112 21088 12124
rect 21140 12112 21146 12164
rect 21450 12084 21456 12096
rect 20395 12056 20944 12084
rect 21411 12056 21456 12084
rect 20395 12053 20407 12056
rect 20349 12047 20407 12053
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 2314 11880 2320 11892
rect 1964 11852 2320 11880
rect 1964 11753 1992 11852
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 2682 11880 2688 11892
rect 2464 11852 2688 11880
rect 2464 11840 2470 11852
rect 2682 11840 2688 11852
rect 2740 11840 2746 11892
rect 3237 11883 3295 11889
rect 3237 11849 3249 11883
rect 3283 11880 3295 11883
rect 3418 11880 3424 11892
rect 3283 11852 3424 11880
rect 3283 11849 3295 11852
rect 3237 11843 3295 11849
rect 3418 11840 3424 11852
rect 3476 11840 3482 11892
rect 3605 11883 3663 11889
rect 3605 11849 3617 11883
rect 3651 11880 3663 11883
rect 4338 11880 4344 11892
rect 3651 11852 4344 11880
rect 3651 11849 3663 11852
rect 3605 11843 3663 11849
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 5350 11880 5356 11892
rect 5311 11852 5356 11880
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 5767 11852 6469 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 7190 11880 7196 11892
rect 6457 11843 6515 11849
rect 6748 11852 7196 11880
rect 2774 11812 2780 11824
rect 2240 11784 2780 11812
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11713 2007 11747
rect 1949 11707 2007 11713
rect 2240 11688 2268 11784
rect 2774 11772 2780 11784
rect 2832 11772 2838 11824
rect 2866 11772 2872 11824
rect 2924 11812 2930 11824
rect 3697 11815 3755 11821
rect 3697 11812 3709 11815
rect 2924 11784 3709 11812
rect 2924 11772 2930 11784
rect 3697 11781 3709 11784
rect 3743 11781 3755 11815
rect 3697 11775 3755 11781
rect 4798 11772 4804 11824
rect 4856 11772 4862 11824
rect 4893 11815 4951 11821
rect 4893 11781 4905 11815
rect 4939 11812 4951 11815
rect 5534 11812 5540 11824
rect 4939 11784 5540 11812
rect 4939 11781 4951 11784
rect 4893 11775 4951 11781
rect 5534 11772 5540 11784
rect 5592 11772 5598 11824
rect 6178 11772 6184 11824
rect 6236 11812 6242 11824
rect 6748 11812 6776 11852
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7742 11880 7748 11892
rect 7361 11852 7512 11880
rect 7703 11852 7748 11880
rect 6236 11784 6776 11812
rect 6825 11815 6883 11821
rect 6236 11772 6242 11784
rect 6825 11781 6837 11815
rect 6871 11812 6883 11815
rect 7361 11812 7389 11852
rect 6871 11784 7389 11812
rect 6871 11781 6883 11784
rect 6825 11775 6883 11781
rect 2406 11704 2412 11756
rect 2464 11744 2470 11756
rect 2685 11747 2743 11753
rect 2685 11744 2697 11747
rect 2464 11716 2697 11744
rect 2464 11704 2470 11716
rect 2685 11713 2697 11716
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 3418 11704 3424 11756
rect 3476 11744 3482 11756
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 3476 11716 4261 11744
rect 3476 11704 3482 11716
rect 4249 11713 4261 11716
rect 4295 11744 4307 11747
rect 4522 11744 4528 11756
rect 4295 11716 4384 11744
rect 4435 11716 4528 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 2222 11676 2228 11688
rect 2183 11648 2228 11676
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 2961 11679 3019 11685
rect 2832 11648 2877 11676
rect 2832 11636 2838 11648
rect 2961 11645 2973 11679
rect 3007 11645 3019 11679
rect 3878 11676 3884 11688
rect 3839 11648 3884 11676
rect 2961 11639 3019 11645
rect 1854 11568 1860 11620
rect 1912 11608 1918 11620
rect 1912 11580 2452 11608
rect 1912 11568 1918 11580
rect 1394 11500 1400 11552
rect 1452 11540 1458 11552
rect 2317 11543 2375 11549
rect 2317 11540 2329 11543
rect 1452 11512 2329 11540
rect 1452 11500 1458 11512
rect 2317 11509 2329 11512
rect 2363 11509 2375 11543
rect 2424 11540 2452 11580
rect 2498 11568 2504 11620
rect 2556 11608 2562 11620
rect 2976 11608 3004 11639
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 4062 11608 4068 11620
rect 2556 11580 3004 11608
rect 4023 11580 4068 11608
rect 2556 11568 2562 11580
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 4356 11617 4384 11716
rect 4522 11704 4528 11716
rect 4580 11744 4586 11756
rect 4816 11744 4844 11772
rect 4982 11744 4988 11756
rect 4580 11716 4844 11744
rect 4943 11716 4988 11744
rect 4580 11704 4586 11716
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 5810 11744 5816 11756
rect 5771 11716 5816 11744
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 7484 11744 7512 11852
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 8113 11883 8171 11889
rect 8113 11880 8125 11883
rect 7852 11852 8125 11880
rect 7650 11772 7656 11824
rect 7708 11812 7714 11824
rect 7708 11784 7753 11812
rect 7708 11772 7714 11784
rect 7852 11744 7880 11852
rect 8113 11849 8125 11852
rect 8159 11849 8171 11883
rect 8113 11843 8171 11849
rect 8573 11883 8631 11889
rect 8573 11849 8585 11883
rect 8619 11880 8631 11883
rect 9030 11880 9036 11892
rect 8619 11852 9036 11880
rect 8619 11849 8631 11852
rect 8573 11843 8631 11849
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 9140 11852 11192 11880
rect 8481 11815 8539 11821
rect 8481 11781 8493 11815
rect 8527 11812 8539 11815
rect 8938 11812 8944 11824
rect 8527 11784 8944 11812
rect 8527 11781 8539 11784
rect 8481 11775 8539 11781
rect 8938 11772 8944 11784
rect 8996 11772 9002 11824
rect 7484 11716 7880 11744
rect 8018 11704 8024 11756
rect 8076 11744 8082 11756
rect 9140 11744 9168 11852
rect 9306 11772 9312 11824
rect 9364 11812 9370 11824
rect 9401 11815 9459 11821
rect 9401 11812 9413 11815
rect 9364 11784 9413 11812
rect 9364 11772 9370 11784
rect 9401 11781 9413 11784
rect 9447 11781 9459 11815
rect 11054 11812 11060 11824
rect 9401 11775 9459 11781
rect 9968 11784 11060 11812
rect 8076 11716 9168 11744
rect 9493 11747 9551 11753
rect 8076 11704 8082 11716
rect 9493 11713 9505 11747
rect 9539 11744 9551 11747
rect 9766 11744 9772 11756
rect 9539 11716 9772 11744
rect 9539 11713 9551 11716
rect 9493 11707 9551 11713
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 9968 11753 9996 11784
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10220 11747 10278 11753
rect 10220 11713 10232 11747
rect 10266 11744 10278 11747
rect 10502 11744 10508 11756
rect 10266 11716 10508 11744
rect 10266 11713 10278 11716
rect 10220 11707 10278 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 11164 11744 11192 11852
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11333 11883 11391 11889
rect 11333 11880 11345 11883
rect 11296 11852 11345 11880
rect 11296 11840 11302 11852
rect 11333 11849 11345 11852
rect 11379 11849 11391 11883
rect 11333 11843 11391 11849
rect 12161 11883 12219 11889
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 12526 11880 12532 11892
rect 12207 11852 12532 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 12526 11840 12532 11852
rect 12584 11840 12590 11892
rect 12618 11840 12624 11892
rect 12676 11880 12682 11892
rect 12986 11880 12992 11892
rect 12676 11852 12992 11880
rect 12676 11840 12682 11852
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 13449 11883 13507 11889
rect 13449 11849 13461 11883
rect 13495 11880 13507 11883
rect 13909 11883 13967 11889
rect 13909 11880 13921 11883
rect 13495 11852 13921 11880
rect 13495 11849 13507 11852
rect 13449 11843 13507 11849
rect 13909 11849 13921 11852
rect 13955 11849 13967 11883
rect 15102 11880 15108 11892
rect 15063 11852 15108 11880
rect 13909 11843 13967 11849
rect 15102 11840 15108 11852
rect 15160 11840 15166 11892
rect 16022 11840 16028 11892
rect 16080 11880 16086 11892
rect 16669 11883 16727 11889
rect 16669 11880 16681 11883
rect 16080 11852 16681 11880
rect 16080 11840 16086 11852
rect 16669 11849 16681 11852
rect 16715 11849 16727 11883
rect 16669 11843 16727 11849
rect 17037 11883 17095 11889
rect 17037 11849 17049 11883
rect 17083 11880 17095 11883
rect 17126 11880 17132 11892
rect 17083 11852 17132 11880
rect 17083 11849 17095 11852
rect 17037 11843 17095 11849
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 17402 11840 17408 11892
rect 17460 11880 17466 11892
rect 17865 11883 17923 11889
rect 17865 11880 17877 11883
rect 17460 11852 17877 11880
rect 17460 11840 17466 11852
rect 17865 11849 17877 11852
rect 17911 11849 17923 11883
rect 18230 11880 18236 11892
rect 18191 11852 18236 11880
rect 17865 11843 17923 11849
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 20346 11880 20352 11892
rect 20307 11852 20352 11880
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 20496 11852 20541 11880
rect 20496 11840 20502 11852
rect 22830 11840 22836 11892
rect 22888 11840 22894 11892
rect 11422 11772 11428 11824
rect 11480 11812 11486 11824
rect 12894 11812 12900 11824
rect 11480 11784 12900 11812
rect 11480 11772 11486 11784
rect 12894 11772 12900 11784
rect 12952 11772 12958 11824
rect 13170 11772 13176 11824
rect 13228 11812 13234 11824
rect 13228 11784 14127 11812
rect 13228 11772 13234 11784
rect 12253 11747 12311 11753
rect 11164 11716 12204 11744
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11645 4859 11679
rect 5626 11676 5632 11688
rect 5587 11648 5632 11676
rect 4801 11639 4859 11645
rect 4341 11611 4399 11617
rect 4341 11577 4353 11611
rect 4387 11577 4399 11611
rect 4816 11608 4844 11639
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 6917 11679 6975 11685
rect 6917 11645 6929 11679
rect 6963 11645 6975 11679
rect 6917 11639 6975 11645
rect 5644 11608 5672 11636
rect 4816 11580 5672 11608
rect 6181 11611 6239 11617
rect 4341 11571 4399 11577
rect 6181 11577 6193 11611
rect 6227 11608 6239 11611
rect 6730 11608 6736 11620
rect 6227 11580 6736 11608
rect 6227 11577 6239 11580
rect 6181 11571 6239 11577
rect 6730 11568 6736 11580
rect 6788 11568 6794 11620
rect 3786 11540 3792 11552
rect 2424 11512 3792 11540
rect 2317 11503 2375 11509
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 5994 11540 6000 11552
rect 4764 11512 6000 11540
rect 4764 11500 4770 11512
rect 5994 11500 6000 11512
rect 6052 11500 6058 11552
rect 6932 11540 6960 11639
rect 7006 11636 7012 11688
rect 7064 11685 7070 11688
rect 7064 11679 7113 11685
rect 7064 11645 7067 11679
rect 7101 11645 7113 11679
rect 7064 11639 7113 11645
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11676 7987 11679
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 7975 11648 8677 11676
rect 7975 11645 7987 11648
rect 7929 11639 7987 11645
rect 7064 11636 7070 11639
rect 7285 11543 7343 11549
rect 7285 11540 7297 11543
rect 6932 11512 7297 11540
rect 7285 11509 7297 11512
rect 7331 11509 7343 11543
rect 7285 11503 7343 11509
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8303 11540 8331 11648
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11645 9275 11679
rect 9217 11639 9275 11645
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11645 12127 11679
rect 12176 11676 12204 11716
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12342 11744 12348 11756
rect 12299 11716 12348 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 12618 11704 12624 11756
rect 12676 11704 12682 11756
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 13354 11744 13360 11756
rect 13127 11716 13360 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 13354 11704 13360 11716
rect 13412 11744 13418 11756
rect 13630 11744 13636 11756
rect 13412 11716 13636 11744
rect 13412 11704 13418 11716
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 12636 11676 12664 11704
rect 12176 11648 12664 11676
rect 12805 11679 12863 11685
rect 12069 11639 12127 11645
rect 12805 11645 12817 11679
rect 12851 11645 12863 11679
rect 12805 11639 12863 11645
rect 12989 11679 13047 11685
rect 12989 11645 13001 11679
rect 13035 11645 13047 11679
rect 12989 11639 13047 11645
rect 8478 11568 8484 11620
rect 8536 11608 8542 11620
rect 9232 11608 9260 11639
rect 11422 11608 11428 11620
rect 8536 11580 9260 11608
rect 9692 11580 9996 11608
rect 8536 11568 8542 11580
rect 7892 11512 8331 11540
rect 7892 11500 7898 11512
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 9692 11540 9720 11580
rect 9858 11540 9864 11552
rect 8904 11512 9720 11540
rect 9819 11512 9864 11540
rect 8904 11500 8910 11512
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 9968 11540 9996 11580
rect 10980 11580 11428 11608
rect 10980 11540 11008 11580
rect 11422 11568 11428 11580
rect 11480 11568 11486 11620
rect 12084 11608 12112 11639
rect 12158 11608 12164 11620
rect 12084 11580 12164 11608
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 12250 11568 12256 11620
rect 12308 11608 12314 11620
rect 12820 11608 12848 11639
rect 12308 11580 12848 11608
rect 13004 11608 13032 11639
rect 13170 11636 13176 11688
rect 13228 11676 13234 11688
rect 14099 11685 14127 11784
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 15657 11815 15715 11821
rect 15657 11812 15669 11815
rect 14516 11784 15669 11812
rect 14516 11772 14522 11784
rect 15657 11781 15669 11784
rect 15703 11781 15715 11815
rect 15657 11775 15715 11781
rect 18322 11772 18328 11824
rect 18380 11812 18386 11824
rect 18782 11812 18788 11824
rect 18380 11784 18788 11812
rect 18380 11772 18386 11784
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11744 14795 11747
rect 15470 11744 15476 11756
rect 14783 11716 15476 11744
rect 14783 11713 14795 11716
rect 14737 11707 14795 11713
rect 15470 11704 15476 11716
rect 15528 11704 15534 11756
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 16390 11744 16396 11756
rect 15611 11716 16396 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 16632 11716 17141 11744
rect 16632 11704 16638 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 17494 11704 17500 11756
rect 17552 11744 17558 11756
rect 17678 11744 17684 11756
rect 17552 11716 17684 11744
rect 17552 11704 17558 11716
rect 17678 11704 17684 11716
rect 17736 11744 17742 11756
rect 18046 11744 18052 11756
rect 17736 11716 18052 11744
rect 17736 11704 17742 11716
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 18432 11753 18460 11784
rect 18782 11772 18788 11784
rect 18840 11812 18846 11824
rect 18840 11784 19012 11812
rect 18840 11772 18846 11784
rect 18984 11753 19012 11784
rect 19334 11772 19340 11824
rect 19392 11812 19398 11824
rect 21266 11812 21272 11824
rect 19392 11784 21272 11812
rect 19392 11772 19398 11784
rect 21266 11772 21272 11784
rect 21324 11772 21330 11824
rect 18417 11747 18475 11753
rect 18417 11713 18429 11747
rect 18463 11713 18475 11747
rect 18417 11707 18475 11713
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11713 18935 11747
rect 18877 11707 18935 11713
rect 18969 11747 19027 11753
rect 18969 11713 18981 11747
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 14001 11679 14059 11685
rect 14001 11676 14013 11679
rect 13228 11648 14013 11676
rect 13228 11636 13234 11648
rect 14001 11645 14013 11648
rect 14047 11645 14059 11679
rect 14001 11639 14059 11645
rect 14093 11679 14151 11685
rect 14093 11645 14105 11679
rect 14139 11645 14151 11679
rect 14093 11639 14151 11645
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 14332 11648 14473 11676
rect 14332 11636 14338 11648
rect 14461 11645 14473 11648
rect 14507 11645 14519 11679
rect 14642 11676 14648 11688
rect 14603 11648 14648 11676
rect 14461 11639 14519 11645
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 14918 11636 14924 11688
rect 14976 11676 14982 11688
rect 15194 11676 15200 11688
rect 14976 11648 15200 11676
rect 14976 11636 14982 11648
rect 15194 11636 15200 11648
rect 15252 11636 15258 11688
rect 15841 11679 15899 11685
rect 15841 11645 15853 11679
rect 15887 11676 15899 11679
rect 16206 11676 16212 11688
rect 15887 11648 16212 11676
rect 15887 11645 15899 11648
rect 15841 11639 15899 11645
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 16301 11679 16359 11685
rect 16301 11645 16313 11679
rect 16347 11676 16359 11679
rect 16758 11676 16764 11688
rect 16347 11648 16764 11676
rect 16347 11645 16359 11648
rect 16301 11639 16359 11645
rect 16758 11636 16764 11648
rect 16816 11636 16822 11688
rect 17221 11679 17279 11685
rect 17221 11645 17233 11679
rect 17267 11645 17279 11679
rect 17586 11676 17592 11688
rect 17547 11648 17592 11676
rect 17221 11639 17279 11645
rect 14366 11608 14372 11620
rect 13004 11580 14372 11608
rect 12308 11568 12314 11580
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 16114 11568 16120 11620
rect 16172 11608 16178 11620
rect 17236 11608 17264 11639
rect 17586 11636 17592 11648
rect 17644 11636 17650 11688
rect 17770 11676 17776 11688
rect 17731 11648 17776 11676
rect 17770 11636 17776 11648
rect 17828 11636 17834 11688
rect 16172 11580 17264 11608
rect 16172 11568 16178 11580
rect 17678 11568 17684 11620
rect 17736 11608 17742 11620
rect 18693 11611 18751 11617
rect 18693 11608 18705 11611
rect 17736 11580 18705 11608
rect 17736 11568 17742 11580
rect 18693 11577 18705 11580
rect 18739 11577 18751 11611
rect 18693 11571 18751 11577
rect 9968 11512 11008 11540
rect 11054 11500 11060 11552
rect 11112 11540 11118 11552
rect 11517 11543 11575 11549
rect 11517 11540 11529 11543
rect 11112 11512 11529 11540
rect 11112 11500 11118 11512
rect 11517 11509 11529 11512
rect 11563 11509 11575 11543
rect 11517 11503 11575 11509
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 11664 11512 11713 11540
rect 11664 11500 11670 11512
rect 11701 11509 11713 11512
rect 11747 11509 11759 11543
rect 11701 11503 11759 11509
rect 12621 11543 12679 11549
rect 12621 11509 12633 11543
rect 12667 11540 12679 11543
rect 12894 11540 12900 11552
rect 12667 11512 12900 11540
rect 12667 11509 12679 11512
rect 12621 11503 12679 11509
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 13541 11543 13599 11549
rect 13541 11540 13553 11543
rect 13320 11512 13553 11540
rect 13320 11500 13326 11512
rect 13541 11509 13553 11512
rect 13587 11509 13599 11543
rect 13541 11503 13599 11509
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 16390 11540 16396 11552
rect 15252 11512 15297 11540
rect 16351 11512 16396 11540
rect 15252 11500 15258 11512
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 17310 11540 17316 11552
rect 16908 11512 17316 11540
rect 16908 11500 16914 11512
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 18138 11540 18144 11552
rect 17460 11512 18144 11540
rect 17460 11500 17466 11512
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 18601 11543 18659 11549
rect 18601 11509 18613 11543
rect 18647 11540 18659 11543
rect 18892 11540 18920 11707
rect 19058 11704 19064 11756
rect 19116 11744 19122 11756
rect 19225 11747 19283 11753
rect 19225 11744 19237 11747
rect 19116 11716 19237 11744
rect 19116 11704 19122 11716
rect 19225 11713 19237 11716
rect 19271 11713 19283 11747
rect 19225 11707 19283 11713
rect 20254 11704 20260 11756
rect 20312 11744 20318 11756
rect 20625 11747 20683 11753
rect 20625 11744 20637 11747
rect 20312 11716 20637 11744
rect 20312 11704 20318 11716
rect 20625 11713 20637 11716
rect 20671 11713 20683 11747
rect 20625 11707 20683 11713
rect 20806 11636 20812 11688
rect 20864 11676 20870 11688
rect 21269 11679 21327 11685
rect 21269 11676 21281 11679
rect 20864 11648 21281 11676
rect 20864 11636 20870 11648
rect 21269 11645 21281 11648
rect 21315 11645 21327 11679
rect 21542 11676 21548 11688
rect 21503 11648 21548 11676
rect 21269 11639 21327 11645
rect 21542 11636 21548 11648
rect 21600 11636 21606 11688
rect 22848 11620 22876 11840
rect 22738 11608 22744 11620
rect 21284 11580 22744 11608
rect 18966 11540 18972 11552
rect 18647 11512 18972 11540
rect 18647 11509 18659 11512
rect 18601 11503 18659 11509
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 19150 11500 19156 11552
rect 19208 11540 19214 11552
rect 21284 11540 21312 11580
rect 22738 11568 22744 11580
rect 22796 11568 22802 11620
rect 22830 11568 22836 11620
rect 22888 11568 22894 11620
rect 19208 11512 21312 11540
rect 19208 11500 19214 11512
rect 21358 11500 21364 11552
rect 21416 11540 21422 11552
rect 22094 11540 22100 11552
rect 21416 11512 22100 11540
rect 21416 11500 21422 11512
rect 22094 11500 22100 11512
rect 22152 11500 22158 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1946 11296 1952 11348
rect 2004 11336 2010 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 2004 11308 3801 11336
rect 2004 11296 2010 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 3789 11299 3847 11305
rect 4430 11296 4436 11348
rect 4488 11296 4494 11348
rect 5258 11296 5264 11348
rect 5316 11336 5322 11348
rect 5316 11308 5580 11336
rect 5316 11296 5322 11308
rect 1670 11268 1676 11280
rect 1631 11240 1676 11268
rect 1670 11228 1676 11240
rect 1728 11228 1734 11280
rect 3602 11268 3608 11280
rect 3563 11240 3608 11268
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 3326 11160 3332 11212
rect 3384 11200 3390 11212
rect 4448 11209 4476 11296
rect 4433 11203 4491 11209
rect 3384 11172 4384 11200
rect 3384 11160 3390 11172
rect 1486 11132 1492 11144
rect 1447 11104 1492 11132
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 2498 11141 2504 11144
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11101 2283 11135
rect 2492 11132 2504 11141
rect 2459 11104 2504 11132
rect 2225 11095 2283 11101
rect 2492 11095 2504 11104
rect 1854 11064 1860 11076
rect 1815 11036 1860 11064
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 2038 11064 2044 11076
rect 1999 11036 2044 11064
rect 2038 11024 2044 11036
rect 2096 11024 2102 11076
rect 2240 11064 2268 11095
rect 2498 11092 2504 11095
rect 2556 11092 2562 11144
rect 3970 11132 3976 11144
rect 3931 11104 3976 11132
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 4356 11132 4384 11172
rect 4433 11169 4445 11203
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 4522 11160 4528 11212
rect 4580 11200 4586 11212
rect 5552 11200 5580 11308
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 5868 11308 6745 11336
rect 5868 11296 5874 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 6733 11299 6791 11305
rect 6840 11308 6960 11336
rect 5626 11228 5632 11280
rect 5684 11268 5690 11280
rect 5905 11271 5963 11277
rect 5905 11268 5917 11271
rect 5684 11240 5917 11268
rect 5684 11228 5690 11240
rect 5905 11237 5917 11240
rect 5951 11237 5963 11271
rect 6641 11271 6699 11277
rect 6641 11268 6653 11271
rect 5905 11231 5963 11237
rect 6012 11240 6653 11268
rect 6012 11200 6040 11240
rect 6641 11237 6653 11240
rect 6687 11268 6699 11271
rect 6840 11268 6868 11308
rect 6687 11240 6868 11268
rect 6932 11268 6960 11308
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 7561 11339 7619 11345
rect 7561 11336 7573 11339
rect 7524 11308 7573 11336
rect 7524 11296 7530 11308
rect 7561 11305 7573 11308
rect 7607 11305 7619 11339
rect 8754 11336 8760 11348
rect 8715 11308 8760 11336
rect 7561 11299 7619 11305
rect 8754 11296 8760 11308
rect 8812 11296 8818 11348
rect 8864 11308 10180 11336
rect 7006 11268 7012 11280
rect 6932 11240 7012 11268
rect 6687 11237 6699 11240
rect 6641 11231 6699 11237
rect 7006 11228 7012 11240
rect 7064 11268 7070 11280
rect 8864 11268 8892 11308
rect 7064 11240 8892 11268
rect 7064 11228 7070 11240
rect 4580 11172 4625 11200
rect 5552 11172 6040 11200
rect 4580 11160 4586 11172
rect 6086 11160 6092 11212
rect 6144 11200 6150 11212
rect 6362 11200 6368 11212
rect 6144 11172 6189 11200
rect 6323 11172 6368 11200
rect 6144 11160 6150 11172
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 7098 11200 7104 11212
rect 7024 11172 7104 11200
rect 6914 11132 6920 11144
rect 4356 11104 6920 11132
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7024 11132 7052 11172
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 7377 11203 7435 11209
rect 7377 11200 7389 11203
rect 7361 11169 7389 11200
rect 7423 11169 7435 11203
rect 7361 11163 7435 11169
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11200 8263 11203
rect 9030 11200 9036 11212
rect 8251 11172 9036 11200
rect 8251 11169 8263 11172
rect 8205 11163 8263 11169
rect 7361 11132 7389 11163
rect 9030 11160 9036 11172
rect 9088 11160 9094 11212
rect 9122 11160 9128 11212
rect 9180 11200 9186 11212
rect 10152 11200 10180 11308
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 11241 11339 11299 11345
rect 11241 11336 11253 11339
rect 10744 11308 11253 11336
rect 10744 11296 10750 11308
rect 11241 11305 11253 11308
rect 11287 11336 11299 11339
rect 11422 11336 11428 11348
rect 11287 11308 11428 11336
rect 11287 11305 11299 11308
rect 11241 11299 11299 11305
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 11517 11339 11575 11345
rect 11517 11305 11529 11339
rect 11563 11336 11575 11339
rect 11698 11336 11704 11348
rect 11563 11308 11704 11336
rect 11563 11305 11575 11308
rect 11517 11299 11575 11305
rect 11698 11296 11704 11308
rect 11756 11336 11762 11348
rect 12342 11336 12348 11348
rect 11756 11308 12204 11336
rect 12303 11308 12348 11336
rect 11756 11296 11762 11308
rect 10870 11268 10876 11280
rect 10831 11240 10876 11268
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 12176 11268 12204 11308
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 13170 11336 13176 11348
rect 13131 11308 13176 11336
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 13354 11336 13360 11348
rect 13315 11308 13360 11336
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13814 11336 13820 11348
rect 13775 11308 13820 11336
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 14553 11339 14611 11345
rect 14553 11336 14565 11339
rect 14516 11308 14565 11336
rect 14516 11296 14522 11308
rect 14553 11305 14565 11308
rect 14599 11305 14611 11339
rect 14553 11299 14611 11305
rect 14642 11296 14648 11348
rect 14700 11336 14706 11348
rect 14737 11339 14795 11345
rect 14737 11336 14749 11339
rect 14700 11308 14749 11336
rect 14700 11296 14706 11308
rect 14737 11305 14749 11308
rect 14783 11305 14795 11339
rect 14737 11299 14795 11305
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 15565 11339 15623 11345
rect 15565 11336 15577 11339
rect 15528 11308 15577 11336
rect 15528 11296 15534 11308
rect 15565 11305 15577 11308
rect 15611 11305 15623 11339
rect 15565 11299 15623 11305
rect 15930 11296 15936 11348
rect 15988 11336 15994 11348
rect 16393 11339 16451 11345
rect 16393 11336 16405 11339
rect 15988 11308 16405 11336
rect 15988 11296 15994 11308
rect 16393 11305 16405 11308
rect 16439 11305 16451 11339
rect 16393 11299 16451 11305
rect 17126 11296 17132 11348
rect 17184 11336 17190 11348
rect 17221 11339 17279 11345
rect 17221 11336 17233 11339
rect 17184 11308 17233 11336
rect 17184 11296 17190 11308
rect 17221 11305 17233 11308
rect 17267 11305 17279 11339
rect 17221 11299 17279 11305
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 17368 11308 17417 11336
rect 17368 11296 17374 11308
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 17862 11336 17868 11348
rect 17405 11299 17463 11305
rect 17696 11308 17868 11336
rect 14369 11271 14427 11277
rect 14369 11268 14381 11271
rect 10980 11240 11928 11268
rect 12176 11240 14381 11268
rect 10980 11200 11008 11240
rect 11790 11200 11796 11212
rect 9180 11172 9225 11200
rect 10152 11172 11008 11200
rect 11751 11172 11796 11200
rect 9180 11160 9186 11172
rect 11790 11160 11796 11172
rect 11848 11160 11854 11212
rect 11900 11200 11928 11240
rect 11900 11172 12204 11200
rect 7024 11104 7389 11132
rect 7929 11135 7987 11141
rect 2958 11064 2964 11076
rect 2240 11036 2964 11064
rect 2958 11024 2964 11036
rect 3016 11064 3022 11076
rect 3418 11064 3424 11076
rect 3016 11036 3424 11064
rect 3016 11024 3022 11036
rect 3418 11024 3424 11036
rect 3476 11024 3482 11076
rect 4157 11067 4215 11073
rect 4157 11033 4169 11067
rect 4203 11064 4215 11067
rect 4522 11064 4528 11076
rect 4203 11036 4528 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 4522 11024 4528 11036
rect 4580 11024 4586 11076
rect 4798 11073 4804 11076
rect 4792 11064 4804 11073
rect 4759 11036 4804 11064
rect 4792 11027 4804 11036
rect 4798 11024 4804 11027
rect 4856 11024 4862 11076
rect 5626 11024 5632 11076
rect 5684 11064 5690 11076
rect 6362 11064 6368 11076
rect 5684 11036 6368 11064
rect 5684 11024 5690 11036
rect 6362 11024 6368 11036
rect 6420 11024 6426 11076
rect 6546 11024 6552 11076
rect 6604 11064 6610 11076
rect 7024 11064 7052 11104
rect 7929 11101 7941 11135
rect 7975 11132 7987 11135
rect 8294 11132 8300 11144
rect 7975 11104 8300 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11132 8447 11135
rect 8570 11132 8576 11144
rect 8435 11104 8576 11132
rect 8435 11101 8447 11104
rect 8389 11095 8447 11101
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 8938 11132 8944 11144
rect 8851 11104 8944 11132
rect 8938 11092 8944 11104
rect 8996 11132 9002 11144
rect 8996 11104 10180 11132
rect 8996 11092 9002 11104
rect 7558 11064 7564 11076
rect 6604 11036 7052 11064
rect 7300 11036 7564 11064
rect 6604 11024 6610 11036
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 6178 10996 6184 11008
rect 3200 10968 6184 10996
rect 3200 10956 3206 10968
rect 6178 10956 6184 10968
rect 6236 10956 6242 11008
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 7101 10999 7159 11005
rect 7101 10996 7113 10999
rect 7064 10968 7113 10996
rect 7064 10956 7070 10968
rect 7101 10965 7113 10968
rect 7147 10965 7159 10999
rect 7101 10959 7159 10965
rect 7193 10999 7251 11005
rect 7193 10965 7205 10999
rect 7239 10996 7251 10999
rect 7300 10996 7328 11036
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 8478 11024 8484 11076
rect 8536 11064 8542 11076
rect 9370 11067 9428 11073
rect 9370 11064 9382 11067
rect 8536 11036 9382 11064
rect 8536 11024 8542 11036
rect 9370 11033 9382 11036
rect 9416 11033 9428 11067
rect 10152 11064 10180 11104
rect 11698 11092 11704 11144
rect 11756 11132 11762 11144
rect 11977 11135 12035 11141
rect 11756 11104 11937 11132
rect 11756 11092 11762 11104
rect 11909 11064 11937 11104
rect 11977 11101 11989 11135
rect 12023 11132 12035 11135
rect 12066 11132 12072 11144
rect 12023 11104 12072 11132
rect 12023 11101 12035 11104
rect 11977 11095 12035 11101
rect 12066 11092 12072 11104
rect 12124 11092 12130 11144
rect 12176 11132 12204 11172
rect 12342 11160 12348 11212
rect 12400 11200 12406 11212
rect 12529 11203 12587 11209
rect 12529 11200 12541 11203
rect 12400 11172 12541 11200
rect 12400 11160 12406 11172
rect 12529 11169 12541 11172
rect 12575 11169 12587 11203
rect 12774 11200 12802 11240
rect 14369 11237 14381 11240
rect 14415 11268 14427 11271
rect 17696 11268 17724 11308
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 18046 11296 18052 11348
rect 18104 11336 18110 11348
rect 18104 11308 18736 11336
rect 18104 11296 18110 11308
rect 14415 11240 17080 11268
rect 14415 11237 14427 11240
rect 14369 11231 14427 11237
rect 12774 11172 12848 11200
rect 12529 11163 12587 11169
rect 12710 11132 12716 11144
rect 12176 11104 12716 11132
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12820 11141 12848 11172
rect 14458 11160 14464 11212
rect 14516 11200 14522 11212
rect 15010 11200 15016 11212
rect 14516 11172 15016 11200
rect 14516 11160 14522 11172
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 15194 11200 15200 11212
rect 15155 11172 15200 11200
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 15286 11160 15292 11212
rect 15344 11200 15350 11212
rect 16114 11200 16120 11212
rect 15344 11172 16120 11200
rect 15344 11160 15350 11172
rect 16114 11160 16120 11172
rect 16172 11200 16178 11212
rect 16945 11203 17003 11209
rect 16945 11200 16957 11203
rect 16172 11172 16957 11200
rect 16172 11160 16178 11172
rect 16945 11169 16957 11172
rect 16991 11169 17003 11203
rect 16945 11163 17003 11169
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11101 12863 11135
rect 16022 11132 16028 11144
rect 12805 11095 12863 11101
rect 14200 11104 16028 11132
rect 13630 11064 13636 11076
rect 10152 11036 11744 11064
rect 11909 11036 12296 11064
rect 13591 11036 13636 11064
rect 9370 11027 9428 11033
rect 11716 11008 11744 11036
rect 7239 10968 7328 10996
rect 7239 10965 7251 10968
rect 7193 10959 7251 10965
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 8202 10996 8208 11008
rect 7708 10968 8208 10996
rect 7708 10956 7714 10968
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 10502 10996 10508 11008
rect 10463 10968 10508 10996
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 11146 10996 11152 11008
rect 10652 10968 10697 10996
rect 11107 10968 11152 10996
rect 10652 10956 10658 10968
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 11698 10956 11704 11008
rect 11756 10956 11762 11008
rect 11885 10999 11943 11005
rect 11885 10965 11897 10999
rect 11931 10996 11943 10999
rect 11974 10996 11980 11008
rect 11931 10968 11980 10996
rect 11931 10965 11943 10968
rect 11885 10959 11943 10965
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 12268 10996 12296 11036
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 12713 10999 12771 11005
rect 12713 10996 12725 10999
rect 12268 10968 12725 10996
rect 12713 10965 12725 10968
rect 12759 10996 12771 10999
rect 13170 10996 13176 11008
rect 12759 10968 13176 10996
rect 12759 10965 12771 10968
rect 12713 10959 12771 10965
rect 13170 10956 13176 10968
rect 13228 10996 13234 11008
rect 14200 10996 14228 11104
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 16758 11132 16764 11144
rect 16719 11104 16764 11132
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 16908 11104 16953 11132
rect 16908 11092 16914 11104
rect 14277 11067 14335 11073
rect 14277 11033 14289 11067
rect 14323 11064 14335 11067
rect 15010 11064 15016 11076
rect 14323 11036 15016 11064
rect 14323 11033 14335 11036
rect 14277 11027 14335 11033
rect 15010 11024 15016 11036
rect 15068 11024 15074 11076
rect 15105 11067 15163 11073
rect 15105 11033 15117 11067
rect 15151 11064 15163 11067
rect 16942 11064 16948 11076
rect 15151 11036 16948 11064
rect 15151 11033 15163 11036
rect 15105 11027 15163 11033
rect 16942 11024 16948 11036
rect 17000 11024 17006 11076
rect 17052 11064 17080 11240
rect 17144 11240 17724 11268
rect 17144 11212 17172 11240
rect 17126 11160 17132 11212
rect 17184 11160 17190 11212
rect 17678 11200 17684 11212
rect 17639 11172 17684 11200
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 18708 11200 18736 11308
rect 18782 11296 18788 11348
rect 18840 11336 18846 11348
rect 18840 11308 20668 11336
rect 18840 11296 18846 11308
rect 19058 11268 19064 11280
rect 18971 11240 19064 11268
rect 19058 11228 19064 11240
rect 19116 11268 19122 11280
rect 19242 11268 19248 11280
rect 19116 11240 19248 11268
rect 19116 11228 19122 11240
rect 19242 11228 19248 11240
rect 19300 11228 19306 11280
rect 20640 11209 20668 11308
rect 20625 11203 20683 11209
rect 18708 11172 19380 11200
rect 17310 11092 17316 11144
rect 17368 11132 17374 11144
rect 17368 11104 19288 11132
rect 17368 11092 17374 11104
rect 17586 11064 17592 11076
rect 17052 11036 17592 11064
rect 17586 11024 17592 11036
rect 17644 11024 17650 11076
rect 17948 11067 18006 11073
rect 17948 11033 17960 11067
rect 17994 11064 18006 11067
rect 18690 11064 18696 11076
rect 17994 11036 18696 11064
rect 17994 11033 18006 11036
rect 17948 11027 18006 11033
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 15930 10996 15936 11008
rect 13228 10968 14228 10996
rect 15891 10968 15936 10996
rect 13228 10956 13234 10968
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 16022 10956 16028 11008
rect 16080 10996 16086 11008
rect 16080 10968 16125 10996
rect 16080 10956 16086 10968
rect 16206 10956 16212 11008
rect 16264 10996 16270 11008
rect 17310 10996 17316 11008
rect 16264 10968 17316 10996
rect 16264 10956 16270 10968
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 18230 10956 18236 11008
rect 18288 10996 18294 11008
rect 18506 10996 18512 11008
rect 18288 10968 18512 10996
rect 18288 10956 18294 10968
rect 18506 10956 18512 10968
rect 18564 10956 18570 11008
rect 19260 11005 19288 11104
rect 19352 11064 19380 11172
rect 20625 11169 20637 11203
rect 20671 11169 20683 11203
rect 21266 11200 21272 11212
rect 21227 11172 21272 11200
rect 20625 11163 20683 11169
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 20346 11092 20352 11144
rect 20404 11141 20410 11144
rect 20404 11132 20416 11141
rect 20404 11104 20449 11132
rect 20404 11095 20416 11104
rect 20404 11092 20410 11095
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 21177 11135 21235 11141
rect 21177 11132 21189 11135
rect 20772 11104 21189 11132
rect 20772 11092 20778 11104
rect 21177 11101 21189 11104
rect 21223 11101 21235 11135
rect 21177 11095 21235 11101
rect 21085 11067 21143 11073
rect 21085 11064 21097 11067
rect 19352 11036 21097 11064
rect 21085 11033 21097 11036
rect 21131 11033 21143 11067
rect 21085 11027 21143 11033
rect 19245 10999 19303 11005
rect 19245 10965 19257 10999
rect 19291 10965 19303 10999
rect 19245 10959 19303 10965
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 20346 10996 20352 11008
rect 19852 10968 20352 10996
rect 19852 10956 19858 10968
rect 20346 10956 20352 10968
rect 20404 10956 20410 11008
rect 20717 10999 20775 11005
rect 20717 10965 20729 10999
rect 20763 10996 20775 10999
rect 20806 10996 20812 11008
rect 20763 10968 20812 10996
rect 20763 10965 20775 10968
rect 20717 10959 20775 10965
rect 20806 10956 20812 10968
rect 20864 10956 20870 11008
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 2498 10792 2504 10804
rect 1627 10764 2504 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3421 10795 3479 10801
rect 3421 10792 3433 10795
rect 2832 10764 3433 10792
rect 2832 10752 2838 10764
rect 3421 10761 3433 10764
rect 3467 10761 3479 10795
rect 3421 10755 3479 10761
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 5166 10792 5172 10804
rect 4856 10764 5172 10792
rect 4856 10752 4862 10764
rect 5166 10752 5172 10764
rect 5224 10792 5230 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5224 10764 5641 10792
rect 5224 10752 5230 10764
rect 5629 10761 5641 10764
rect 5675 10792 5687 10795
rect 6546 10792 6552 10804
rect 5675 10764 6552 10792
rect 5675 10761 5687 10764
rect 5629 10755 5687 10761
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 6733 10795 6791 10801
rect 6733 10761 6745 10795
rect 6779 10792 6791 10795
rect 6822 10792 6828 10804
rect 6779 10764 6828 10792
rect 6779 10761 6791 10764
rect 6733 10755 6791 10761
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 7009 10795 7067 10801
rect 7009 10761 7021 10795
rect 7055 10792 7067 10795
rect 7558 10792 7564 10804
rect 7055 10764 7564 10792
rect 7055 10761 7067 10764
rect 7009 10755 7067 10761
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 7742 10752 7748 10804
rect 7800 10792 7806 10804
rect 7926 10792 7932 10804
rect 7800 10764 7932 10792
rect 7800 10752 7806 10764
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 8294 10792 8300 10804
rect 8255 10764 8300 10792
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 8386 10752 8392 10804
rect 8444 10792 8450 10804
rect 8662 10792 8668 10804
rect 8444 10764 8668 10792
rect 8444 10752 8450 10764
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 9766 10792 9772 10804
rect 9727 10764 9772 10792
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 10137 10795 10195 10801
rect 10137 10761 10149 10795
rect 10183 10792 10195 10795
rect 10594 10792 10600 10804
rect 10183 10764 10600 10792
rect 10183 10761 10195 10764
rect 10137 10755 10195 10761
rect 10594 10752 10600 10764
rect 10652 10752 10658 10804
rect 11793 10795 11851 10801
rect 11793 10761 11805 10795
rect 11839 10792 11851 10795
rect 11882 10792 11888 10804
rect 11839 10764 11888 10792
rect 11839 10761 11851 10764
rect 11793 10755 11851 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12066 10752 12072 10804
rect 12124 10792 12130 10804
rect 12342 10792 12348 10804
rect 12124 10764 12348 10792
rect 12124 10752 12130 10764
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 13078 10752 13084 10804
rect 13136 10792 13142 10804
rect 13538 10792 13544 10804
rect 13136 10764 13544 10792
rect 13136 10752 13142 10764
rect 13538 10752 13544 10764
rect 13596 10792 13602 10804
rect 14185 10795 14243 10801
rect 14185 10792 14197 10795
rect 13596 10764 14197 10792
rect 13596 10752 13602 10764
rect 14185 10761 14197 10764
rect 14231 10761 14243 10795
rect 14366 10792 14372 10804
rect 14327 10764 14372 10792
rect 14185 10755 14243 10761
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 15930 10792 15936 10804
rect 14467 10764 15936 10792
rect 1762 10684 1768 10736
rect 1820 10724 1826 10736
rect 1820 10696 3280 10724
rect 1820 10684 1826 10696
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 3252 10665 3280 10696
rect 3602 10684 3608 10736
rect 3660 10724 3666 10736
rect 4516 10727 4574 10733
rect 4516 10724 4528 10727
rect 3660 10696 4528 10724
rect 3660 10684 3666 10696
rect 4516 10693 4528 10696
rect 4562 10724 4574 10727
rect 6917 10727 6975 10733
rect 4562 10696 6868 10724
rect 4562 10693 4574 10696
rect 4516 10687 4574 10693
rect 2694 10659 2752 10665
rect 2694 10656 2706 10659
rect 1912 10628 2706 10656
rect 1912 10616 1918 10628
rect 2694 10625 2706 10628
rect 2740 10656 2752 10659
rect 3237 10659 3295 10665
rect 2740 10628 3188 10656
rect 2740 10625 2752 10628
rect 2694 10619 2752 10625
rect 2958 10588 2964 10600
rect 2919 10560 2964 10588
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 3160 10520 3188 10628
rect 3237 10625 3249 10659
rect 3283 10625 3295 10659
rect 3237 10619 3295 10625
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10656 3847 10659
rect 4338 10656 4344 10668
rect 3835 10628 4344 10656
rect 3835 10625 3847 10628
rect 3789 10619 3847 10625
rect 4338 10616 4344 10628
rect 4396 10616 4402 10668
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5408 10628 5733 10656
rect 5408 10616 5414 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10656 6055 10659
rect 6730 10656 6736 10668
rect 6043 10628 6736 10656
rect 6043 10625 6055 10628
rect 5997 10619 6055 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 3878 10588 3884 10600
rect 3839 10560 3884 10588
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10557 4031 10591
rect 4246 10588 4252 10600
rect 4207 10560 4252 10588
rect 3973 10551 4031 10557
rect 3988 10520 4016 10551
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 6365 10591 6423 10597
rect 6365 10588 6377 10591
rect 5960 10560 6377 10588
rect 5960 10548 5966 10560
rect 6365 10557 6377 10560
rect 6411 10557 6423 10591
rect 6840 10588 6868 10696
rect 6917 10693 6929 10727
rect 6963 10724 6975 10727
rect 7374 10724 7380 10736
rect 6963 10696 7380 10724
rect 6963 10693 6975 10696
rect 6917 10687 6975 10693
rect 7374 10684 7380 10696
rect 7432 10684 7438 10736
rect 7469 10727 7527 10733
rect 7469 10693 7481 10727
rect 7515 10724 7527 10727
rect 8938 10724 8944 10736
rect 7515 10696 7972 10724
rect 7515 10693 7527 10696
rect 7469 10687 7527 10693
rect 7006 10616 7012 10668
rect 7064 10656 7070 10668
rect 7282 10656 7288 10668
rect 7064 10628 7288 10656
rect 7064 10616 7070 10628
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7834 10660 7840 10668
rect 7576 10656 7687 10660
rect 7760 10656 7840 10660
rect 7576 10632 7840 10656
rect 7576 10597 7604 10632
rect 7659 10628 7788 10632
rect 7834 10616 7840 10632
rect 7892 10616 7898 10668
rect 7944 10665 7972 10696
rect 8128 10696 8944 10724
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 8018 10656 8024 10668
rect 7975 10628 8024 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 6840 10560 7573 10588
rect 6365 10551 6423 10557
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 8128 10588 8156 10696
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 9030 10684 9036 10736
rect 9088 10724 9094 10736
rect 9306 10724 9312 10736
rect 9088 10696 9312 10724
rect 9088 10684 9094 10696
rect 9306 10684 9312 10696
rect 9364 10724 9370 10736
rect 9410 10727 9468 10733
rect 9410 10724 9422 10727
rect 9364 10696 9422 10724
rect 9364 10684 9370 10696
rect 9410 10693 9422 10696
rect 9456 10724 9468 10727
rect 9456 10696 10456 10724
rect 9456 10693 9468 10696
rect 9410 10687 9468 10693
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10656 8263 10659
rect 9582 10656 9588 10668
rect 8251 10628 9588 10656
rect 8251 10625 8263 10628
rect 8205 10619 8263 10625
rect 7561 10551 7619 10557
rect 7760 10560 8156 10588
rect 6178 10520 6184 10532
rect 3160 10492 4016 10520
rect 5175 10492 6184 10520
rect 1486 10452 1492 10464
rect 1447 10424 1492 10452
rect 1486 10412 1492 10424
rect 1544 10412 1550 10464
rect 2222 10412 2228 10464
rect 2280 10452 2286 10464
rect 3053 10455 3111 10461
rect 3053 10452 3065 10455
rect 2280 10424 3065 10452
rect 2280 10412 2286 10424
rect 3053 10421 3065 10424
rect 3099 10421 3111 10455
rect 3053 10415 3111 10421
rect 3418 10412 3424 10464
rect 3476 10452 3482 10464
rect 5175 10452 5203 10492
rect 6178 10480 6184 10492
rect 6236 10480 6242 10532
rect 6454 10480 6460 10532
rect 6512 10520 6518 10532
rect 7650 10520 7656 10532
rect 6512 10492 7656 10520
rect 6512 10480 6518 10492
rect 7650 10480 7656 10492
rect 7708 10480 7714 10532
rect 3476 10424 5203 10452
rect 3476 10412 3482 10424
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6089 10455 6147 10461
rect 6089 10452 6101 10455
rect 6052 10424 6101 10452
rect 6052 10412 6058 10424
rect 6089 10421 6101 10424
rect 6135 10421 6147 10455
rect 6089 10415 6147 10421
rect 6362 10412 6368 10464
rect 6420 10452 6426 10464
rect 6822 10452 6828 10464
rect 6420 10424 6828 10452
rect 6420 10412 6426 10424
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7760 10452 7788 10560
rect 8018 10520 8024 10532
rect 7979 10492 8024 10520
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 7156 10424 7788 10452
rect 7156 10412 7162 10424
rect 7926 10412 7932 10464
rect 7984 10452 7990 10464
rect 8220 10452 8248 10619
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 8352 10560 8524 10588
rect 8352 10548 8358 10560
rect 7984 10424 8248 10452
rect 8496 10452 8524 10560
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 10229 10591 10287 10597
rect 9732 10560 9777 10588
rect 9732 10548 9738 10560
rect 10229 10557 10241 10591
rect 10275 10588 10287 10591
rect 10318 10588 10324 10600
rect 10275 10560 10324 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 10244 10520 10272 10551
rect 10318 10548 10324 10560
rect 10376 10548 10382 10600
rect 10428 10597 10456 10696
rect 11698 10684 11704 10736
rect 11756 10724 11762 10736
rect 11974 10724 11980 10736
rect 11756 10696 11980 10724
rect 11756 10684 11762 10696
rect 11974 10684 11980 10696
rect 12032 10684 12038 10736
rect 12158 10684 12164 10736
rect 12216 10724 12222 10736
rect 12590 10727 12648 10733
rect 12590 10724 12602 10727
rect 12216 10696 12602 10724
rect 12216 10684 12222 10696
rect 12590 10693 12602 10696
rect 12636 10693 12648 10727
rect 12590 10687 12648 10693
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 14467 10724 14495 10764
rect 15930 10752 15936 10764
rect 15988 10752 15994 10804
rect 16114 10792 16120 10804
rect 16075 10764 16120 10792
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 16669 10795 16727 10801
rect 16669 10761 16681 10795
rect 16715 10792 16727 10795
rect 16942 10792 16948 10804
rect 16715 10764 16948 10792
rect 16715 10761 16727 10764
rect 16669 10755 16727 10761
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 17586 10752 17592 10804
rect 17644 10792 17650 10804
rect 18046 10792 18052 10804
rect 17644 10764 18052 10792
rect 17644 10752 17650 10764
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 18414 10752 18420 10804
rect 18472 10792 18478 10804
rect 18509 10795 18567 10801
rect 18509 10792 18521 10795
rect 18472 10764 18521 10792
rect 18472 10752 18478 10764
rect 18509 10761 18521 10764
rect 18555 10761 18567 10795
rect 18509 10755 18567 10761
rect 19886 10752 19892 10804
rect 19944 10792 19950 10804
rect 20165 10795 20223 10801
rect 20165 10792 20177 10795
rect 19944 10764 20177 10792
rect 19944 10752 19950 10764
rect 20165 10761 20177 10764
rect 20211 10761 20223 10795
rect 20165 10755 20223 10761
rect 20254 10752 20260 10804
rect 20312 10792 20318 10804
rect 20312 10764 20357 10792
rect 20312 10752 20318 10764
rect 12768 10696 14495 10724
rect 15004 10727 15062 10733
rect 12768 10684 12774 10696
rect 15004 10693 15016 10727
rect 15050 10724 15062 10727
rect 15194 10724 15200 10736
rect 15050 10696 15200 10724
rect 15050 10693 15062 10696
rect 15004 10687 15062 10693
rect 15194 10684 15200 10696
rect 15252 10724 15258 10736
rect 16206 10724 16212 10736
rect 15252 10696 16212 10724
rect 15252 10684 15258 10696
rect 16206 10684 16212 10696
rect 16264 10684 16270 10736
rect 17862 10724 17868 10736
rect 17052 10696 17868 10724
rect 11146 10616 11152 10668
rect 11204 10656 11210 10668
rect 11333 10659 11391 10665
rect 11333 10656 11345 10659
rect 11204 10628 11345 10656
rect 11204 10616 11210 10628
rect 11333 10625 11345 10628
rect 11379 10656 11391 10659
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 11379 10628 11897 10656
rect 11379 10625 11391 10628
rect 11333 10619 11391 10625
rect 11885 10625 11897 10628
rect 11931 10656 11943 10659
rect 12250 10656 12256 10668
rect 11931 10628 12256 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 12345 10659 12403 10665
rect 12345 10625 12357 10659
rect 12391 10656 12403 10659
rect 12434 10656 12440 10668
rect 12391 10628 12440 10656
rect 12391 10625 12403 10628
rect 12345 10619 12403 10625
rect 12434 10616 12440 10628
rect 12492 10656 12498 10668
rect 14274 10656 14280 10668
rect 12492 10628 14280 10656
rect 12492 10616 12498 10628
rect 14274 10616 14280 10628
rect 14332 10656 14338 10668
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 14332 10628 14749 10656
rect 14332 10616 14338 10628
rect 14737 10625 14749 10628
rect 14783 10656 14795 10659
rect 15746 10656 15752 10668
rect 14783 10628 15752 10656
rect 14783 10625 14795 10628
rect 14737 10619 14795 10625
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 16942 10616 16948 10668
rect 17000 10656 17006 10668
rect 17052 10665 17080 10696
rect 17862 10684 17868 10696
rect 17920 10684 17926 10736
rect 17954 10684 17960 10736
rect 18012 10724 18018 10736
rect 20625 10727 20683 10733
rect 18012 10696 19196 10724
rect 18012 10684 18018 10696
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 17000 10628 17049 10656
rect 17000 10616 17006 10628
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17497 10659 17555 10665
rect 17497 10656 17509 10659
rect 17037 10619 17095 10625
rect 17144 10628 17509 10656
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10557 10471 10591
rect 10413 10551 10471 10557
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 11609 10591 11667 10597
rect 11609 10588 11621 10591
rect 11296 10560 11621 10588
rect 11296 10548 11302 10560
rect 11609 10557 11621 10560
rect 11655 10588 11667 10591
rect 12066 10588 12072 10600
rect 11655 10560 12072 10588
rect 11655 10557 11667 10560
rect 11609 10551 11667 10557
rect 12066 10548 12072 10560
rect 12124 10548 12130 10600
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10588 13967 10591
rect 14642 10588 14648 10600
rect 13955 10560 14648 10588
rect 13955 10557 13967 10560
rect 13909 10551 13967 10557
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 15930 10548 15936 10600
rect 15988 10588 15994 10600
rect 16209 10591 16267 10597
rect 16209 10588 16221 10591
rect 15988 10560 16221 10588
rect 15988 10548 15994 10560
rect 16209 10557 16221 10560
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 16850 10548 16856 10600
rect 16908 10588 16914 10600
rect 17144 10597 17172 10628
rect 17497 10625 17509 10628
rect 17543 10625 17555 10659
rect 17497 10619 17555 10625
rect 17129 10591 17187 10597
rect 17129 10588 17141 10591
rect 16908 10560 17141 10588
rect 16908 10548 16914 10560
rect 17129 10557 17141 10560
rect 17175 10557 17187 10591
rect 17310 10588 17316 10600
rect 17271 10560 17316 10588
rect 17129 10551 17187 10557
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 17972 10597 18000 10684
rect 18141 10659 18199 10665
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 18598 10656 18604 10668
rect 18187 10628 18604 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 18966 10656 18972 10668
rect 18708 10628 18972 10656
rect 17957 10591 18015 10597
rect 17957 10557 17969 10591
rect 18003 10557 18015 10591
rect 17957 10551 18015 10557
rect 18322 10548 18328 10600
rect 18380 10588 18386 10600
rect 18708 10588 18736 10628
rect 18966 10616 18972 10628
rect 19024 10616 19030 10668
rect 18380 10560 18736 10588
rect 18380 10548 18386 10560
rect 18782 10548 18788 10600
rect 18840 10588 18846 10600
rect 19168 10597 19196 10696
rect 20625 10693 20637 10727
rect 20671 10724 20683 10727
rect 20714 10724 20720 10736
rect 20671 10696 20720 10724
rect 20671 10693 20683 10696
rect 20625 10687 20683 10693
rect 20714 10684 20720 10696
rect 20772 10684 20778 10736
rect 21174 10684 21180 10736
rect 21232 10724 21238 10736
rect 21269 10727 21327 10733
rect 21269 10724 21281 10727
rect 21232 10696 21281 10724
rect 21232 10684 21238 10696
rect 21269 10693 21281 10696
rect 21315 10693 21327 10727
rect 21269 10687 21327 10693
rect 19794 10656 19800 10668
rect 19755 10628 19800 10656
rect 19794 10616 19800 10628
rect 19852 10616 19858 10668
rect 21082 10656 21088 10668
rect 21043 10628 21088 10656
rect 21082 10616 21088 10628
rect 21140 10616 21146 10668
rect 21450 10656 21456 10668
rect 21411 10628 21456 10656
rect 21450 10616 21456 10628
rect 21508 10616 21514 10668
rect 19061 10591 19119 10597
rect 19061 10588 19073 10591
rect 18840 10560 19073 10588
rect 18840 10548 18846 10560
rect 19061 10557 19073 10560
rect 19107 10557 19119 10591
rect 19061 10551 19119 10557
rect 19153 10591 19211 10597
rect 19153 10557 19165 10591
rect 19199 10557 19211 10591
rect 19153 10551 19211 10557
rect 19242 10548 19248 10600
rect 19300 10588 19306 10600
rect 19613 10591 19671 10597
rect 19613 10588 19625 10591
rect 19300 10560 19625 10588
rect 19300 10548 19306 10560
rect 19613 10557 19625 10560
rect 19659 10557 19671 10591
rect 19613 10551 19671 10557
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10588 19763 10591
rect 20162 10588 20168 10600
rect 19751 10560 20168 10588
rect 19751 10557 19763 10560
rect 19705 10551 19763 10557
rect 10781 10523 10839 10529
rect 10781 10520 10793 10523
rect 9824 10492 10272 10520
rect 10336 10492 10793 10520
rect 9824 10480 9830 10492
rect 10336 10464 10364 10492
rect 10781 10489 10793 10492
rect 10827 10489 10839 10523
rect 14001 10523 14059 10529
rect 14001 10520 14013 10523
rect 10781 10483 10839 10489
rect 10980 10492 12388 10520
rect 10226 10452 10232 10464
rect 8496 10424 10232 10452
rect 7984 10412 7990 10424
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 10318 10412 10324 10464
rect 10376 10412 10382 10464
rect 10410 10412 10416 10464
rect 10468 10452 10474 10464
rect 10597 10455 10655 10461
rect 10597 10452 10609 10455
rect 10468 10424 10609 10452
rect 10468 10412 10474 10424
rect 10597 10421 10609 10424
rect 10643 10421 10655 10455
rect 10597 10415 10655 10421
rect 10686 10412 10692 10464
rect 10744 10452 10750 10464
rect 10980 10452 11008 10492
rect 10744 10424 11008 10452
rect 11057 10455 11115 10461
rect 10744 10412 10750 10424
rect 11057 10421 11069 10455
rect 11103 10452 11115 10455
rect 11698 10452 11704 10464
rect 11103 10424 11704 10452
rect 11103 10421 11115 10424
rect 11057 10415 11115 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 12250 10452 12256 10464
rect 12211 10424 12256 10452
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 12360 10452 12388 10492
rect 13280 10492 14013 10520
rect 13280 10452 13308 10492
rect 14001 10489 14013 10492
rect 14047 10520 14059 10523
rect 14458 10520 14464 10532
rect 14047 10492 14464 10520
rect 14047 10489 14059 10492
rect 14001 10483 14059 10489
rect 14458 10480 14464 10492
rect 14516 10480 14522 10532
rect 16040 10492 17724 10520
rect 13722 10452 13728 10464
rect 12360 10424 13308 10452
rect 13683 10424 13728 10452
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 14645 10455 14703 10461
rect 14645 10421 14657 10455
rect 14691 10452 14703 10455
rect 16040 10452 16068 10492
rect 14691 10424 16068 10452
rect 14691 10421 14703 10424
rect 14645 10415 14703 10421
rect 16114 10412 16120 10464
rect 16172 10452 16178 10464
rect 16390 10452 16396 10464
rect 16172 10424 16396 10452
rect 16172 10412 16178 10424
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 17696 10452 17724 10492
rect 17770 10480 17776 10532
rect 17828 10520 17834 10532
rect 18601 10523 18659 10529
rect 18601 10520 18613 10523
rect 17828 10492 18613 10520
rect 17828 10480 17834 10492
rect 18601 10489 18613 10492
rect 18647 10489 18659 10523
rect 19628 10520 19656 10551
rect 20162 10548 20168 10560
rect 20220 10548 20226 10600
rect 20254 10548 20260 10600
rect 20312 10588 20318 10600
rect 20717 10591 20775 10597
rect 20717 10588 20729 10591
rect 20312 10560 20729 10588
rect 20312 10548 20318 10560
rect 20717 10557 20729 10560
rect 20763 10557 20775 10591
rect 20717 10551 20775 10557
rect 20809 10591 20867 10597
rect 20809 10557 20821 10591
rect 20855 10557 20867 10591
rect 20809 10551 20867 10557
rect 20824 10520 20852 10551
rect 19628 10492 20852 10520
rect 18601 10483 18659 10489
rect 20622 10452 20628 10464
rect 17696 10424 20628 10452
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 2958 10208 2964 10260
rect 3016 10248 3022 10260
rect 4709 10251 4767 10257
rect 3016 10220 3280 10248
rect 3016 10208 3022 10220
rect 1486 10072 1492 10124
rect 1544 10072 1550 10124
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 2038 10112 2044 10124
rect 1719 10084 2044 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 2038 10072 2044 10084
rect 2096 10072 2102 10124
rect 3252 10121 3280 10220
rect 4709 10217 4721 10251
rect 4755 10248 4767 10251
rect 4982 10248 4988 10260
rect 4755 10220 4988 10248
rect 4755 10217 4767 10220
rect 4709 10211 4767 10217
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5813 10251 5871 10257
rect 5813 10248 5825 10251
rect 5592 10220 5825 10248
rect 5592 10208 5598 10220
rect 5813 10217 5825 10220
rect 5859 10217 5871 10251
rect 7190 10248 7196 10260
rect 5813 10211 5871 10217
rect 5920 10220 7196 10248
rect 5920 10180 5948 10220
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 10413 10251 10471 10257
rect 10413 10248 10425 10251
rect 7300 10220 10425 10248
rect 6641 10183 6699 10189
rect 6641 10180 6653 10183
rect 3712 10152 5948 10180
rect 6012 10152 6653 10180
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10081 3295 10115
rect 3602 10112 3608 10124
rect 3563 10084 3608 10112
rect 3237 10075 3295 10081
rect 3602 10072 3608 10084
rect 3660 10072 3666 10124
rect 1504 10044 1532 10072
rect 1504 10016 3464 10044
rect 1489 9979 1547 9985
rect 1489 9945 1501 9979
rect 1535 9976 1547 9979
rect 1946 9976 1952 9988
rect 1535 9948 1952 9976
rect 1535 9945 1547 9948
rect 1489 9939 1547 9945
rect 1946 9936 1952 9948
rect 2004 9936 2010 9988
rect 2958 9976 2964 9988
rect 3016 9985 3022 9988
rect 3436 9985 3464 10016
rect 2928 9948 2964 9976
rect 2958 9936 2964 9948
rect 3016 9939 3028 9985
rect 3421 9979 3479 9985
rect 3421 9945 3433 9979
rect 3467 9945 3479 9979
rect 3421 9939 3479 9945
rect 3016 9936 3022 9939
rect 1854 9908 1860 9920
rect 1815 9880 1860 9908
rect 1854 9868 1860 9880
rect 1912 9868 1918 9920
rect 2038 9868 2044 9920
rect 2096 9908 2102 9920
rect 3712 9908 3740 10152
rect 5166 10072 5172 10124
rect 5224 10112 5230 10124
rect 5261 10115 5319 10121
rect 5261 10112 5273 10115
rect 5224 10084 5273 10112
rect 5224 10072 5230 10084
rect 5261 10081 5273 10084
rect 5307 10081 5319 10115
rect 5261 10075 5319 10081
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 6012 10112 6040 10152
rect 6641 10149 6653 10152
rect 6687 10149 6699 10183
rect 7098 10180 7104 10192
rect 7059 10152 7104 10180
rect 6641 10143 6699 10149
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 5500 10084 6040 10112
rect 6273 10115 6331 10121
rect 5500 10072 5506 10084
rect 6273 10081 6285 10115
rect 6319 10112 6331 10115
rect 6362 10112 6368 10124
rect 6319 10084 6368 10112
rect 6319 10081 6331 10084
rect 6273 10075 6331 10081
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 6457 10115 6515 10121
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 6546 10112 6552 10124
rect 6503 10084 6552 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 3786 10004 3792 10056
rect 3844 10044 3850 10056
rect 4062 10044 4068 10056
rect 3844 10016 3937 10044
rect 4023 10016 4068 10044
rect 3844 10004 3863 10016
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 4430 10004 4436 10056
rect 4488 10044 4494 10056
rect 5077 10047 5135 10053
rect 5077 10044 5089 10047
rect 4488 10016 5089 10044
rect 4488 10004 4494 10016
rect 5077 10013 5089 10016
rect 5123 10013 5135 10047
rect 6822 10044 6828 10056
rect 6783 10016 6828 10044
rect 5077 10007 5135 10013
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 3835 9976 3863 10004
rect 5442 9976 5448 9988
rect 3835 9948 5448 9976
rect 5442 9936 5448 9948
rect 5500 9936 5506 9988
rect 7300 9976 7328 10220
rect 10413 10217 10425 10220
rect 10459 10217 10471 10251
rect 10413 10211 10471 10217
rect 10870 10208 10876 10260
rect 10928 10248 10934 10260
rect 13541 10251 13599 10257
rect 10928 10220 12296 10248
rect 10928 10208 10934 10220
rect 9398 10180 9404 10192
rect 7392 10152 9404 10180
rect 7392 10121 7420 10152
rect 9398 10140 9404 10152
rect 9456 10180 9462 10192
rect 9674 10180 9680 10192
rect 9456 10152 9680 10180
rect 9456 10140 9462 10152
rect 9674 10140 9680 10152
rect 9732 10140 9738 10192
rect 12158 10180 12164 10192
rect 11992 10152 12164 10180
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10081 7435 10115
rect 7377 10075 7435 10081
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10112 8263 10115
rect 8386 10112 8392 10124
rect 8251 10084 8392 10112
rect 8251 10081 8263 10084
rect 8205 10075 8263 10081
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 9585 10115 9643 10121
rect 9585 10081 9597 10115
rect 9631 10112 9643 10115
rect 10502 10112 10508 10124
rect 9631 10084 10508 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10594 10072 10600 10124
rect 10652 10112 10658 10124
rect 11992 10121 12020 10152
rect 12158 10140 12164 10152
rect 12216 10140 12222 10192
rect 12268 10180 12296 10220
rect 13541 10217 13553 10251
rect 13587 10248 13599 10251
rect 14366 10248 14372 10260
rect 13587 10220 14372 10248
rect 13587 10217 13599 10220
rect 13541 10211 13599 10217
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 15657 10251 15715 10257
rect 15657 10217 15669 10251
rect 15703 10248 15715 10251
rect 16022 10248 16028 10260
rect 15703 10220 16028 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 16206 10248 16212 10260
rect 16167 10220 16212 10248
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 17678 10248 17684 10260
rect 17328 10220 17684 10248
rect 13817 10183 13875 10189
rect 13817 10180 13829 10183
rect 12268 10152 13829 10180
rect 13817 10149 13829 10152
rect 13863 10180 13875 10183
rect 14829 10183 14887 10189
rect 13863 10152 14412 10180
rect 13863 10149 13875 10152
rect 13817 10143 13875 10149
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 10652 10084 11253 10112
rect 10652 10072 10658 10084
rect 11241 10081 11253 10084
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 11977 10115 12035 10121
rect 11977 10081 11989 10115
rect 12023 10081 12035 10115
rect 11977 10075 12035 10081
rect 12069 10115 12127 10121
rect 12069 10081 12081 10115
rect 12115 10112 12127 10115
rect 12802 10112 12808 10124
rect 12115 10084 12808 10112
rect 12115 10081 12127 10084
rect 12069 10075 12127 10081
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10112 13047 10115
rect 13722 10112 13728 10124
rect 13035 10084 13728 10112
rect 13035 10081 13047 10084
rect 12989 10075 13047 10081
rect 13722 10072 13728 10084
rect 13780 10072 13786 10124
rect 14182 10112 14188 10124
rect 14143 10084 14188 10112
rect 14182 10072 14188 10084
rect 14240 10072 14246 10124
rect 14384 10121 14412 10152
rect 14829 10149 14841 10183
rect 14875 10180 14887 10183
rect 14875 10152 17172 10180
rect 14875 10149 14887 10152
rect 14829 10143 14887 10149
rect 14369 10115 14427 10121
rect 14369 10081 14381 10115
rect 14415 10081 14427 10115
rect 15010 10112 15016 10124
rect 14971 10084 15016 10112
rect 14369 10075 14427 10081
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 16577 10115 16635 10121
rect 16577 10112 16589 10115
rect 15120 10084 16589 10112
rect 7558 10004 7564 10056
rect 7616 10044 7622 10056
rect 7616 10016 7661 10044
rect 7616 10004 7622 10016
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 8662 10044 8668 10056
rect 8076 10016 8668 10044
rect 8076 10004 8082 10016
rect 8662 10004 8668 10016
rect 8720 10044 8726 10056
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8720 10016 8953 10044
rect 8720 10004 8726 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9030 10004 9036 10056
rect 9088 10044 9094 10056
rect 9088 10016 9812 10044
rect 9088 10004 9094 10016
rect 6564 9948 7328 9976
rect 2096 9880 3740 9908
rect 2096 9868 2102 9880
rect 4430 9868 4436 9920
rect 4488 9908 4494 9920
rect 5169 9911 5227 9917
rect 5169 9908 5181 9911
rect 4488 9880 5181 9908
rect 4488 9868 4494 9880
rect 5169 9877 5181 9880
rect 5215 9877 5227 9911
rect 5169 9871 5227 9877
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 5629 9911 5687 9917
rect 5629 9908 5641 9911
rect 5592 9880 5641 9908
rect 5592 9868 5598 9880
rect 5629 9877 5641 9880
rect 5675 9877 5687 9911
rect 5629 9871 5687 9877
rect 5810 9868 5816 9920
rect 5868 9908 5874 9920
rect 6181 9911 6239 9917
rect 6181 9908 6193 9911
rect 5868 9880 6193 9908
rect 5868 9868 5874 9880
rect 6181 9877 6193 9880
rect 6227 9877 6239 9911
rect 6181 9871 6239 9877
rect 6270 9868 6276 9920
rect 6328 9908 6334 9920
rect 6564 9908 6592 9948
rect 7834 9936 7840 9988
rect 7892 9976 7898 9988
rect 8846 9976 8852 9988
rect 7892 9948 8852 9976
rect 7892 9936 7898 9948
rect 8846 9936 8852 9948
rect 8904 9936 8910 9988
rect 9677 9979 9735 9985
rect 9677 9976 9689 9979
rect 9048 9948 9689 9976
rect 6328 9880 6592 9908
rect 6328 9868 6334 9880
rect 7374 9868 7380 9920
rect 7432 9908 7438 9920
rect 7469 9911 7527 9917
rect 7469 9908 7481 9911
rect 7432 9880 7481 9908
rect 7432 9868 7438 9880
rect 7469 9877 7481 9880
rect 7515 9877 7527 9911
rect 7469 9871 7527 9877
rect 7929 9911 7987 9917
rect 7929 9877 7941 9911
rect 7975 9908 7987 9911
rect 8297 9911 8355 9917
rect 8297 9908 8309 9911
rect 7975 9880 8309 9908
rect 7975 9877 7987 9880
rect 7929 9871 7987 9877
rect 8297 9877 8309 9880
rect 8343 9877 8355 9911
rect 8297 9871 8355 9877
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 8757 9911 8815 9917
rect 8444 9880 8489 9908
rect 8444 9868 8450 9880
rect 8757 9877 8769 9911
rect 8803 9908 8815 9911
rect 9048 9908 9076 9948
rect 9677 9945 9689 9948
rect 9723 9945 9735 9979
rect 9784 9976 9812 10016
rect 11882 10004 11888 10056
rect 11940 10044 11946 10056
rect 12621 10047 12679 10053
rect 12621 10044 12633 10047
rect 11940 10016 12633 10044
rect 11940 10004 11946 10016
rect 12621 10013 12633 10016
rect 12667 10013 12679 10047
rect 12621 10007 12679 10013
rect 12894 10004 12900 10056
rect 12952 10044 12958 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12952 10016 13185 10044
rect 12952 10004 12958 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10044 14519 10047
rect 14550 10044 14556 10056
rect 14507 10016 14556 10044
rect 14507 10013 14519 10016
rect 14461 10007 14519 10013
rect 14550 10004 14556 10016
rect 14608 10004 14614 10056
rect 10229 9979 10287 9985
rect 10229 9976 10241 9979
rect 9784 9948 10241 9976
rect 9677 9939 9735 9945
rect 10229 9945 10241 9948
rect 10275 9945 10287 9979
rect 11514 9976 11520 9988
rect 11475 9948 11520 9976
rect 10229 9939 10287 9945
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 13081 9979 13139 9985
rect 13081 9976 13093 9979
rect 12544 9948 13093 9976
rect 8803 9880 9076 9908
rect 9125 9911 9183 9917
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9214 9908 9220 9920
rect 9171 9880 9220 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 9309 9911 9367 9917
rect 9309 9877 9321 9911
rect 9355 9908 9367 9911
rect 9490 9908 9496 9920
rect 9355 9880 9496 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 9769 9911 9827 9917
rect 9769 9877 9781 9911
rect 9815 9908 9827 9911
rect 9858 9908 9864 9920
rect 9815 9880 9864 9908
rect 9815 9877 9827 9880
rect 9769 9871 9827 9877
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 10134 9908 10140 9920
rect 10095 9880 10140 9908
rect 10134 9868 10140 9880
rect 10192 9868 10198 9920
rect 10686 9908 10692 9920
rect 10647 9880 10692 9908
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 11054 9908 11060 9920
rect 11015 9880 11060 9908
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 12158 9908 12164 9920
rect 11204 9880 11249 9908
rect 12119 9880 12164 9908
rect 11204 9868 11210 9880
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 12544 9917 12572 9948
rect 13081 9945 13093 9948
rect 13127 9945 13139 9979
rect 13081 9939 13139 9945
rect 14182 9936 14188 9988
rect 14240 9976 14246 9988
rect 15120 9976 15148 10084
rect 16577 10081 16589 10084
rect 16623 10112 16635 10115
rect 16623 10084 16896 10112
rect 16623 10081 16635 10084
rect 16577 10075 16635 10081
rect 15286 10044 15292 10056
rect 15247 10016 15292 10044
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 15746 10044 15752 10056
rect 15707 10016 15752 10044
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 16206 10004 16212 10056
rect 16264 10044 16270 10056
rect 16761 10047 16819 10053
rect 16761 10044 16773 10047
rect 16264 10016 16773 10044
rect 16264 10004 16270 10016
rect 16761 10013 16773 10016
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 14240 9948 15148 9976
rect 15304 9976 15332 10004
rect 16025 9979 16083 9985
rect 16025 9976 16037 9979
rect 15304 9948 16037 9976
rect 14240 9936 14246 9948
rect 16025 9945 16037 9948
rect 16071 9945 16083 9979
rect 16868 9976 16896 10084
rect 17144 10044 17172 10152
rect 17328 10124 17356 10220
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 18690 10248 18696 10260
rect 18651 10220 18696 10248
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 19610 10208 19616 10260
rect 19668 10248 19674 10260
rect 19886 10248 19892 10260
rect 19668 10220 19892 10248
rect 19668 10208 19674 10220
rect 19886 10208 19892 10220
rect 19944 10208 19950 10260
rect 20254 10248 20260 10260
rect 20215 10220 20260 10248
rect 20254 10208 20260 10220
rect 20312 10208 20318 10260
rect 17310 10112 17316 10124
rect 17223 10084 17316 10112
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 18708 10112 18736 10208
rect 19334 10140 19340 10192
rect 19392 10180 19398 10192
rect 20438 10180 20444 10192
rect 19392 10152 20444 10180
rect 19392 10140 19398 10152
rect 20438 10140 20444 10152
rect 20496 10140 20502 10192
rect 20625 10183 20683 10189
rect 20625 10149 20637 10183
rect 20671 10180 20683 10183
rect 21266 10180 21272 10192
rect 20671 10152 21272 10180
rect 20671 10149 20683 10152
rect 20625 10143 20683 10149
rect 21266 10140 21272 10152
rect 21324 10140 21330 10192
rect 19610 10112 19616 10124
rect 18708 10084 19616 10112
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 20806 10112 20812 10124
rect 19904 10084 20812 10112
rect 19702 10044 19708 10056
rect 17144 10016 19708 10044
rect 19702 10004 19708 10016
rect 19760 10004 19766 10056
rect 19904 10053 19932 10084
rect 20806 10072 20812 10084
rect 20864 10072 20870 10124
rect 20990 10112 20996 10124
rect 20951 10084 20996 10112
rect 20990 10072 20996 10084
rect 21048 10072 21054 10124
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10013 19947 10047
rect 19889 10007 19947 10013
rect 20622 10004 20628 10056
rect 20680 10044 20686 10056
rect 20717 10047 20775 10053
rect 20717 10044 20729 10047
rect 20680 10016 20729 10044
rect 20680 10004 20686 10016
rect 20717 10013 20729 10016
rect 20763 10013 20775 10047
rect 20717 10007 20775 10013
rect 17558 9979 17616 9985
rect 17558 9976 17570 9979
rect 16868 9948 17570 9976
rect 16025 9939 16083 9945
rect 17558 9945 17570 9948
rect 17604 9976 17616 9979
rect 17678 9976 17684 9988
rect 17604 9948 17684 9976
rect 17604 9945 17616 9948
rect 17558 9939 17616 9945
rect 17678 9936 17684 9948
rect 17736 9936 17742 9988
rect 17770 9936 17776 9988
rect 17828 9976 17834 9988
rect 18785 9979 18843 9985
rect 18785 9976 18797 9979
rect 17828 9948 18797 9976
rect 17828 9936 17834 9948
rect 18785 9945 18797 9948
rect 18831 9945 18843 9979
rect 18966 9976 18972 9988
rect 18927 9948 18972 9976
rect 18785 9939 18843 9945
rect 18966 9936 18972 9948
rect 19024 9936 19030 9988
rect 19429 9979 19487 9985
rect 19429 9945 19441 9979
rect 19475 9976 19487 9979
rect 20346 9976 20352 9988
rect 19475 9948 20352 9976
rect 19475 9945 19487 9948
rect 19429 9939 19487 9945
rect 20346 9936 20352 9948
rect 20404 9936 20410 9988
rect 20438 9936 20444 9988
rect 20496 9976 20502 9988
rect 20496 9948 20541 9976
rect 20496 9936 20502 9948
rect 12529 9911 12587 9917
rect 12529 9877 12541 9911
rect 12575 9877 12587 9911
rect 12529 9871 12587 9877
rect 12618 9868 12624 9920
rect 12676 9908 12682 9920
rect 13633 9911 13691 9917
rect 13633 9908 13645 9911
rect 12676 9880 13645 9908
rect 12676 9868 12682 9880
rect 13633 9877 13645 9880
rect 13679 9908 13691 9911
rect 13906 9908 13912 9920
rect 13679 9880 13912 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 15010 9908 15016 9920
rect 14792 9880 15016 9908
rect 14792 9868 14798 9880
rect 15010 9868 15016 9880
rect 15068 9868 15074 9920
rect 15197 9911 15255 9917
rect 15197 9877 15209 9911
rect 15243 9908 15255 9911
rect 15470 9908 15476 9920
rect 15243 9880 15476 9908
rect 15243 9877 15255 9880
rect 15197 9871 15255 9877
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 15933 9911 15991 9917
rect 15933 9877 15945 9911
rect 15979 9908 15991 9911
rect 16298 9908 16304 9920
rect 15979 9880 16304 9908
rect 15979 9877 15991 9880
rect 15933 9871 15991 9877
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 16853 9911 16911 9917
rect 16853 9877 16865 9911
rect 16899 9908 16911 9911
rect 17126 9908 17132 9920
rect 16899 9880 17132 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 17126 9868 17132 9880
rect 17184 9868 17190 9920
rect 17221 9911 17279 9917
rect 17221 9877 17233 9911
rect 17267 9908 17279 9911
rect 17862 9908 17868 9920
rect 17267 9880 17868 9908
rect 17267 9877 17279 9880
rect 17221 9871 17279 9877
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 19150 9868 19156 9920
rect 19208 9908 19214 9920
rect 19797 9911 19855 9917
rect 19797 9908 19809 9911
rect 19208 9880 19809 9908
rect 19208 9868 19214 9880
rect 19797 9877 19809 9880
rect 19843 9877 19855 9911
rect 19797 9871 19855 9877
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 1581 9707 1639 9713
rect 1581 9673 1593 9707
rect 1627 9704 1639 9707
rect 1762 9704 1768 9716
rect 1627 9676 1768 9704
rect 1627 9673 1639 9676
rect 1581 9667 1639 9673
rect 1762 9664 1768 9676
rect 1820 9664 1826 9716
rect 2130 9664 2136 9716
rect 2188 9704 2194 9716
rect 3326 9704 3332 9716
rect 2188 9676 3332 9704
rect 2188 9664 2194 9676
rect 3326 9664 3332 9676
rect 3384 9664 3390 9716
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 4617 9707 4675 9713
rect 4617 9704 4629 9707
rect 4396 9676 4629 9704
rect 4396 9664 4402 9676
rect 4617 9673 4629 9676
rect 4663 9673 4675 9707
rect 4617 9667 4675 9673
rect 5350 9664 5356 9716
rect 5408 9704 5414 9716
rect 6178 9704 6184 9716
rect 5408 9676 6184 9704
rect 5408 9664 5414 9676
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 7098 9704 7104 9716
rect 6748 9676 7104 9704
rect 3786 9596 3792 9648
rect 3844 9645 3850 9648
rect 3844 9636 3856 9645
rect 3844 9608 3889 9636
rect 3844 9599 3856 9608
rect 3844 9596 3850 9599
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 6748 9645 6776 9676
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 7561 9707 7619 9713
rect 7561 9673 7573 9707
rect 7607 9704 7619 9707
rect 7742 9704 7748 9716
rect 7607 9676 7748 9704
rect 7607 9673 7619 9676
rect 7561 9667 7619 9673
rect 7742 9664 7748 9676
rect 7800 9664 7806 9716
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 9585 9707 9643 9713
rect 9585 9704 9597 9707
rect 8444 9676 9597 9704
rect 8444 9664 8450 9676
rect 9585 9673 9597 9676
rect 9631 9673 9643 9707
rect 9585 9667 9643 9673
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 10505 9707 10563 9713
rect 10505 9704 10517 9707
rect 9824 9676 10517 9704
rect 9824 9664 9830 9676
rect 10505 9673 10517 9676
rect 10551 9704 10563 9707
rect 10778 9704 10784 9716
rect 10551 9676 10784 9704
rect 10551 9673 10563 9676
rect 10505 9667 10563 9673
rect 10778 9664 10784 9676
rect 10836 9704 10842 9716
rect 10873 9707 10931 9713
rect 10873 9704 10885 9707
rect 10836 9676 10885 9704
rect 10836 9664 10842 9676
rect 10873 9673 10885 9676
rect 10919 9673 10931 9707
rect 10873 9667 10931 9673
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 11333 9707 11391 9713
rect 11333 9704 11345 9707
rect 11112 9676 11345 9704
rect 11112 9664 11118 9676
rect 11333 9673 11345 9676
rect 11379 9673 11391 9707
rect 11333 9667 11391 9673
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 11882 9704 11888 9716
rect 11756 9676 11888 9704
rect 11756 9664 11762 9676
rect 11882 9664 11888 9676
rect 11940 9664 11946 9716
rect 11977 9707 12035 9713
rect 11977 9673 11989 9707
rect 12023 9704 12035 9707
rect 12250 9704 12256 9716
rect 12023 9676 12256 9704
rect 12023 9673 12035 9676
rect 11977 9667 12035 9673
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 12802 9664 12808 9716
rect 12860 9704 12866 9716
rect 13078 9704 13084 9716
rect 12860 9676 13084 9704
rect 12860 9664 12866 9676
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 13265 9707 13323 9713
rect 13265 9673 13277 9707
rect 13311 9704 13323 9707
rect 19150 9704 19156 9716
rect 13311 9676 19156 9704
rect 13311 9673 13323 9676
rect 13265 9667 13323 9673
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 19521 9707 19579 9713
rect 19521 9673 19533 9707
rect 19567 9704 19579 9707
rect 19794 9704 19800 9716
rect 19567 9676 19800 9704
rect 19567 9673 19579 9676
rect 19521 9667 19579 9673
rect 19794 9664 19800 9676
rect 19852 9664 19858 9716
rect 20162 9664 20168 9716
rect 20220 9704 20226 9716
rect 20349 9707 20407 9713
rect 20349 9704 20361 9707
rect 20220 9676 20361 9704
rect 20220 9664 20226 9676
rect 20349 9673 20361 9676
rect 20395 9673 20407 9707
rect 20349 9667 20407 9673
rect 6733 9639 6791 9645
rect 5592 9608 6592 9636
rect 5592 9596 5598 9608
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 4522 9568 4528 9580
rect 4203 9540 4528 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9568 5135 9571
rect 5123 9540 5764 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 1854 9500 1860 9512
rect 1815 9472 1860 9500
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 2130 9500 2136 9512
rect 1995 9472 2136 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9500 4123 9503
rect 4246 9500 4252 9512
rect 4111 9472 4252 9500
rect 4111 9469 4123 9472
rect 4065 9463 4123 9469
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 4338 9460 4344 9512
rect 4396 9500 4402 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 4396 9472 4445 9500
rect 4396 9460 4402 9472
rect 4433 9469 4445 9472
rect 4479 9500 4491 9503
rect 4890 9500 4896 9512
rect 4479 9472 4896 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 2406 9432 2412 9444
rect 2367 9404 2412 9432
rect 2406 9392 2412 9404
rect 2464 9392 2470 9444
rect 2685 9435 2743 9441
rect 2685 9432 2697 9435
rect 2516 9404 2697 9432
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 2516 9364 2544 9404
rect 2685 9401 2697 9404
rect 2731 9432 2743 9435
rect 2958 9432 2964 9444
rect 2731 9404 2964 9432
rect 2731 9401 2743 9404
rect 2685 9395 2743 9401
rect 2958 9392 2964 9404
rect 3016 9392 3022 9444
rect 4798 9432 4804 9444
rect 4080 9404 4804 9432
rect 1728 9336 2544 9364
rect 2593 9367 2651 9373
rect 1728 9324 1734 9336
rect 2593 9333 2605 9367
rect 2639 9364 2651 9367
rect 2866 9364 2872 9376
rect 2639 9336 2872 9364
rect 2639 9333 2651 9336
rect 2593 9327 2651 9333
rect 2866 9324 2872 9336
rect 2924 9324 2930 9376
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 4080 9364 4108 9404
rect 4798 9392 4804 9404
rect 4856 9392 4862 9444
rect 5000 9432 5028 9531
rect 5166 9500 5172 9512
rect 5127 9472 5172 9500
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 5445 9435 5503 9441
rect 5445 9432 5457 9435
rect 5000 9404 5457 9432
rect 5445 9401 5457 9404
rect 5491 9401 5503 9435
rect 5736 9432 5764 9540
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 6564 9568 6592 9608
rect 6733 9605 6745 9639
rect 6779 9605 6791 9639
rect 6733 9599 6791 9605
rect 7834 9596 7840 9648
rect 7892 9636 7898 9648
rect 7892 9608 9251 9636
rect 7892 9596 7898 9608
rect 6822 9568 6828 9580
rect 5868 9540 5913 9568
rect 6564 9540 6828 9568
rect 5868 9528 5874 9540
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 7650 9568 7656 9580
rect 7611 9540 7656 9568
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7926 9528 7932 9580
rect 7984 9568 7990 9580
rect 8386 9577 8392 9580
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 7984 9540 8125 9568
rect 7984 9528 7990 9540
rect 8113 9537 8125 9540
rect 8159 9537 8171 9571
rect 8369 9571 8392 9577
rect 8369 9568 8381 9571
rect 8113 9531 8171 9537
rect 8220 9540 8381 9568
rect 5902 9500 5908 9512
rect 5863 9472 5908 9500
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 6089 9503 6147 9509
rect 6089 9469 6101 9503
rect 6135 9500 6147 9503
rect 6270 9500 6276 9512
rect 6135 9472 6276 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 6270 9460 6276 9472
rect 6328 9500 6334 9512
rect 6932 9500 6960 9528
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 6328 9472 7021 9500
rect 6328 9460 6334 9472
rect 7009 9469 7021 9472
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 7469 9503 7527 9509
rect 7469 9500 7481 9503
rect 7432 9472 7481 9500
rect 7432 9460 7438 9472
rect 7469 9469 7481 9472
rect 7515 9500 7527 9503
rect 8220 9500 8248 9540
rect 8369 9537 8381 9540
rect 8369 9531 8392 9537
rect 8386 9528 8392 9531
rect 8444 9528 8450 9580
rect 9223 9568 9251 9608
rect 9306 9596 9312 9648
rect 9364 9636 9370 9648
rect 12069 9639 12127 9645
rect 9364 9608 11836 9636
rect 9364 9596 9370 9608
rect 9582 9568 9588 9580
rect 9223 9540 9588 9568
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9824 9540 9965 9568
rect 9824 9528 9830 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 10965 9571 11023 9577
rect 10965 9537 10977 9571
rect 11011 9568 11023 9571
rect 11698 9568 11704 9580
rect 11011 9540 11704 9568
rect 11011 9537 11023 9540
rect 10965 9531 11023 9537
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 11808 9568 11836 9608
rect 12069 9605 12081 9639
rect 12115 9636 12127 9639
rect 12434 9636 12440 9648
rect 12115 9608 12440 9636
rect 12115 9605 12127 9608
rect 12069 9599 12127 9605
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 13722 9645 13728 9648
rect 13716 9636 13728 9645
rect 12636 9608 13584 9636
rect 13683 9608 13728 9636
rect 12526 9568 12532 9580
rect 11808 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 7515 9472 8248 9500
rect 10045 9503 10103 9509
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 10045 9469 10057 9503
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9469 10195 9503
rect 10137 9463 10195 9469
rect 6365 9435 6423 9441
rect 6365 9432 6377 9435
rect 5736 9404 6377 9432
rect 5445 9395 5503 9401
rect 6365 9401 6377 9404
rect 6411 9401 6423 9435
rect 10060 9432 10088 9463
rect 6365 9395 6423 9401
rect 9048 9404 10088 9432
rect 4338 9364 4344 9376
rect 3108 9336 4108 9364
rect 4299 9336 4344 9364
rect 3108 9324 3114 9336
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 7926 9364 7932 9376
rect 7616 9336 7932 9364
rect 7616 9324 7622 9336
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 8021 9367 8079 9373
rect 8021 9333 8033 9367
rect 8067 9364 8079 9367
rect 9048 9364 9076 9404
rect 8067 9336 9076 9364
rect 9493 9367 9551 9373
rect 8067 9333 8079 9336
rect 8021 9327 8079 9333
rect 9493 9333 9505 9367
rect 9539 9364 9551 9367
rect 9674 9364 9680 9376
rect 9539 9336 9680 9364
rect 9539 9333 9551 9336
rect 9493 9327 9551 9333
rect 9674 9324 9680 9336
rect 9732 9364 9738 9376
rect 10152 9364 10180 9463
rect 10502 9460 10508 9512
rect 10560 9500 10566 9512
rect 10689 9503 10747 9509
rect 10689 9500 10701 9503
rect 10560 9472 10701 9500
rect 10560 9460 10566 9472
rect 10689 9469 10701 9472
rect 10735 9469 10747 9503
rect 11790 9500 11796 9512
rect 11751 9472 11796 9500
rect 10689 9463 10747 9469
rect 11790 9460 11796 9472
rect 11848 9460 11854 9512
rect 12636 9509 12664 9608
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 12768 9540 12909 9568
rect 12768 9528 12774 9540
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 13170 9528 13176 9580
rect 13228 9528 13234 9580
rect 13556 9568 13584 9608
rect 13716 9599 13728 9608
rect 13722 9596 13728 9599
rect 13780 9596 13786 9648
rect 14458 9596 14464 9648
rect 14516 9636 14522 9648
rect 17586 9645 17592 9648
rect 17558 9639 17592 9645
rect 17558 9636 17570 9639
rect 14516 9608 17570 9636
rect 14516 9596 14522 9608
rect 17558 9605 17570 9608
rect 17558 9599 17592 9605
rect 17586 9596 17592 9599
rect 17644 9596 17650 9648
rect 17678 9596 17684 9648
rect 17736 9596 17742 9648
rect 17862 9596 17868 9648
rect 17920 9636 17926 9648
rect 19981 9639 20039 9645
rect 19981 9636 19993 9639
rect 17920 9608 19993 9636
rect 17920 9596 17926 9608
rect 19981 9605 19993 9608
rect 20027 9605 20039 9639
rect 19981 9599 20039 9605
rect 20438 9596 20444 9648
rect 20496 9636 20502 9648
rect 20990 9636 20996 9648
rect 20496 9608 20996 9636
rect 20496 9596 20502 9608
rect 20990 9596 20996 9608
rect 21048 9596 21054 9648
rect 21266 9596 21272 9648
rect 21324 9636 21330 9648
rect 21453 9639 21511 9645
rect 21453 9636 21465 9639
rect 21324 9608 21465 9636
rect 21324 9596 21330 9608
rect 21453 9605 21465 9608
rect 21499 9605 21511 9639
rect 21453 9599 21511 9605
rect 14182 9568 14188 9580
rect 13556 9540 14188 9568
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 14550 9528 14556 9580
rect 14608 9568 14614 9580
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 14608 9540 15301 9568
rect 14608 9528 14614 9540
rect 15289 9537 15301 9540
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 17034 9568 17040 9580
rect 16163 9540 17040 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 17034 9528 17040 9540
rect 17092 9528 17098 9580
rect 17126 9528 17132 9580
rect 17184 9528 17190 9580
rect 17221 9571 17279 9577
rect 17221 9537 17233 9571
rect 17267 9568 17279 9571
rect 17310 9568 17316 9580
rect 17267 9540 17316 9568
rect 17267 9537 17279 9540
rect 17221 9531 17279 9537
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 17696 9568 17724 9596
rect 18785 9571 18843 9577
rect 18785 9568 18797 9571
rect 17696 9540 18797 9568
rect 18785 9537 18797 9540
rect 18831 9537 18843 9571
rect 18785 9531 18843 9537
rect 18969 9571 19027 9577
rect 18969 9537 18981 9571
rect 19015 9568 19027 9571
rect 19334 9568 19340 9580
rect 19015 9540 19340 9568
rect 19015 9537 19027 9540
rect 18969 9531 19027 9537
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9469 12679 9503
rect 12621 9463 12679 9469
rect 12805 9503 12863 9509
rect 12805 9469 12817 9503
rect 12851 9500 12863 9503
rect 13078 9500 13084 9512
rect 12851 9472 13084 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 12158 9392 12164 9444
rect 12216 9432 12222 9444
rect 12437 9435 12495 9441
rect 12437 9432 12449 9435
rect 12216 9404 12449 9432
rect 12216 9392 12222 9404
rect 12437 9401 12449 9404
rect 12483 9401 12495 9435
rect 13188 9432 13216 9528
rect 13446 9500 13452 9512
rect 13407 9472 13452 9500
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 15102 9500 15108 9512
rect 15063 9472 15108 9500
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9500 15255 9503
rect 15470 9500 15476 9512
rect 15243 9472 15476 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 15470 9460 15476 9472
rect 15528 9460 15534 9512
rect 15930 9500 15936 9512
rect 15891 9472 15936 9500
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 16025 9503 16083 9509
rect 16025 9469 16037 9503
rect 16071 9469 16083 9503
rect 16025 9463 16083 9469
rect 13354 9432 13360 9444
rect 13188 9404 13360 9432
rect 12437 9395 12495 9401
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 14918 9392 14924 9444
rect 14976 9432 14982 9444
rect 16040 9432 16068 9463
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 17144 9500 17172 9528
rect 16724 9472 17172 9500
rect 16724 9460 16730 9472
rect 14976 9404 16068 9432
rect 16485 9435 16543 9441
rect 14976 9392 14982 9404
rect 16485 9401 16497 9435
rect 16531 9432 16543 9435
rect 17126 9432 17132 9444
rect 16531 9404 17132 9432
rect 16531 9401 16543 9404
rect 16485 9395 16543 9401
rect 17126 9392 17132 9404
rect 17184 9392 17190 9444
rect 18693 9435 18751 9441
rect 18693 9401 18705 9435
rect 18739 9432 18751 9435
rect 18984 9432 19012 9531
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 19484 9540 19529 9568
rect 19484 9528 19490 9540
rect 19702 9528 19708 9580
rect 19760 9528 19766 9580
rect 19794 9528 19800 9580
rect 19852 9568 19858 9580
rect 19889 9571 19947 9577
rect 19889 9568 19901 9571
rect 19852 9540 19901 9568
rect 19852 9528 19858 9540
rect 19889 9537 19901 9540
rect 19935 9537 19947 9571
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 19889 9531 19947 9537
rect 19996 9540 20729 9568
rect 19720 9500 19748 9528
rect 19996 9500 20024 9540
rect 20717 9537 20729 9540
rect 20763 9537 20775 9571
rect 20717 9531 20775 9537
rect 19720 9472 20024 9500
rect 20073 9503 20131 9509
rect 20073 9469 20085 9503
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 18739 9404 19012 9432
rect 18739 9401 18751 9404
rect 18693 9395 18751 9401
rect 19610 9392 19616 9444
rect 19668 9432 19674 9444
rect 20088 9432 20116 9463
rect 20254 9460 20260 9512
rect 20312 9500 20318 9512
rect 20438 9500 20444 9512
rect 20312 9472 20444 9500
rect 20312 9460 20318 9472
rect 20438 9460 20444 9472
rect 20496 9460 20502 9512
rect 20806 9500 20812 9512
rect 20767 9472 20812 9500
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 20901 9503 20959 9509
rect 20901 9469 20913 9503
rect 20947 9469 20959 9503
rect 20901 9463 20959 9469
rect 20622 9432 20628 9444
rect 19668 9404 20628 9432
rect 19668 9392 19674 9404
rect 20622 9392 20628 9404
rect 20680 9432 20686 9444
rect 20916 9432 20944 9463
rect 20680 9404 20944 9432
rect 20680 9392 20686 9404
rect 21082 9392 21088 9444
rect 21140 9432 21146 9444
rect 21269 9435 21327 9441
rect 21269 9432 21281 9435
rect 21140 9404 21281 9432
rect 21140 9392 21146 9404
rect 21269 9401 21281 9404
rect 21315 9401 21327 9435
rect 21269 9395 21327 9401
rect 9732 9336 10180 9364
rect 9732 9324 9738 9336
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 10468 9336 11529 9364
rect 10468 9324 10474 9336
rect 11517 9333 11529 9336
rect 11563 9364 11575 9367
rect 12710 9364 12716 9376
rect 11563 9336 12716 9364
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 14792 9336 14841 9364
rect 14792 9324 14798 9336
rect 14829 9333 14841 9336
rect 14875 9333 14887 9367
rect 14829 9327 14887 9333
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 15344 9336 15669 9364
rect 15344 9324 15350 9336
rect 15657 9333 15669 9336
rect 15703 9333 15715 9367
rect 16666 9364 16672 9376
rect 16627 9336 16672 9364
rect 15657 9327 15715 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 16853 9367 16911 9373
rect 16853 9364 16865 9367
rect 16816 9336 16865 9364
rect 16816 9324 16822 9336
rect 16853 9333 16865 9336
rect 16899 9333 16911 9367
rect 16853 9327 16911 9333
rect 17037 9367 17095 9373
rect 17037 9333 17049 9367
rect 17083 9364 17095 9367
rect 17218 9364 17224 9376
rect 17083 9336 17224 9364
rect 17083 9333 17095 9336
rect 17037 9327 17095 9333
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 18782 9324 18788 9376
rect 18840 9364 18846 9376
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 18840 9336 19257 9364
rect 18840 9324 18846 9336
rect 19245 9333 19257 9336
rect 19291 9333 19303 9367
rect 19245 9327 19303 9333
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 2130 9160 2136 9172
rect 2091 9132 2136 9160
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 3418 9160 3424 9172
rect 3283 9132 3424 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 3936 9132 4077 9160
rect 3936 9120 3942 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 4212 9132 5304 9160
rect 4212 9120 4218 9132
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 2682 9092 2688 9104
rect 2556 9064 2688 9092
rect 2556 9052 2562 9064
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 3605 9095 3663 9101
rect 3605 9061 3617 9095
rect 3651 9092 3663 9095
rect 3970 9092 3976 9104
rect 3651 9064 3976 9092
rect 3651 9061 3663 9064
rect 3605 9055 3663 9061
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 5166 9092 5172 9104
rect 4632 9064 5172 9092
rect 1581 9027 1639 9033
rect 1581 8993 1593 9027
rect 1627 9024 1639 9027
rect 1670 9024 1676 9036
rect 1627 8996 1676 9024
rect 1627 8993 1639 8996
rect 1581 8987 1639 8993
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 2406 8984 2412 9036
rect 2464 9024 2470 9036
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 2464 8996 2881 9024
rect 2464 8984 2470 8996
rect 2869 8993 2881 8996
rect 2915 9024 2927 9027
rect 4062 9024 4068 9036
rect 2915 8996 4068 9024
rect 2915 8993 2927 8996
rect 2869 8987 2927 8993
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4632 9033 4660 9064
rect 5166 9052 5172 9064
rect 5224 9052 5230 9104
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 4172 8996 4629 9024
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 2682 8956 2688 8968
rect 2639 8928 2688 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 3418 8956 3424 8968
rect 3379 8928 3424 8956
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 1673 8891 1731 8897
rect 1673 8857 1685 8891
rect 1719 8888 1731 8891
rect 1719 8860 2268 8888
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 2240 8829 2268 8860
rect 2958 8848 2964 8900
rect 3016 8888 3022 8900
rect 4172 8888 4200 8996
rect 4617 8993 4629 8996
rect 4663 8993 4675 9027
rect 5276 9024 5304 9132
rect 5902 9120 5908 9172
rect 5960 9160 5966 9172
rect 6638 9160 6644 9172
rect 5960 9132 6644 9160
rect 5960 9120 5966 9132
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 7374 9160 7380 9172
rect 7335 9132 7380 9160
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 7800 9132 8953 9160
rect 7800 9120 7806 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 9122 9160 9128 9172
rect 9083 9132 9128 9160
rect 8941 9123 8999 9129
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 9401 9163 9459 9169
rect 9401 9129 9413 9163
rect 9447 9160 9459 9163
rect 9582 9160 9588 9172
rect 9447 9132 9588 9160
rect 9447 9129 9459 9132
rect 9401 9123 9459 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 10229 9163 10287 9169
rect 10229 9129 10241 9163
rect 10275 9160 10287 9163
rect 11054 9160 11060 9172
rect 10275 9132 11060 9160
rect 10275 9129 10287 9132
rect 10229 9123 10287 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 13078 9160 13084 9172
rect 13039 9132 13084 9160
rect 13078 9120 13084 9132
rect 13136 9120 13142 9172
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 13228 9132 13273 9160
rect 13228 9120 13234 9132
rect 13814 9120 13820 9172
rect 13872 9160 13878 9172
rect 14550 9160 14556 9172
rect 13872 9132 14556 9160
rect 13872 9120 13878 9132
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 15930 9120 15936 9172
rect 15988 9160 15994 9172
rect 16209 9163 16267 9169
rect 16209 9160 16221 9163
rect 15988 9132 16221 9160
rect 15988 9120 15994 9132
rect 16209 9129 16221 9132
rect 16255 9129 16267 9163
rect 16209 9123 16267 9129
rect 10321 9095 10379 9101
rect 10321 9061 10333 9095
rect 10367 9092 10379 9095
rect 10594 9092 10600 9104
rect 10367 9064 10600 9092
rect 10367 9061 10379 9064
rect 10321 9055 10379 9061
rect 10594 9052 10600 9064
rect 10652 9052 10658 9104
rect 11698 9052 11704 9104
rect 11756 9092 11762 9104
rect 14458 9092 14464 9104
rect 11756 9064 11836 9092
rect 11756 9052 11762 9064
rect 5350 9024 5356 9036
rect 5263 8996 5356 9024
rect 4617 8987 4675 8993
rect 5350 8984 5356 8996
rect 5408 9024 5414 9036
rect 5445 9027 5503 9033
rect 5445 9024 5457 9027
rect 5408 8996 5457 9024
rect 5408 8984 5414 8996
rect 5445 8993 5457 8996
rect 5491 8993 5503 9027
rect 6270 9024 6276 9036
rect 6231 8996 6276 9024
rect 5445 8987 5503 8993
rect 6270 8984 6276 8996
rect 6328 9024 6334 9036
rect 6638 9024 6644 9036
rect 6328 8996 6644 9024
rect 6328 8984 6334 8996
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 6788 8996 7113 9024
rect 6788 8984 6794 8996
rect 7101 8993 7113 8996
rect 7147 8993 7159 9027
rect 7101 8987 7159 8993
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 10502 9024 10508 9036
rect 9723 8996 10508 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 11808 9033 11836 9064
rect 12452 9064 14464 9092
rect 12452 9033 12480 9064
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 11793 9027 11851 9033
rect 11793 8993 11805 9027
rect 11839 8993 11851 9027
rect 11793 8987 11851 8993
rect 12437 9027 12495 9033
rect 12437 8993 12449 9027
rect 12483 8993 12495 9027
rect 12618 9024 12624 9036
rect 12579 8996 12624 9024
rect 12437 8987 12495 8993
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 13354 9024 13360 9036
rect 12820 8996 13360 9024
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8956 4491 8959
rect 5166 8956 5172 8968
rect 4479 8928 5172 8956
rect 4479 8925 4491 8928
rect 4433 8919 4491 8925
rect 5166 8916 5172 8928
rect 5224 8916 5230 8968
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 6086 8956 6092 8968
rect 5316 8928 5361 8956
rect 6047 8928 6092 8956
rect 5316 8916 5322 8928
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8956 6975 8959
rect 7466 8956 7472 8968
rect 6963 8928 7472 8956
rect 6963 8925 6975 8928
rect 6917 8919 6975 8925
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 8662 8956 8668 8968
rect 7800 8928 8668 8956
rect 7800 8916 7806 8928
rect 8662 8916 8668 8928
rect 8720 8956 8726 8968
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 8720 8928 8769 8956
rect 8720 8916 8726 8928
rect 8757 8925 8769 8928
rect 8803 8925 8815 8959
rect 8757 8919 8815 8925
rect 9582 8916 9588 8968
rect 9640 8956 9646 8968
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 9640 8928 9781 8956
rect 9640 8916 9646 8928
rect 9769 8925 9781 8928
rect 9815 8925 9827 8959
rect 10520 8956 10548 8984
rect 11146 8956 11152 8968
rect 10520 8928 11152 8956
rect 9769 8919 9827 8925
rect 11146 8916 11152 8928
rect 11204 8956 11210 8968
rect 11434 8959 11492 8965
rect 11434 8956 11446 8959
rect 11204 8928 11446 8956
rect 11204 8916 11210 8928
rect 11434 8925 11446 8928
rect 11480 8925 11492 8959
rect 11698 8956 11704 8968
rect 11659 8928 11704 8956
rect 11434 8919 11492 8925
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 12820 8956 12848 8996
rect 13354 8984 13360 8996
rect 13412 9024 13418 9036
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13412 8996 13645 9024
rect 13412 8984 13418 8996
rect 13633 8993 13645 8996
rect 13679 8993 13691 9027
rect 13633 8987 13691 8993
rect 14274 8984 14280 9036
rect 14332 9024 14338 9036
rect 14829 9027 14887 9033
rect 14829 9024 14841 9027
rect 14332 8996 14841 9024
rect 14332 8984 14338 8996
rect 14829 8993 14841 8996
rect 14875 8993 14887 9027
rect 16224 9024 16252 9123
rect 17034 9120 17040 9172
rect 17092 9160 17098 9172
rect 17773 9163 17831 9169
rect 17773 9160 17785 9163
rect 17092 9132 17785 9160
rect 17092 9120 17098 9132
rect 17773 9129 17785 9132
rect 17819 9129 17831 9163
rect 17773 9123 17831 9129
rect 18874 9120 18880 9172
rect 18932 9160 18938 9172
rect 19061 9163 19119 9169
rect 19061 9160 19073 9163
rect 18932 9132 19073 9160
rect 18932 9120 18938 9132
rect 19061 9129 19073 9132
rect 19107 9129 19119 9163
rect 20714 9160 20720 9172
rect 20675 9132 20720 9160
rect 19061 9123 19119 9129
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 17494 9052 17500 9104
rect 17552 9092 17558 9104
rect 18046 9092 18052 9104
rect 17552 9064 18052 9092
rect 17552 9052 17558 9064
rect 18046 9052 18052 9064
rect 18104 9052 18110 9104
rect 18601 9095 18659 9101
rect 18601 9092 18613 9095
rect 18248 9064 18613 9092
rect 18248 9033 18276 9064
rect 18601 9061 18613 9064
rect 18647 9061 18659 9095
rect 18601 9055 18659 9061
rect 18233 9027 18291 9033
rect 18233 9024 18245 9027
rect 16224 8996 16436 9024
rect 14829 8987 14887 8993
rect 12584 8928 12848 8956
rect 12584 8916 12590 8928
rect 12894 8916 12900 8968
rect 12952 8956 12958 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 12952 8928 13461 8956
rect 12952 8916 12958 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 13817 8959 13875 8965
rect 13817 8956 13829 8959
rect 13780 8928 13829 8956
rect 13780 8916 13786 8928
rect 13817 8925 13829 8928
rect 13863 8956 13875 8959
rect 14369 8959 14427 8965
rect 14369 8956 14381 8959
rect 13863 8928 14381 8956
rect 13863 8925 13875 8928
rect 13817 8919 13875 8925
rect 14369 8925 14381 8928
rect 14415 8956 14427 8959
rect 15470 8956 15476 8968
rect 14415 8928 15476 8956
rect 14415 8925 14427 8928
rect 14369 8919 14427 8925
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 16298 8956 16304 8968
rect 16259 8928 16304 8956
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 16408 8956 16436 8996
rect 17328 8996 18245 9024
rect 16557 8959 16615 8965
rect 16557 8956 16569 8959
rect 16408 8928 16569 8956
rect 16557 8925 16569 8928
rect 16603 8925 16615 8959
rect 16557 8919 16615 8925
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17328 8956 17356 8996
rect 18233 8993 18245 8996
rect 18279 8993 18291 9027
rect 18233 8987 18291 8993
rect 18417 9027 18475 9033
rect 18417 8993 18429 9027
rect 18463 9024 18475 9027
rect 18463 8996 19380 9024
rect 18463 8993 18475 8996
rect 18417 8987 18475 8993
rect 18432 8956 18460 8987
rect 19352 8968 19380 8996
rect 20622 8984 20628 9036
rect 20680 9024 20686 9036
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 20680 8996 21281 9024
rect 20680 8984 20686 8996
rect 21269 8993 21281 8996
rect 21315 8993 21327 9027
rect 21269 8987 21327 8993
rect 18874 8956 18880 8968
rect 17092 8928 17356 8956
rect 17420 8928 18460 8956
rect 18835 8928 18880 8956
rect 17092 8916 17098 8928
rect 3016 8860 4200 8888
rect 4525 8891 4583 8897
rect 3016 8848 3022 8860
rect 4525 8857 4537 8891
rect 4571 8888 4583 8891
rect 6564 8888 6592 8916
rect 7926 8888 7932 8900
rect 4571 8860 5764 8888
rect 6564 8860 7932 8888
rect 4571 8857 4583 8860
rect 4525 8851 4583 8857
rect 2225 8823 2283 8829
rect 2225 8789 2237 8823
rect 2271 8789 2283 8823
rect 2225 8783 2283 8789
rect 2498 8780 2504 8832
rect 2556 8820 2562 8832
rect 2685 8823 2743 8829
rect 2685 8820 2697 8823
rect 2556 8792 2697 8820
rect 2556 8780 2562 8792
rect 2685 8789 2697 8792
rect 2731 8789 2743 8823
rect 2685 8783 2743 8789
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3384 8792 3801 8820
rect 3384 8780 3390 8792
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 4798 8780 4804 8832
rect 4856 8820 4862 8832
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 4856 8792 4905 8820
rect 4856 8780 4862 8792
rect 4893 8789 4905 8792
rect 4939 8789 4951 8823
rect 4893 8783 4951 8789
rect 5353 8823 5411 8829
rect 5353 8789 5365 8823
rect 5399 8820 5411 8823
rect 5534 8820 5540 8832
rect 5399 8792 5540 8820
rect 5399 8789 5411 8792
rect 5353 8783 5411 8789
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 5736 8829 5764 8860
rect 7926 8848 7932 8860
rect 7984 8848 7990 8900
rect 8501 8891 8559 8897
rect 8501 8857 8513 8891
rect 8547 8888 8559 8891
rect 9674 8888 9680 8900
rect 8547 8860 9680 8888
rect 8547 8857 8559 8860
rect 8501 8851 8559 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 9858 8888 9864 8900
rect 9819 8860 9864 8888
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 12161 8891 12219 8897
rect 12161 8857 12173 8891
rect 12207 8857 12219 8891
rect 12161 8851 12219 8857
rect 5721 8823 5779 8829
rect 5721 8789 5733 8823
rect 5767 8789 5779 8823
rect 5721 8783 5779 8789
rect 6181 8823 6239 8829
rect 6181 8789 6193 8823
rect 6227 8820 6239 8823
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 6227 8792 6561 8820
rect 6227 8789 6239 8792
rect 6181 8783 6239 8789
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 6549 8783 6607 8789
rect 6822 8780 6828 8832
rect 6880 8820 6886 8832
rect 7009 8823 7067 8829
rect 7009 8820 7021 8823
rect 6880 8792 7021 8820
rect 6880 8780 6886 8792
rect 7009 8789 7021 8792
rect 7055 8789 7067 8823
rect 7009 8783 7067 8789
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 9490 8820 9496 8832
rect 8076 8792 9496 8820
rect 8076 8780 8082 8792
rect 9490 8780 9496 8792
rect 9548 8820 9554 8832
rect 12176 8820 12204 8851
rect 12250 8848 12256 8900
rect 12308 8888 12314 8900
rect 15102 8897 15108 8900
rect 12308 8860 14679 8888
rect 12308 8848 12314 8860
rect 12713 8823 12771 8829
rect 12713 8820 12725 8823
rect 9548 8792 12725 8820
rect 9548 8780 9554 8792
rect 12713 8789 12725 8792
rect 12759 8820 12771 8823
rect 13170 8820 13176 8832
rect 12759 8792 13176 8820
rect 12759 8789 12771 8792
rect 12713 8783 12771 8789
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13446 8780 13452 8832
rect 13504 8820 13510 8832
rect 14090 8820 14096 8832
rect 13504 8792 14096 8820
rect 13504 8780 13510 8792
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 14185 8823 14243 8829
rect 14185 8789 14197 8823
rect 14231 8820 14243 8823
rect 14550 8820 14556 8832
rect 14231 8792 14556 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 14651 8820 14679 8860
rect 15096 8851 15108 8897
rect 15160 8888 15166 8900
rect 17420 8888 17448 8928
rect 18874 8916 18880 8928
rect 18932 8916 18938 8968
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 19116 8928 19257 8956
rect 19116 8916 19122 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 19334 8916 19340 8968
rect 19392 8916 19398 8968
rect 19518 8965 19524 8968
rect 19512 8919 19524 8965
rect 19576 8956 19582 8968
rect 19576 8928 19612 8956
rect 19518 8916 19524 8919
rect 19576 8916 19582 8928
rect 19426 8888 19432 8900
rect 15160 8860 17448 8888
rect 17481 8860 19432 8888
rect 15102 8848 15108 8851
rect 15160 8848 15166 8860
rect 17481 8820 17509 8860
rect 19426 8848 19432 8860
rect 19484 8848 19490 8900
rect 17678 8820 17684 8832
rect 14651 8792 17509 8820
rect 17639 8792 17684 8820
rect 17678 8780 17684 8792
rect 17736 8780 17742 8832
rect 18138 8820 18144 8832
rect 18099 8792 18144 8820
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 19334 8780 19340 8832
rect 19392 8820 19398 8832
rect 20530 8820 20536 8832
rect 19392 8792 20536 8820
rect 19392 8780 19398 8792
rect 20530 8780 20536 8792
rect 20588 8820 20594 8832
rect 20625 8823 20683 8829
rect 20625 8820 20637 8823
rect 20588 8792 20637 8820
rect 20588 8780 20594 8792
rect 20625 8789 20637 8792
rect 20671 8789 20683 8823
rect 21082 8820 21088 8832
rect 21043 8792 21088 8820
rect 20625 8783 20683 8789
rect 21082 8780 21088 8792
rect 21140 8780 21146 8832
rect 21174 8780 21180 8832
rect 21232 8820 21238 8832
rect 21232 8792 21277 8820
rect 21232 8780 21238 8792
rect 22002 8780 22008 8832
rect 22060 8820 22066 8832
rect 22060 8792 22140 8820
rect 22060 8780 22066 8792
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 2317 8619 2375 8625
rect 2317 8616 2329 8619
rect 2188 8588 2329 8616
rect 2188 8576 2194 8588
rect 2317 8585 2329 8588
rect 2363 8616 2375 8619
rect 3421 8619 3479 8625
rect 2363 8588 3372 8616
rect 2363 8585 2375 8588
rect 2317 8579 2375 8585
rect 3344 8548 3372 8588
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 3467 8588 3893 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 3881 8579 3939 8585
rect 3973 8619 4031 8625
rect 3973 8585 3985 8619
rect 4019 8616 4031 8619
rect 4341 8619 4399 8625
rect 4341 8616 4353 8619
rect 4019 8588 4353 8616
rect 4019 8585 4031 8588
rect 3973 8579 4031 8585
rect 4341 8585 4353 8588
rect 4387 8585 4399 8619
rect 4341 8579 4399 8585
rect 4709 8619 4767 8625
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 4890 8616 4896 8628
rect 4755 8588 4896 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5166 8616 5172 8628
rect 5127 8588 5172 8616
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 5537 8619 5595 8625
rect 5537 8616 5549 8619
rect 5316 8588 5549 8616
rect 5316 8576 5322 8588
rect 5537 8585 5549 8588
rect 5583 8616 5595 8619
rect 6270 8616 6276 8628
rect 5583 8588 6276 8616
rect 5583 8585 5595 8588
rect 5537 8579 5595 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6365 8619 6423 8625
rect 6365 8585 6377 8619
rect 6411 8616 6423 8619
rect 6638 8616 6644 8628
rect 6411 8588 6644 8616
rect 6411 8585 6423 8588
rect 6365 8579 6423 8585
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 7929 8619 7987 8625
rect 7929 8616 7941 8619
rect 7340 8588 7941 8616
rect 7340 8576 7346 8588
rect 7929 8585 7941 8588
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 8757 8619 8815 8625
rect 8757 8616 8769 8619
rect 8168 8588 8769 8616
rect 8168 8576 8174 8588
rect 8757 8585 8769 8588
rect 8803 8585 8815 8619
rect 8757 8579 8815 8585
rect 8846 8576 8852 8628
rect 8904 8616 8910 8628
rect 9125 8619 9183 8625
rect 8904 8588 9076 8616
rect 8904 8576 8910 8588
rect 4614 8548 4620 8560
rect 3344 8520 4620 8548
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 5629 8551 5687 8557
rect 5629 8517 5641 8551
rect 5675 8548 5687 8551
rect 5994 8548 6000 8560
rect 5675 8520 6000 8548
rect 5675 8517 5687 8520
rect 5629 8511 5687 8517
rect 5994 8508 6000 8520
rect 6052 8548 6058 8560
rect 8297 8551 8355 8557
rect 6052 8520 6132 8548
rect 6052 8508 6058 8520
rect 1394 8480 1400 8492
rect 1355 8452 1400 8480
rect 1394 8440 1400 8452
rect 1452 8440 1458 8492
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8480 2283 8483
rect 2866 8480 2872 8492
rect 2271 8452 2872 8480
rect 2271 8449 2283 8452
rect 2225 8443 2283 8449
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3234 8480 3240 8492
rect 3099 8452 3240 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 4798 8440 4804 8492
rect 4856 8480 4862 8492
rect 4856 8452 4901 8480
rect 4856 8440 4862 8452
rect 2406 8372 2412 8424
rect 2464 8412 2470 8424
rect 2464 8384 2509 8412
rect 2464 8372 2470 8384
rect 2590 8372 2596 8424
rect 2648 8412 2654 8424
rect 2648 8384 2737 8412
rect 2648 8372 2654 8384
rect 2709 8344 2737 8384
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 2958 8412 2964 8424
rect 2832 8384 2877 8412
rect 2919 8384 2964 8412
rect 2832 8372 2838 8384
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 3878 8372 3884 8424
rect 3936 8412 3942 8424
rect 4065 8415 4123 8421
rect 4065 8412 4077 8415
rect 3936 8384 4077 8412
rect 3936 8372 3942 8384
rect 4065 8381 4077 8384
rect 4111 8381 4123 8415
rect 4893 8415 4951 8421
rect 4893 8412 4905 8415
rect 4065 8375 4123 8381
rect 4172 8384 4905 8412
rect 3513 8347 3571 8353
rect 3513 8344 3525 8347
rect 2709 8316 3525 8344
rect 3513 8313 3525 8316
rect 3559 8313 3571 8347
rect 3513 8307 3571 8313
rect 1854 8276 1860 8288
rect 1815 8248 1860 8276
rect 1854 8236 1860 8248
rect 1912 8236 1918 8288
rect 2866 8236 2872 8288
rect 2924 8276 2930 8288
rect 4062 8276 4068 8288
rect 2924 8248 4068 8276
rect 2924 8236 2930 8248
rect 4062 8236 4068 8248
rect 4120 8276 4126 8288
rect 4172 8276 4200 8384
rect 4893 8381 4905 8384
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 5442 8372 5448 8424
rect 5500 8412 5506 8424
rect 5721 8415 5779 8421
rect 5721 8412 5733 8415
rect 5500 8384 5733 8412
rect 5500 8372 5506 8384
rect 5721 8381 5733 8384
rect 5767 8381 5779 8415
rect 6104 8412 6132 8520
rect 6196 8520 7696 8548
rect 6196 8489 6224 8520
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 7478 8483 7536 8489
rect 7478 8480 7490 8483
rect 6788 8452 7490 8480
rect 6788 8440 6794 8452
rect 7478 8449 7490 8452
rect 7524 8449 7536 8483
rect 7478 8443 7536 8449
rect 6546 8412 6552 8424
rect 6104 8384 6552 8412
rect 5721 8375 5779 8381
rect 6546 8372 6552 8384
rect 6604 8372 6610 8424
rect 7668 8412 7696 8520
rect 8297 8517 8309 8551
rect 8343 8548 8355 8551
rect 8938 8548 8944 8560
rect 8343 8520 8944 8548
rect 8343 8517 8355 8520
rect 8297 8511 8355 8517
rect 8938 8508 8944 8520
rect 8996 8508 9002 8560
rect 9048 8548 9076 8588
rect 9125 8585 9137 8619
rect 9171 8616 9183 8619
rect 9398 8616 9404 8628
rect 9171 8588 9404 8616
rect 9171 8585 9183 8588
rect 9125 8579 9183 8585
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9585 8619 9643 8625
rect 9585 8585 9597 8619
rect 9631 8616 9643 8619
rect 9674 8616 9680 8628
rect 9631 8588 9680 8616
rect 9631 8585 9643 8588
rect 9585 8579 9643 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 11609 8619 11667 8625
rect 11609 8616 11621 8619
rect 10100 8588 11621 8616
rect 10100 8576 10106 8588
rect 11609 8585 11621 8588
rect 11655 8616 11667 8619
rect 11790 8616 11796 8628
rect 11655 8588 11796 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 12710 8616 12716 8628
rect 12671 8588 12716 8616
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 13265 8619 13323 8625
rect 13265 8616 13277 8619
rect 13228 8588 13277 8616
rect 13228 8576 13234 8588
rect 13265 8585 13277 8588
rect 13311 8616 13323 8619
rect 13722 8616 13728 8628
rect 13311 8588 13728 8616
rect 13311 8585 13323 8588
rect 13265 8579 13323 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14553 8619 14611 8625
rect 14553 8616 14565 8619
rect 14056 8588 14565 8616
rect 14056 8576 14062 8588
rect 14553 8585 14565 8588
rect 14599 8585 14611 8619
rect 14918 8616 14924 8628
rect 14879 8588 14924 8616
rect 14553 8579 14611 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15286 8576 15292 8628
rect 15344 8616 15350 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 15344 8588 16037 8616
rect 15344 8576 15350 8588
rect 16025 8585 16037 8588
rect 16071 8585 16083 8619
rect 16025 8579 16083 8585
rect 16485 8619 16543 8625
rect 16485 8585 16497 8619
rect 16531 8616 16543 8619
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 16531 8588 16957 8616
rect 16531 8585 16543 8588
rect 16485 8579 16543 8585
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 16945 8579 17003 8585
rect 17037 8619 17095 8625
rect 17037 8585 17049 8619
rect 17083 8616 17095 8619
rect 17126 8616 17132 8628
rect 17083 8588 17132 8616
rect 17083 8585 17095 8588
rect 17037 8579 17095 8585
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 17402 8616 17408 8628
rect 17363 8588 17408 8616
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17681 8619 17739 8625
rect 17681 8585 17693 8619
rect 17727 8616 17739 8619
rect 18138 8616 18144 8628
rect 17727 8588 18144 8616
rect 17727 8585 17739 8588
rect 17681 8579 17739 8585
rect 18138 8576 18144 8588
rect 18196 8576 18202 8628
rect 19426 8616 19432 8628
rect 19387 8588 19432 8616
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 19702 8576 19708 8628
rect 19760 8616 19766 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 19760 8588 20085 8616
rect 19760 8576 19766 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 20073 8579 20131 8585
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20441 8619 20499 8625
rect 20441 8616 20453 8619
rect 20404 8588 20453 8616
rect 20404 8576 20410 8588
rect 20441 8585 20453 8588
rect 20487 8585 20499 8619
rect 20441 8579 20499 8585
rect 20714 8576 20720 8628
rect 20772 8616 20778 8628
rect 20993 8619 21051 8625
rect 20993 8616 21005 8619
rect 20772 8588 21005 8616
rect 20772 8576 20778 8588
rect 20993 8585 21005 8588
rect 21039 8585 21051 8619
rect 22112 8616 22140 8792
rect 20993 8579 21051 8585
rect 21468 8588 22140 8616
rect 9217 8551 9275 8557
rect 9217 8548 9229 8551
rect 9048 8520 9229 8548
rect 9217 8517 9229 8520
rect 9263 8548 9275 8551
rect 9263 8520 10548 8548
rect 9263 8517 9275 8520
rect 9217 8511 9275 8517
rect 9490 8480 9496 8492
rect 8516 8452 9496 8480
rect 7742 8412 7748 8424
rect 7668 8384 7748 8412
rect 7742 8372 7748 8384
rect 7800 8412 7806 8424
rect 8389 8415 8447 8421
rect 7800 8384 7893 8412
rect 7800 8372 7806 8384
rect 8389 8381 8401 8415
rect 8435 8381 8447 8415
rect 8516 8412 8544 8452
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 10520 8480 10548 8520
rect 10594 8508 10600 8560
rect 10652 8548 10658 8560
rect 10698 8551 10756 8557
rect 10698 8548 10710 8551
rect 10652 8520 10710 8548
rect 10652 8508 10658 8520
rect 10698 8517 10710 8520
rect 10744 8517 10756 8551
rect 10698 8511 10756 8517
rect 10870 8508 10876 8560
rect 10928 8548 10934 8560
rect 11149 8551 11207 8557
rect 11149 8548 11161 8551
rect 10928 8520 11161 8548
rect 10928 8508 10934 8520
rect 11149 8517 11161 8520
rect 11195 8548 11207 8551
rect 12250 8548 12256 8560
rect 11195 8520 12256 8548
rect 11195 8517 11207 8520
rect 11149 8511 11207 8517
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 11241 8483 11299 8489
rect 11241 8480 11253 8483
rect 10520 8452 11253 8480
rect 11241 8449 11253 8452
rect 11287 8480 11299 8483
rect 11330 8480 11336 8492
rect 11287 8452 11336 8480
rect 11287 8449 11299 8452
rect 11241 8443 11299 8449
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 12158 8480 12164 8492
rect 12119 8452 12164 8480
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 12728 8480 12756 8576
rect 14461 8551 14519 8557
rect 14461 8548 14473 8551
rect 14016 8520 14473 8548
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12728 8452 12909 8480
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13044 8452 13645 8480
rect 13044 8440 13050 8452
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 8389 8375 8447 8381
rect 8496 8384 8544 8412
rect 8573 8415 8631 8421
rect 4798 8304 4804 8356
rect 4856 8344 4862 8356
rect 4856 8316 6868 8344
rect 4856 8304 4862 8316
rect 4120 8248 4200 8276
rect 4120 8236 4126 8248
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5997 8279 6055 8285
rect 5997 8276 6009 8279
rect 5224 8248 6009 8276
rect 5224 8236 5230 8248
rect 5997 8245 6009 8248
rect 6043 8245 6055 8279
rect 6840 8276 6868 8316
rect 8110 8304 8116 8356
rect 8168 8344 8174 8356
rect 8404 8344 8432 8375
rect 8496 8344 8524 8384
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 8662 8412 8668 8424
rect 8619 8384 8668 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 8662 8372 8668 8384
rect 8720 8412 8726 8424
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 8720 8384 9321 8412
rect 8720 8372 8726 8384
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 10965 8415 11023 8421
rect 10965 8381 10977 8415
rect 11011 8412 11023 8415
rect 11698 8412 11704 8424
rect 11011 8384 11704 8412
rect 11011 8381 11023 8384
rect 10965 8375 11023 8381
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 12250 8412 12256 8424
rect 12211 8384 12256 8412
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 12345 8415 12403 8421
rect 12345 8381 12357 8415
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 9582 8344 9588 8356
rect 8168 8316 8524 8344
rect 8864 8316 9588 8344
rect 8168 8304 8174 8316
rect 7466 8276 7472 8288
rect 6840 8248 7472 8276
rect 5997 8239 6055 8245
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 7558 8236 7564 8288
rect 7616 8276 7622 8288
rect 8864 8276 8892 8316
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 12360 8344 12388 8375
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 13170 8412 13176 8424
rect 12492 8384 13176 8412
rect 12492 8372 12498 8384
rect 13170 8372 13176 8384
rect 13228 8372 13234 8424
rect 13538 8412 13544 8424
rect 13499 8384 13544 8412
rect 13538 8372 13544 8384
rect 13596 8412 13602 8424
rect 14016 8412 14044 8520
rect 14461 8517 14473 8520
rect 14507 8517 14519 8551
rect 14461 8511 14519 8517
rect 15381 8551 15439 8557
rect 15381 8517 15393 8551
rect 15427 8548 15439 8551
rect 15470 8548 15476 8560
rect 15427 8520 15476 8548
rect 15427 8517 15439 8520
rect 15381 8511 15439 8517
rect 15470 8508 15476 8520
rect 15528 8508 15534 8560
rect 15657 8551 15715 8557
rect 15657 8517 15669 8551
rect 15703 8548 15715 8551
rect 17954 8548 17960 8560
rect 15703 8520 17960 8548
rect 15703 8517 15715 8520
rect 15657 8511 15715 8517
rect 17954 8508 17960 8520
rect 18012 8508 18018 8560
rect 18966 8508 18972 8560
rect 19024 8557 19030 8560
rect 19024 8548 19036 8557
rect 19024 8520 19069 8548
rect 19024 8511 19036 8520
rect 19024 8508 19030 8511
rect 19150 8508 19156 8560
rect 19208 8548 19214 8560
rect 21085 8551 21143 8557
rect 21085 8548 21097 8551
rect 19208 8520 21097 8548
rect 19208 8508 19214 8520
rect 21085 8517 21097 8520
rect 21131 8548 21143 8551
rect 21266 8548 21272 8560
rect 21131 8520 21272 8548
rect 21131 8517 21143 8520
rect 21085 8511 21143 8517
rect 21266 8508 21272 8520
rect 21324 8508 21330 8560
rect 14090 8440 14096 8492
rect 14148 8480 14154 8492
rect 14148 8452 16068 8480
rect 14148 8440 14154 8452
rect 13596 8384 14044 8412
rect 14277 8415 14335 8421
rect 13596 8372 13602 8384
rect 14277 8381 14289 8415
rect 14323 8381 14335 8415
rect 15010 8412 15016 8424
rect 14971 8384 15016 8412
rect 14277 8375 14335 8381
rect 11204 8316 12388 8344
rect 11204 8304 11210 8316
rect 13078 8304 13084 8356
rect 13136 8344 13142 8356
rect 13136 8316 13181 8344
rect 13136 8304 13142 8316
rect 13814 8304 13820 8356
rect 13872 8344 13878 8356
rect 14292 8344 14320 8375
rect 15010 8372 15016 8384
rect 15068 8372 15074 8424
rect 15930 8412 15936 8424
rect 15891 8384 15936 8412
rect 15930 8372 15936 8384
rect 15988 8372 15994 8424
rect 16040 8412 16068 8452
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 16172 8452 16217 8480
rect 16172 8440 16178 8452
rect 17494 8440 17500 8492
rect 17552 8480 17558 8492
rect 19245 8483 19303 8489
rect 19245 8480 19257 8483
rect 17552 8452 19257 8480
rect 17552 8440 17558 8452
rect 19245 8449 19257 8452
rect 19291 8449 19303 8483
rect 19245 8443 19303 8449
rect 19521 8483 19579 8489
rect 19521 8449 19533 8483
rect 19567 8480 19579 8483
rect 19610 8480 19616 8492
rect 19567 8452 19616 8480
rect 19567 8449 19579 8452
rect 19521 8443 19579 8449
rect 19610 8440 19616 8452
rect 19668 8440 19674 8492
rect 19886 8480 19892 8492
rect 19847 8452 19892 8480
rect 19886 8440 19892 8452
rect 19944 8440 19950 8492
rect 21468 8489 21496 8588
rect 21453 8483 21511 8489
rect 21453 8449 21465 8483
rect 21499 8449 21511 8483
rect 21453 8443 21511 8449
rect 16298 8412 16304 8424
rect 16040 8384 16304 8412
rect 16298 8372 16304 8384
rect 16356 8372 16362 8424
rect 16853 8415 16911 8421
rect 16853 8381 16865 8415
rect 16899 8412 16911 8415
rect 17034 8412 17040 8424
rect 16899 8384 17040 8412
rect 16899 8381 16911 8384
rect 16853 8375 16911 8381
rect 17034 8372 17040 8384
rect 17092 8412 17098 8424
rect 17678 8412 17684 8424
rect 17092 8384 17684 8412
rect 17092 8372 17098 8384
rect 17678 8372 17684 8384
rect 17736 8372 17742 8424
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 19705 8415 19763 8421
rect 19705 8412 19717 8415
rect 19392 8384 19717 8412
rect 19392 8372 19398 8384
rect 19705 8381 19717 8384
rect 19751 8381 19763 8415
rect 19705 8375 19763 8381
rect 20438 8372 20444 8424
rect 20496 8412 20502 8424
rect 20533 8415 20591 8421
rect 20533 8412 20545 8415
rect 20496 8384 20545 8412
rect 20496 8372 20502 8384
rect 20533 8381 20545 8384
rect 20579 8381 20591 8415
rect 20533 8375 20591 8381
rect 20625 8415 20683 8421
rect 20625 8381 20637 8415
rect 20671 8412 20683 8415
rect 20714 8412 20720 8424
rect 20671 8384 20720 8412
rect 20671 8381 20683 8384
rect 20625 8375 20683 8381
rect 20714 8372 20720 8384
rect 20772 8412 20778 8424
rect 21358 8412 21364 8424
rect 20772 8384 21364 8412
rect 20772 8372 20778 8384
rect 21358 8372 21364 8384
rect 21416 8372 21422 8424
rect 15102 8344 15108 8356
rect 13872 8316 13917 8344
rect 14292 8316 15108 8344
rect 13872 8304 13878 8316
rect 15102 8304 15108 8316
rect 15160 8304 15166 8356
rect 15194 8304 15200 8356
rect 15252 8344 15258 8356
rect 17126 8344 17132 8356
rect 15252 8316 17132 8344
rect 15252 8304 15258 8316
rect 17126 8304 17132 8316
rect 17184 8304 17190 8356
rect 17586 8304 17592 8356
rect 17644 8344 17650 8356
rect 17865 8347 17923 8353
rect 17865 8344 17877 8347
rect 17644 8316 17877 8344
rect 17644 8304 17650 8316
rect 17865 8313 17877 8316
rect 17911 8313 17923 8347
rect 21468 8344 21496 8443
rect 17865 8307 17923 8313
rect 19260 8316 21496 8344
rect 7616 8248 8892 8276
rect 7616 8236 7622 8248
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 9950 8276 9956 8288
rect 9088 8248 9956 8276
rect 9088 8236 9094 8248
rect 9950 8236 9956 8248
rect 10008 8236 10014 8288
rect 11790 8276 11796 8288
rect 11751 8248 11796 8276
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 13909 8279 13967 8285
rect 13909 8276 13921 8279
rect 13044 8248 13921 8276
rect 13044 8236 13050 8248
rect 13909 8245 13921 8248
rect 13955 8245 13967 8279
rect 13909 8239 13967 8245
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 15212 8276 15240 8304
rect 14608 8248 15240 8276
rect 14608 8236 14614 8248
rect 17218 8236 17224 8288
rect 17276 8276 17282 8288
rect 17494 8276 17500 8288
rect 17276 8248 17500 8276
rect 17276 8236 17282 8248
rect 17494 8236 17500 8248
rect 17552 8236 17558 8288
rect 17678 8236 17684 8288
rect 17736 8276 17742 8288
rect 19260 8276 19288 8316
rect 21358 8276 21364 8288
rect 17736 8248 19288 8276
rect 21319 8248 21364 8276
rect 17736 8236 17742 8248
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2409 8075 2467 8081
rect 2409 8072 2421 8075
rect 2096 8044 2421 8072
rect 2096 8032 2102 8044
rect 2409 8041 2421 8044
rect 2455 8041 2467 8075
rect 2409 8035 2467 8041
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 2958 8072 2964 8084
rect 2915 8044 2964 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 4890 8032 4896 8084
rect 4948 8072 4954 8084
rect 5261 8075 5319 8081
rect 5261 8072 5273 8075
rect 4948 8044 5273 8072
rect 4948 8032 4954 8044
rect 5261 8041 5273 8044
rect 5307 8041 5319 8075
rect 5261 8035 5319 8041
rect 5810 8032 5816 8084
rect 5868 8072 5874 8084
rect 6086 8072 6092 8084
rect 5868 8044 5948 8072
rect 6047 8044 6092 8072
rect 5868 8032 5874 8044
rect 14 7964 20 8016
rect 72 8004 78 8016
rect 934 8004 940 8016
rect 72 7976 940 8004
rect 72 7964 78 7976
rect 934 7964 940 7976
rect 992 7964 998 8016
rect 1118 7964 1124 8016
rect 1176 8004 1182 8016
rect 2777 8007 2835 8013
rect 1176 7976 2084 8004
rect 1176 7964 1182 7976
rect 1670 7896 1676 7948
rect 1728 7936 1734 7948
rect 1765 7939 1823 7945
rect 1765 7936 1777 7939
rect 1728 7908 1777 7936
rect 1728 7896 1734 7908
rect 1765 7905 1777 7908
rect 1811 7905 1823 7939
rect 1765 7899 1823 7905
rect 1854 7896 1860 7948
rect 1912 7936 1918 7948
rect 1949 7939 2007 7945
rect 1949 7936 1961 7939
rect 1912 7908 1961 7936
rect 1912 7896 1918 7908
rect 1949 7905 1961 7908
rect 1995 7905 2007 7939
rect 2056 7936 2084 7976
rect 2777 7973 2789 8007
rect 2823 8004 2835 8007
rect 3142 8004 3148 8016
rect 2823 7976 3148 8004
rect 2823 7973 2835 7976
rect 2777 7967 2835 7973
rect 3142 7964 3148 7976
rect 3200 7964 3206 8016
rect 5350 7964 5356 8016
rect 5408 8004 5414 8016
rect 5920 8004 5948 8044
rect 6086 8032 6092 8044
rect 6144 8032 6150 8084
rect 7193 8075 7251 8081
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7374 8072 7380 8084
rect 7239 8044 7380 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 7374 8032 7380 8044
rect 7432 8072 7438 8084
rect 10410 8072 10416 8084
rect 7432 8044 10416 8072
rect 7432 8032 7438 8044
rect 6917 8007 6975 8013
rect 6917 8004 6929 8007
rect 5408 7976 5856 8004
rect 5920 7976 6929 8004
rect 5408 7964 5414 7976
rect 2958 7936 2964 7948
rect 2056 7908 2964 7936
rect 1949 7899 2007 7905
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 3513 7939 3571 7945
rect 3513 7905 3525 7939
rect 3559 7936 3571 7939
rect 3602 7936 3608 7948
rect 3559 7908 3608 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 3602 7896 3608 7908
rect 3660 7936 3666 7948
rect 4154 7936 4160 7948
rect 3660 7908 4160 7936
rect 3660 7896 3666 7908
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 5828 7945 5856 7976
rect 6917 7973 6929 7976
rect 6963 8004 6975 8007
rect 7282 8004 7288 8016
rect 6963 7976 7288 8004
rect 6963 7973 6975 7976
rect 6917 7967 6975 7973
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 7466 7964 7472 8016
rect 7524 8004 7530 8016
rect 7524 7976 8156 8004
rect 7524 7964 7530 7976
rect 5813 7939 5871 7945
rect 5813 7905 5825 7939
rect 5859 7905 5871 7939
rect 5813 7899 5871 7905
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 1486 7868 1492 7880
rect 1443 7840 1492 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 1486 7828 1492 7840
rect 1544 7828 1550 7880
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2866 7868 2872 7880
rect 2639 7840 2872 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2866 7828 2872 7840
rect 2924 7868 2930 7880
rect 3970 7868 3976 7880
rect 2924 7840 3976 7868
rect 2924 7828 2930 7840
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4902 7871 4960 7877
rect 4902 7868 4914 7871
rect 4120 7840 4914 7868
rect 4120 7828 4126 7840
rect 4902 7837 4914 7840
rect 4948 7837 4960 7871
rect 5166 7868 5172 7880
rect 5127 7840 5172 7868
rect 4902 7831 4960 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 5718 7868 5724 7880
rect 5408 7840 5724 7868
rect 5408 7828 5414 7840
rect 5718 7828 5724 7840
rect 5776 7868 5782 7880
rect 6656 7868 6684 7899
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 8018 7936 8024 7948
rect 6880 7908 8024 7936
rect 6880 7896 6886 7908
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 8128 7945 8156 7976
rect 8113 7939 8171 7945
rect 8113 7905 8125 7939
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 7098 7868 7104 7880
rect 5776 7840 6684 7868
rect 7059 7840 7104 7868
rect 5776 7828 5782 7840
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 7558 7828 7564 7880
rect 7616 7828 7622 7880
rect 7834 7868 7840 7880
rect 7795 7840 7840 7868
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 8036 7868 8064 7896
rect 8384 7877 8412 8044
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 11146 8072 11152 8084
rect 10836 8044 11152 8072
rect 10836 8032 10842 8044
rect 11146 8032 11152 8044
rect 11204 8072 11210 8084
rect 11425 8075 11483 8081
rect 11425 8072 11437 8075
rect 11204 8044 11437 8072
rect 11204 8032 11210 8044
rect 11425 8041 11437 8044
rect 11471 8041 11483 8075
rect 11425 8035 11483 8041
rect 11698 8032 11704 8084
rect 11756 8072 11762 8084
rect 12986 8072 12992 8084
rect 11756 8044 12992 8072
rect 11756 8032 11762 8044
rect 8757 8007 8815 8013
rect 8757 7973 8769 8007
rect 8803 8004 8815 8007
rect 9030 8004 9036 8016
rect 8803 7976 9036 8004
rect 8803 7973 8815 7976
rect 8757 7967 8815 7973
rect 9030 7964 9036 7976
rect 9088 7964 9094 8016
rect 9766 7964 9772 8016
rect 9824 8004 9830 8016
rect 10134 8004 10140 8016
rect 9824 7976 10140 8004
rect 9824 7964 9830 7976
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 10505 8007 10563 8013
rect 10505 7973 10517 8007
rect 10551 8004 10563 8007
rect 10870 8004 10876 8016
rect 10551 7976 10876 8004
rect 10551 7973 10563 7976
rect 10505 7967 10563 7973
rect 10870 7964 10876 7976
rect 10928 7964 10934 8016
rect 8662 7896 8668 7948
rect 8720 7936 8726 7948
rect 9398 7936 9404 7948
rect 8720 7908 9404 7936
rect 8720 7896 8726 7908
rect 9398 7896 9404 7908
rect 9456 7936 9462 7948
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 9456 7908 9505 7936
rect 9456 7896 9462 7908
rect 9493 7905 9505 7908
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 9861 7939 9919 7945
rect 9861 7936 9873 7939
rect 9732 7908 9873 7936
rect 9732 7896 9738 7908
rect 9861 7905 9873 7908
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 10042 7896 10048 7948
rect 10100 7896 10106 7948
rect 10594 7896 10600 7948
rect 10652 7936 10658 7948
rect 12811 7945 12839 8044
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 13998 8072 14004 8084
rect 13372 8044 14004 8072
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 10652 7908 11161 7936
rect 10652 7896 10658 7908
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 11149 7899 11207 7905
rect 12805 7939 12863 7945
rect 12805 7905 12817 7939
rect 12851 7905 12863 7939
rect 12805 7899 12863 7905
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 8036 7840 8309 7868
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8384 7871 8447 7877
rect 8384 7840 8401 7871
rect 8297 7831 8355 7837
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 8496 7840 8984 7868
rect 2498 7760 2504 7812
rect 2556 7800 2562 7812
rect 3237 7803 3295 7809
rect 3237 7800 3249 7803
rect 2556 7772 3249 7800
rect 2556 7760 2562 7772
rect 3237 7769 3249 7772
rect 3283 7800 3295 7803
rect 3283 7772 4660 7800
rect 3283 7769 3295 7772
rect 3237 7763 3295 7769
rect 1578 7732 1584 7744
rect 1539 7704 1584 7732
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 2038 7732 2044 7744
rect 1999 7704 2044 7732
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 3329 7735 3387 7741
rect 3329 7701 3341 7735
rect 3375 7732 3387 7735
rect 3694 7732 3700 7744
rect 3375 7704 3700 7732
rect 3375 7701 3387 7704
rect 3329 7695 3387 7701
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 3789 7735 3847 7741
rect 3789 7701 3801 7735
rect 3835 7732 3847 7735
rect 3878 7732 3884 7744
rect 3835 7704 3884 7732
rect 3835 7701 3847 7704
rect 3789 7695 3847 7701
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 4632 7732 4660 7772
rect 4706 7760 4712 7812
rect 4764 7800 4770 7812
rect 6457 7803 6515 7809
rect 6457 7800 6469 7803
rect 4764 7772 6469 7800
rect 4764 7760 4770 7772
rect 6457 7769 6469 7772
rect 6503 7800 6515 7803
rect 7576 7800 7604 7828
rect 6503 7772 7604 7800
rect 6503 7769 6515 7772
rect 6457 7763 6515 7769
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 8496 7800 8524 7840
rect 8846 7800 8852 7812
rect 8168 7772 8524 7800
rect 8588 7772 8852 7800
rect 8168 7760 8174 7772
rect 5074 7732 5080 7744
rect 4632 7704 5080 7732
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 5626 7732 5632 7744
rect 5587 7704 5632 7732
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 5721 7735 5779 7741
rect 5721 7701 5733 7735
rect 5767 7732 5779 7735
rect 5810 7732 5816 7744
rect 5767 7704 5816 7732
rect 5767 7701 5779 7704
rect 5721 7695 5779 7701
rect 5810 7692 5816 7704
rect 5868 7692 5874 7744
rect 6549 7735 6607 7741
rect 6549 7701 6561 7735
rect 6595 7732 6607 7735
rect 7006 7732 7012 7744
rect 6595 7704 7012 7732
rect 6595 7701 6607 7704
rect 6549 7695 6607 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 7745 7735 7803 7741
rect 7745 7701 7757 7735
rect 7791 7732 7803 7735
rect 7834 7732 7840 7744
rect 7791 7704 7840 7732
rect 7791 7701 7803 7704
rect 7745 7695 7803 7701
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 8588 7732 8616 7772
rect 8846 7760 8852 7772
rect 8904 7760 8910 7812
rect 8956 7800 8984 7840
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 9180 7840 9321 7868
rect 9180 7828 9186 7840
rect 9309 7837 9321 7840
rect 9355 7868 9367 7871
rect 10060 7868 10088 7896
rect 9355 7840 10088 7868
rect 10137 7871 10195 7877
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 10137 7837 10149 7871
rect 10183 7868 10195 7871
rect 10686 7868 10692 7880
rect 10183 7840 10692 7868
rect 10183 7837 10195 7840
rect 10137 7831 10195 7837
rect 10686 7828 10692 7840
rect 10744 7828 10750 7880
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7868 11115 7871
rect 11790 7868 11796 7880
rect 11103 7840 11796 7868
rect 11103 7837 11115 7840
rect 11057 7831 11115 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7868 13323 7871
rect 13372 7868 13400 8044
rect 13998 8032 14004 8044
rect 14056 8072 14062 8084
rect 15194 8072 15200 8084
rect 14056 8044 15200 8072
rect 14056 8032 14062 8044
rect 15194 8032 15200 8044
rect 15252 8032 15258 8084
rect 16206 8032 16212 8084
rect 16264 8072 16270 8084
rect 16301 8075 16359 8081
rect 16301 8072 16313 8075
rect 16264 8044 16313 8072
rect 16264 8032 16270 8044
rect 16301 8041 16313 8044
rect 16347 8041 16359 8075
rect 16301 8035 16359 8041
rect 16577 8075 16635 8081
rect 16577 8041 16589 8075
rect 16623 8072 16635 8075
rect 17402 8072 17408 8084
rect 16623 8044 17408 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 18874 8032 18880 8084
rect 18932 8072 18938 8084
rect 19245 8075 19303 8081
rect 19245 8072 19257 8075
rect 18932 8044 19257 8072
rect 18932 8032 18938 8044
rect 19245 8041 19257 8044
rect 19291 8041 19303 8075
rect 20162 8072 20168 8084
rect 20123 8044 20168 8072
rect 19245 8035 19303 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 21082 8032 21088 8084
rect 21140 8072 21146 8084
rect 21361 8075 21419 8081
rect 21361 8072 21373 8075
rect 21140 8044 21373 8072
rect 21140 8032 21146 8044
rect 21361 8041 21373 8044
rect 21407 8041 21419 8075
rect 21361 8035 21419 8041
rect 21450 8032 21456 8084
rect 21508 8072 21514 8084
rect 21508 8044 21553 8072
rect 21508 8032 21514 8044
rect 13909 8007 13967 8013
rect 13909 7973 13921 8007
rect 13955 8004 13967 8007
rect 15102 8004 15108 8016
rect 13955 7976 15108 8004
rect 13955 7973 13967 7976
rect 13909 7967 13967 7973
rect 15102 7964 15108 7976
rect 15160 7964 15166 8016
rect 16761 8007 16819 8013
rect 16761 7973 16773 8007
rect 16807 8004 16819 8007
rect 17586 8004 17592 8016
rect 16807 7976 17448 8004
rect 17547 7976 17592 8004
rect 16807 7973 16819 7976
rect 16761 7967 16819 7973
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7905 13507 7939
rect 14734 7936 14740 7948
rect 14695 7908 14740 7936
rect 13449 7899 13507 7905
rect 13311 7840 13400 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 9214 7800 9220 7812
rect 8956 7772 9220 7800
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 10045 7803 10103 7809
rect 10045 7769 10057 7803
rect 10091 7800 10103 7803
rect 10091 7772 10640 7800
rect 10091 7769 10103 7772
rect 10045 7763 10103 7769
rect 8076 7704 8616 7732
rect 8076 7692 8082 7704
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8720 7704 8953 7732
rect 8720 7692 8726 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 8941 7695 8999 7701
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 10226 7732 10232 7744
rect 9447 7704 10232 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 10612 7741 10640 7772
rect 12342 7760 12348 7812
rect 12400 7800 12406 7812
rect 12560 7803 12618 7809
rect 12560 7800 12572 7803
rect 12400 7772 12572 7800
rect 12400 7760 12406 7772
rect 12560 7769 12572 7772
rect 12606 7800 12618 7803
rect 13464 7800 13492 7899
rect 14734 7896 14740 7908
rect 14792 7936 14798 7948
rect 15565 7939 15623 7945
rect 15565 7936 15577 7939
rect 14792 7908 15577 7936
rect 14792 7896 14798 7908
rect 15565 7905 15577 7908
rect 15611 7905 15623 7939
rect 15565 7899 15623 7905
rect 17037 7939 17095 7945
rect 17037 7905 17049 7939
rect 17083 7936 17095 7939
rect 17126 7936 17132 7948
rect 17083 7908 17132 7936
rect 17083 7905 17095 7908
rect 17037 7899 17095 7905
rect 17126 7896 17132 7908
rect 17184 7896 17190 7948
rect 13722 7868 13728 7880
rect 13683 7840 13728 7868
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 15010 7868 15016 7880
rect 14599 7840 15016 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15470 7868 15476 7880
rect 15431 7840 15476 7868
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7868 17279 7871
rect 17310 7868 17316 7880
rect 17267 7840 17316 7868
rect 17267 7837 17279 7840
rect 17221 7831 17279 7837
rect 17310 7828 17316 7840
rect 17368 7828 17374 7880
rect 17420 7868 17448 7976
rect 17586 7964 17592 7976
rect 17644 7964 17650 8016
rect 18966 7964 18972 8016
rect 19024 8004 19030 8016
rect 19061 8007 19119 8013
rect 19061 8004 19073 8007
rect 19024 7976 19073 8004
rect 19024 7964 19030 7976
rect 19061 7973 19073 7976
rect 19107 8004 19119 8007
rect 20254 8004 20260 8016
rect 19107 7976 19840 8004
rect 20215 7976 20260 8004
rect 19107 7973 19119 7976
rect 19061 7967 19119 7973
rect 17494 7896 17500 7948
rect 17552 7936 17558 7948
rect 19812 7945 19840 7976
rect 20254 7964 20260 7976
rect 20312 7964 20318 8016
rect 20438 7964 20444 8016
rect 20496 7964 20502 8016
rect 17681 7939 17739 7945
rect 17681 7936 17693 7939
rect 17552 7908 17693 7936
rect 17552 7896 17558 7908
rect 17681 7905 17693 7908
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7905 19855 7939
rect 19797 7899 19855 7905
rect 20162 7896 20168 7948
rect 20220 7936 20226 7948
rect 20456 7936 20484 7964
rect 20714 7936 20720 7948
rect 20220 7908 20484 7936
rect 20675 7908 20720 7936
rect 20220 7896 20226 7908
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 21450 7896 21456 7948
rect 21508 7936 21514 7948
rect 21726 7936 21732 7948
rect 21508 7908 21732 7936
rect 21508 7896 21514 7908
rect 21726 7896 21732 7908
rect 21784 7896 21790 7948
rect 22462 7896 22468 7948
rect 22520 7936 22526 7948
rect 22830 7936 22836 7948
rect 22520 7908 22836 7936
rect 22520 7896 22526 7908
rect 22830 7896 22836 7908
rect 22888 7896 22894 7948
rect 17770 7868 17776 7880
rect 17420 7840 17776 7868
rect 17770 7828 17776 7840
rect 17828 7828 17834 7880
rect 20438 7868 20444 7880
rect 17880 7840 20444 7868
rect 15838 7800 15844 7812
rect 12606 7772 13492 7800
rect 15396 7772 15844 7800
rect 12606 7769 12618 7772
rect 12560 7763 12618 7769
rect 15396 7744 15424 7772
rect 15838 7760 15844 7772
rect 15896 7760 15902 7812
rect 16209 7803 16267 7809
rect 16209 7769 16221 7803
rect 16255 7800 16267 7803
rect 17880 7800 17908 7840
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 16255 7772 17908 7800
rect 17948 7803 18006 7809
rect 16255 7769 16267 7772
rect 16209 7763 16267 7769
rect 17948 7769 17960 7803
rect 17994 7800 18006 7803
rect 18506 7800 18512 7812
rect 17994 7772 18512 7800
rect 17994 7769 18006 7772
rect 17948 7763 18006 7769
rect 18506 7760 18512 7772
rect 18564 7760 18570 7812
rect 18690 7760 18696 7812
rect 18748 7800 18754 7812
rect 20901 7803 20959 7809
rect 20901 7800 20913 7803
rect 18748 7772 20913 7800
rect 18748 7760 18754 7772
rect 20901 7769 20913 7772
rect 20947 7800 20959 7803
rect 22830 7800 22836 7812
rect 20947 7772 22836 7800
rect 20947 7769 20959 7772
rect 20901 7763 20959 7769
rect 22830 7760 22836 7772
rect 22888 7760 22894 7812
rect 10597 7735 10655 7741
rect 10597 7701 10609 7735
rect 10643 7701 10655 7735
rect 10962 7732 10968 7744
rect 10923 7704 10968 7732
rect 10597 7695 10655 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11790 7732 11796 7744
rect 11112 7704 11796 7732
rect 11112 7692 11118 7704
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 12897 7735 12955 7741
rect 12897 7732 12909 7735
rect 12308 7704 12909 7732
rect 12308 7692 12314 7704
rect 12897 7701 12909 7704
rect 12943 7701 12955 7735
rect 12897 7695 12955 7701
rect 13078 7692 13084 7744
rect 13136 7732 13142 7744
rect 13357 7735 13415 7741
rect 13357 7732 13369 7735
rect 13136 7704 13369 7732
rect 13136 7692 13142 7704
rect 13357 7701 13369 7704
rect 13403 7701 13415 7735
rect 13357 7695 13415 7701
rect 14185 7735 14243 7741
rect 14185 7701 14197 7735
rect 14231 7732 14243 7735
rect 14458 7732 14464 7744
rect 14231 7704 14464 7732
rect 14231 7701 14243 7704
rect 14185 7695 14243 7701
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 14608 7704 14657 7732
rect 14608 7692 14614 7704
rect 14645 7701 14657 7704
rect 14691 7701 14703 7735
rect 15010 7732 15016 7744
rect 14971 7704 15016 7732
rect 14645 7695 14703 7701
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 15378 7732 15384 7744
rect 15339 7704 15384 7732
rect 15378 7692 15384 7704
rect 15436 7692 15442 7744
rect 17129 7735 17187 7741
rect 17129 7701 17141 7735
rect 17175 7732 17187 7735
rect 18782 7732 18788 7744
rect 17175 7704 18788 7732
rect 17175 7701 17187 7704
rect 17129 7695 17187 7701
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19613 7735 19671 7741
rect 19613 7732 19625 7735
rect 19392 7704 19625 7732
rect 19392 7692 19398 7704
rect 19613 7701 19625 7704
rect 19659 7701 19671 7735
rect 19613 7695 19671 7701
rect 19702 7692 19708 7744
rect 19760 7732 19766 7744
rect 20993 7735 21051 7741
rect 19760 7704 19805 7732
rect 19760 7692 19766 7704
rect 20993 7701 21005 7735
rect 21039 7732 21051 7735
rect 21266 7732 21272 7744
rect 21039 7704 21272 7732
rect 21039 7701 21051 7704
rect 20993 7695 21051 7701
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 1949 7531 2007 7537
rect 1949 7528 1961 7531
rect 1820 7500 1961 7528
rect 1820 7488 1826 7500
rect 1949 7497 1961 7500
rect 1995 7497 2007 7531
rect 1949 7491 2007 7497
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 2498 7528 2504 7540
rect 2455 7500 2504 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 4246 7528 4252 7540
rect 2832 7500 2877 7528
rect 4207 7500 4252 7528
rect 2832 7488 2838 7500
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4706 7528 4712 7540
rect 4667 7500 4712 7528
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 6181 7531 6239 7537
rect 6181 7497 6193 7531
rect 6227 7528 6239 7531
rect 6730 7528 6736 7540
rect 6227 7500 6736 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7101 7531 7159 7537
rect 7101 7497 7113 7531
rect 7147 7497 7159 7531
rect 7558 7528 7564 7540
rect 7519 7500 7564 7528
rect 7101 7491 7159 7497
rect 934 7420 940 7472
rect 992 7460 998 7472
rect 1489 7463 1547 7469
rect 1489 7460 1501 7463
rect 992 7432 1501 7460
rect 992 7420 998 7432
rect 1489 7429 1501 7432
rect 1535 7429 1547 7463
rect 1489 7423 1547 7429
rect 2317 7463 2375 7469
rect 2317 7429 2329 7463
rect 2363 7460 2375 7463
rect 2363 7432 2774 7460
rect 2363 7429 2375 7432
rect 2317 7423 2375 7429
rect 1854 7284 1860 7336
rect 1912 7324 1918 7336
rect 2406 7324 2412 7336
rect 1912 7296 2412 7324
rect 1912 7284 1918 7296
rect 2406 7284 2412 7296
rect 2464 7324 2470 7336
rect 2501 7327 2559 7333
rect 2501 7324 2513 7327
rect 2464 7296 2513 7324
rect 2464 7284 2470 7296
rect 2501 7293 2513 7296
rect 2547 7293 2559 7327
rect 2501 7287 2559 7293
rect 1670 7256 1676 7268
rect 1631 7228 1676 7256
rect 1670 7216 1676 7228
rect 1728 7216 1734 7268
rect 2746 7256 2774 7432
rect 2866 7420 2872 7472
rect 2924 7460 2930 7472
rect 7116 7460 7144 7491
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 8018 7528 8024 7540
rect 7944 7500 8024 7528
rect 7944 7460 7972 7500
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 9030 7488 9036 7540
rect 9088 7528 9094 7540
rect 9953 7531 10011 7537
rect 9953 7528 9965 7531
rect 9088 7500 9965 7528
rect 9088 7488 9094 7500
rect 9953 7497 9965 7500
rect 9999 7497 10011 7531
rect 9953 7491 10011 7497
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 10284 7500 10333 7528
rect 10284 7488 10290 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 11333 7531 11391 7537
rect 11333 7528 11345 7531
rect 10321 7491 10379 7497
rect 11256 7500 11345 7528
rect 8110 7460 8116 7472
rect 2924 7432 6960 7460
rect 7116 7432 7972 7460
rect 8036 7432 8116 7460
rect 2924 7420 2930 7432
rect 2958 7352 2964 7404
rect 3016 7392 3022 7404
rect 3602 7392 3608 7404
rect 3016 7364 3608 7392
rect 3016 7352 3022 7364
rect 3602 7352 3608 7364
rect 3660 7392 3666 7404
rect 3890 7395 3948 7401
rect 3890 7392 3902 7395
rect 3660 7364 3902 7392
rect 3660 7352 3666 7364
rect 3890 7361 3902 7364
rect 3936 7361 3948 7395
rect 3890 7355 3948 7361
rect 4062 7352 4068 7404
rect 4120 7392 4126 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 4120 7364 4169 7392
rect 4120 7352 4126 7364
rect 4157 7361 4169 7364
rect 4203 7392 4215 7395
rect 4246 7392 4252 7404
rect 4203 7364 4252 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 4430 7392 4436 7404
rect 4391 7364 4436 7392
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 4706 7392 4712 7404
rect 4571 7364 4712 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 4890 7352 4896 7404
rect 4948 7392 4954 7404
rect 5057 7395 5115 7401
rect 5057 7392 5069 7395
rect 4948 7364 5069 7392
rect 4948 7352 4954 7364
rect 5057 7361 5069 7364
rect 5103 7361 5115 7395
rect 5057 7355 5115 7361
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 6932 7401 6960 7432
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 5500 7364 6377 7392
rect 5500 7352 5506 7364
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6641 7395 6699 7401
rect 6641 7392 6653 7395
rect 6365 7355 6423 7361
rect 6472 7364 6653 7392
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 2746 7228 2912 7256
rect 1762 7188 1768 7200
rect 1723 7160 1768 7188
rect 1762 7148 1768 7160
rect 1820 7188 1826 7200
rect 2774 7188 2780 7200
rect 1820 7160 2780 7188
rect 1820 7148 1826 7160
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 2884 7188 2912 7228
rect 4430 7216 4436 7268
rect 4488 7256 4494 7268
rect 4816 7256 4844 7287
rect 6472 7256 6500 7364
rect 6641 7361 6653 7364
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 6917 7395 6975 7401
rect 6917 7361 6929 7395
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 7374 7352 7380 7404
rect 7432 7392 7438 7404
rect 8036 7401 8064 7432
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 8277 7463 8335 7469
rect 8277 7429 8289 7463
rect 8323 7429 8335 7463
rect 8277 7423 8335 7429
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 7432 7364 7665 7392
rect 7432 7352 7438 7364
rect 7653 7361 7665 7364
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7361 8079 7395
rect 8303 7392 8331 7423
rect 8386 7420 8392 7472
rect 8444 7460 8450 7472
rect 8662 7460 8668 7472
rect 8444 7432 8668 7460
rect 8444 7420 8450 7432
rect 8662 7420 8668 7432
rect 8720 7420 8726 7472
rect 8846 7420 8852 7472
rect 8904 7460 8910 7472
rect 10042 7460 10048 7472
rect 8904 7432 10048 7460
rect 8904 7420 8910 7432
rect 10042 7420 10048 7432
rect 10100 7460 10106 7472
rect 10594 7460 10600 7472
rect 10100 7432 10600 7460
rect 10100 7420 10106 7432
rect 10594 7420 10600 7432
rect 10652 7420 10658 7472
rect 10778 7460 10784 7472
rect 10704 7432 10784 7460
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 8021 7355 8079 7361
rect 8128 7364 8331 7392
rect 9324 7364 9873 7392
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 7834 7324 7840 7336
rect 6604 7296 7512 7324
rect 7795 7296 7840 7324
rect 6604 7284 6610 7296
rect 7374 7256 7380 7268
rect 4488 7228 4844 7256
rect 4488 7216 4494 7228
rect 4338 7188 4344 7200
rect 2884 7160 4344 7188
rect 4338 7148 4344 7160
rect 4396 7188 4402 7200
rect 4706 7188 4712 7200
rect 4396 7160 4712 7188
rect 4396 7148 4402 7160
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 4816 7188 4844 7228
rect 5736 7228 6500 7256
rect 6748 7228 7380 7256
rect 5166 7188 5172 7200
rect 4816 7160 5172 7188
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 5736 7188 5764 7228
rect 5592 7160 5764 7188
rect 5592 7148 5598 7160
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 5868 7160 6561 7188
rect 5868 7148 5874 7160
rect 6549 7157 6561 7160
rect 6595 7188 6607 7191
rect 6748 7188 6776 7228
rect 7374 7216 7380 7228
rect 7432 7216 7438 7268
rect 6595 7160 6776 7188
rect 6825 7191 6883 7197
rect 6595 7157 6607 7160
rect 6549 7151 6607 7157
rect 6825 7157 6837 7191
rect 6871 7188 6883 7191
rect 6914 7188 6920 7200
rect 6871 7160 6920 7188
rect 6871 7157 6883 7160
rect 6825 7151 6883 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7484 7188 7512 7296
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 8128 7324 8156 7364
rect 9324 7324 9352 7364
rect 9861 7361 9873 7364
rect 9907 7392 9919 7395
rect 10134 7392 10140 7404
rect 9907 7364 10140 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 8036 7296 8156 7324
rect 9039 7296 9352 7324
rect 8036 7268 8064 7296
rect 8018 7216 8024 7268
rect 8076 7216 8082 7268
rect 9039 7188 9067 7296
rect 9398 7284 9404 7336
rect 9456 7324 9462 7336
rect 10704 7333 10732 7432
rect 10778 7420 10784 7432
rect 10836 7420 10842 7472
rect 10873 7463 10931 7469
rect 10873 7429 10885 7463
rect 10919 7429 10931 7463
rect 10873 7423 10931 7429
rect 10965 7463 11023 7469
rect 10965 7429 10977 7463
rect 11011 7460 11023 7463
rect 11146 7460 11152 7472
rect 11011 7432 11152 7460
rect 11011 7429 11023 7432
rect 10965 7423 11023 7429
rect 10888 7392 10916 7423
rect 11146 7420 11152 7432
rect 11204 7420 11210 7472
rect 10888 7364 11008 7392
rect 10045 7327 10103 7333
rect 10045 7324 10057 7327
rect 9456 7296 10057 7324
rect 9456 7284 9462 7296
rect 10045 7293 10057 7296
rect 10091 7293 10103 7327
rect 10045 7287 10103 7293
rect 10689 7327 10747 7333
rect 10689 7293 10701 7327
rect 10735 7293 10747 7327
rect 10980 7324 11008 7364
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 11256 7392 11284 7500
rect 11333 7497 11345 7500
rect 11379 7497 11391 7531
rect 11333 7491 11391 7497
rect 11790 7488 11796 7540
rect 11848 7528 11854 7540
rect 11885 7531 11943 7537
rect 11885 7528 11897 7531
rect 11848 7500 11897 7528
rect 11848 7488 11854 7500
rect 11885 7497 11897 7500
rect 11931 7497 11943 7531
rect 12158 7528 12164 7540
rect 12119 7500 12164 7528
rect 11885 7491 11943 7497
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 12618 7528 12624 7540
rect 12579 7500 12624 7528
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 13998 7528 14004 7540
rect 13004 7500 14004 7528
rect 11422 7420 11428 7472
rect 11480 7460 11486 7472
rect 11609 7463 11667 7469
rect 11609 7460 11621 7463
rect 11480 7432 11621 7460
rect 11480 7420 11486 7432
rect 11609 7429 11621 7432
rect 11655 7460 11667 7463
rect 12250 7460 12256 7472
rect 11655 7432 12256 7460
rect 11655 7429 11667 7432
rect 11609 7423 11667 7429
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 11112 7364 11284 7392
rect 11112 7352 11118 7364
rect 11974 7352 11980 7404
rect 12032 7392 12038 7404
rect 12529 7395 12587 7401
rect 12529 7392 12541 7395
rect 12032 7364 12541 7392
rect 12032 7352 12038 7364
rect 12529 7361 12541 7364
rect 12575 7392 12587 7395
rect 12802 7392 12808 7404
rect 12575 7364 12808 7392
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 11790 7324 11796 7336
rect 10980 7296 11796 7324
rect 10689 7287 10747 7293
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 9122 7216 9128 7268
rect 9180 7256 9186 7268
rect 9493 7259 9551 7265
rect 9493 7256 9505 7259
rect 9180 7228 9505 7256
rect 9180 7216 9186 7228
rect 9493 7225 9505 7228
rect 9539 7225 9551 7259
rect 9493 7219 9551 7225
rect 9858 7216 9864 7268
rect 9916 7256 9922 7268
rect 11146 7256 11152 7268
rect 9916 7228 11152 7256
rect 9916 7216 9922 7228
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 12342 7216 12348 7268
rect 12400 7256 12406 7268
rect 12728 7256 12756 7287
rect 12894 7284 12900 7336
rect 12952 7284 12958 7336
rect 13004 7333 13032 7500
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 15010 7488 15016 7540
rect 15068 7528 15074 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 15068 7500 15301 7528
rect 15068 7488 15074 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 17678 7528 17684 7540
rect 16347 7500 17684 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 19334 7528 19340 7540
rect 19295 7500 19340 7528
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 19429 7531 19487 7537
rect 19429 7497 19441 7531
rect 19475 7528 19487 7531
rect 19702 7528 19708 7540
rect 19475 7500 19708 7528
rect 19475 7497 19487 7500
rect 19429 7491 19487 7497
rect 19702 7488 19708 7500
rect 19760 7488 19766 7540
rect 20346 7528 20352 7540
rect 20307 7500 20352 7528
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 20441 7531 20499 7537
rect 20441 7497 20453 7531
rect 20487 7528 20499 7531
rect 20806 7528 20812 7540
rect 20487 7500 20812 7528
rect 20487 7497 20499 7500
rect 20441 7491 20499 7497
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 14734 7460 14740 7472
rect 14200 7432 14740 7460
rect 13808 7395 13866 7401
rect 13808 7361 13820 7395
rect 13854 7392 13866 7395
rect 14200 7392 14228 7432
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 16117 7463 16175 7469
rect 16117 7429 16129 7463
rect 16163 7460 16175 7463
rect 16390 7460 16396 7472
rect 16163 7432 16396 7460
rect 16163 7429 16175 7432
rect 16117 7423 16175 7429
rect 16390 7420 16396 7432
rect 16448 7420 16454 7472
rect 17037 7463 17095 7469
rect 17037 7429 17049 7463
rect 17083 7460 17095 7463
rect 19518 7460 19524 7472
rect 17083 7432 19524 7460
rect 17083 7429 17095 7432
rect 17037 7423 17095 7429
rect 19518 7420 19524 7432
rect 19576 7420 19582 7472
rect 20622 7420 20628 7472
rect 20680 7460 20686 7472
rect 20901 7463 20959 7469
rect 20901 7460 20913 7463
rect 20680 7432 20913 7460
rect 20680 7420 20686 7432
rect 20901 7429 20913 7432
rect 20947 7429 20959 7463
rect 20901 7423 20959 7429
rect 20990 7420 20996 7472
rect 21048 7420 21054 7472
rect 13854 7364 14228 7392
rect 13854 7361 13866 7364
rect 13808 7355 13866 7361
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 15010 7392 15016 7404
rect 14332 7364 15016 7392
rect 14332 7352 14338 7364
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 15378 7392 15384 7404
rect 15339 7364 15384 7392
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 17218 7392 17224 7404
rect 17175 7364 17224 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 17402 7401 17408 7404
rect 17396 7392 17408 7401
rect 17363 7364 17408 7392
rect 17396 7355 17408 7364
rect 17402 7352 17408 7355
rect 17460 7352 17466 7404
rect 18966 7392 18972 7404
rect 18927 7364 18972 7392
rect 18966 7352 18972 7364
rect 19024 7352 19030 7404
rect 19797 7395 19855 7401
rect 19797 7361 19809 7395
rect 19843 7392 19855 7395
rect 20346 7392 20352 7404
rect 19843 7364 20352 7392
rect 19843 7361 19855 7364
rect 19797 7355 19855 7361
rect 20346 7352 20352 7364
rect 20404 7352 20410 7404
rect 20806 7392 20812 7404
rect 20767 7364 20812 7392
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 12989 7327 13047 7333
rect 12989 7293 13001 7327
rect 13035 7293 13047 7327
rect 12989 7287 13047 7293
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 13541 7327 13599 7333
rect 13541 7324 13553 7327
rect 13504 7296 13553 7324
rect 13504 7284 13510 7296
rect 13541 7293 13553 7296
rect 13587 7293 13599 7327
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 13541 7287 13599 7293
rect 14936 7296 15117 7324
rect 12400 7228 12756 7256
rect 12912 7256 12940 7284
rect 12912 7228 13584 7256
rect 12400 7216 12406 7228
rect 9398 7188 9404 7200
rect 7484 7160 9067 7188
rect 9359 7160 9404 7188
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 11422 7188 11428 7200
rect 10192 7160 11428 7188
rect 10192 7148 10198 7160
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 11698 7188 11704 7200
rect 11659 7160 11704 7188
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 13078 7148 13084 7200
rect 13136 7188 13142 7200
rect 13173 7191 13231 7197
rect 13173 7188 13185 7191
rect 13136 7160 13185 7188
rect 13136 7148 13142 7160
rect 13173 7157 13185 7160
rect 13219 7157 13231 7191
rect 13354 7188 13360 7200
rect 13315 7160 13360 7188
rect 13173 7151 13231 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 13556 7188 13584 7228
rect 13722 7188 13728 7200
rect 13556 7160 13728 7188
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 14274 7148 14280 7200
rect 14332 7188 14338 7200
rect 14936 7197 14964 7296
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 15286 7284 15292 7336
rect 15344 7324 15350 7336
rect 16022 7324 16028 7336
rect 15344 7296 16028 7324
rect 15344 7284 15350 7296
rect 16022 7284 16028 7296
rect 16080 7324 16086 7336
rect 16393 7327 16451 7333
rect 16393 7324 16405 7327
rect 16080 7296 16405 7324
rect 16080 7284 16086 7296
rect 16393 7293 16405 7296
rect 16439 7293 16451 7327
rect 16393 7287 16451 7293
rect 16666 7284 16672 7336
rect 16724 7324 16730 7336
rect 17034 7324 17040 7336
rect 16724 7296 17040 7324
rect 16724 7284 16730 7296
rect 17034 7284 17040 7296
rect 17092 7284 17098 7336
rect 18693 7327 18751 7333
rect 18693 7293 18705 7327
rect 18739 7293 18751 7327
rect 18874 7324 18880 7336
rect 18835 7296 18880 7324
rect 18693 7287 18751 7293
rect 15933 7259 15991 7265
rect 15933 7225 15945 7259
rect 15979 7256 15991 7259
rect 16298 7256 16304 7268
rect 15979 7228 16304 7256
rect 15979 7225 15991 7228
rect 15933 7219 15991 7225
rect 16298 7216 16304 7228
rect 16356 7216 16362 7268
rect 18506 7256 18512 7268
rect 18419 7228 18512 7256
rect 18506 7216 18512 7228
rect 18564 7256 18570 7268
rect 18708 7256 18736 7287
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 19886 7324 19892 7336
rect 19847 7296 19892 7324
rect 19886 7284 19892 7296
rect 19944 7284 19950 7336
rect 21008 7333 21036 7420
rect 21453 7395 21511 7401
rect 21453 7392 21465 7395
rect 21376 7364 21465 7392
rect 19981 7327 20039 7333
rect 19981 7293 19993 7327
rect 20027 7293 20039 7327
rect 19981 7287 20039 7293
rect 20993 7327 21051 7333
rect 20993 7293 21005 7327
rect 21039 7293 21051 7327
rect 20993 7287 21051 7293
rect 19996 7256 20024 7287
rect 18564 7228 20024 7256
rect 18564 7216 18570 7228
rect 20254 7216 20260 7268
rect 20312 7256 20318 7268
rect 21269 7259 21327 7265
rect 21269 7256 21281 7259
rect 20312 7228 21281 7256
rect 20312 7216 20318 7228
rect 21269 7225 21281 7228
rect 21315 7225 21327 7259
rect 21269 7219 21327 7225
rect 14921 7191 14979 7197
rect 14921 7188 14933 7191
rect 14332 7160 14933 7188
rect 14332 7148 14338 7160
rect 14921 7157 14933 7160
rect 14967 7157 14979 7191
rect 15746 7188 15752 7200
rect 15707 7160 15752 7188
rect 14921 7151 14979 7157
rect 15746 7148 15752 7160
rect 15804 7148 15810 7200
rect 16482 7148 16488 7200
rect 16540 7188 16546 7200
rect 16669 7191 16727 7197
rect 16669 7188 16681 7191
rect 16540 7160 16681 7188
rect 16540 7148 16546 7160
rect 16669 7157 16681 7160
rect 16715 7157 16727 7191
rect 16669 7151 16727 7157
rect 17126 7148 17132 7200
rect 17184 7188 17190 7200
rect 21082 7188 21088 7200
rect 17184 7160 21088 7188
rect 17184 7148 17190 7160
rect 21082 7148 21088 7160
rect 21140 7188 21146 7200
rect 21376 7188 21404 7364
rect 21453 7361 21465 7364
rect 21499 7361 21511 7395
rect 21453 7355 21511 7361
rect 21140 7160 21404 7188
rect 21140 7148 21146 7160
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 2038 6944 2044 6996
rect 2096 6984 2102 6996
rect 2409 6987 2467 6993
rect 2409 6984 2421 6987
rect 2096 6956 2421 6984
rect 2096 6944 2102 6956
rect 2409 6953 2421 6956
rect 2455 6953 2467 6987
rect 2409 6947 2467 6953
rect 3050 6944 3056 6996
rect 3108 6984 3114 6996
rect 6822 6984 6828 6996
rect 3108 6956 6828 6984
rect 3108 6944 3114 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7650 6984 7656 6996
rect 6972 6956 7656 6984
rect 6972 6944 6978 6956
rect 7650 6944 7656 6956
rect 7708 6984 7714 6996
rect 9582 6984 9588 6996
rect 7708 6956 9588 6984
rect 7708 6944 7714 6956
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 9858 6984 9864 6996
rect 9784 6956 9864 6984
rect 2774 6916 2780 6928
rect 2700 6888 2780 6916
rect 1854 6848 1860 6860
rect 1815 6820 1860 6848
rect 1854 6808 1860 6820
rect 1912 6808 1918 6860
rect 2700 6857 2728 6888
rect 2774 6876 2780 6888
rect 2832 6876 2838 6928
rect 3234 6916 3240 6928
rect 3195 6888 3240 6916
rect 3234 6876 3240 6888
rect 3292 6876 3298 6928
rect 3605 6919 3663 6925
rect 3605 6885 3617 6919
rect 3651 6916 3663 6919
rect 3970 6916 3976 6928
rect 3651 6888 3976 6916
rect 3651 6885 3663 6888
rect 3605 6879 3663 6885
rect 3970 6876 3976 6888
rect 4028 6876 4034 6928
rect 5353 6919 5411 6925
rect 5353 6885 5365 6919
rect 5399 6885 5411 6919
rect 5353 6879 5411 6885
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6817 2743 6851
rect 2685 6811 2743 6817
rect 3694 6808 3700 6860
rect 3752 6848 3758 6860
rect 4893 6851 4951 6857
rect 4893 6848 4905 6851
rect 3752 6820 4905 6848
rect 3752 6808 3758 6820
rect 4893 6817 4905 6820
rect 4939 6817 4951 6851
rect 4893 6811 4951 6817
rect 5258 6808 5264 6860
rect 5316 6848 5322 6860
rect 5368 6848 5396 6879
rect 6546 6876 6552 6928
rect 6604 6916 6610 6928
rect 7190 6916 7196 6928
rect 6604 6888 7196 6916
rect 6604 6876 6610 6888
rect 7190 6876 7196 6888
rect 7248 6876 7254 6928
rect 9784 6916 9812 6956
rect 9858 6944 9864 6956
rect 9916 6944 9922 6996
rect 9968 6956 10916 6984
rect 9968 6916 9996 6956
rect 8588 6888 9812 6916
rect 9876 6888 9996 6916
rect 5316 6820 5396 6848
rect 5316 6808 5322 6820
rect 5810 6808 5816 6860
rect 5868 6848 5874 6860
rect 6089 6851 6147 6857
rect 6089 6848 6101 6851
rect 5868 6820 6101 6848
rect 5868 6808 5874 6820
rect 6089 6817 6101 6820
rect 6135 6817 6147 6851
rect 6917 6851 6975 6857
rect 6917 6848 6929 6851
rect 6089 6811 6147 6817
rect 6196 6820 6929 6848
rect 106 6740 112 6792
rect 164 6780 170 6792
rect 934 6780 940 6792
rect 164 6752 940 6780
rect 164 6740 170 6752
rect 934 6740 940 6752
rect 992 6740 998 6792
rect 1210 6740 1216 6792
rect 1268 6780 1274 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 1268 6752 1409 6780
rect 1268 6740 1274 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 2774 6780 2780 6792
rect 1995 6752 2780 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 1854 6672 1860 6724
rect 1912 6712 1918 6724
rect 1964 6712 1992 6743
rect 2774 6740 2780 6752
rect 2832 6740 2838 6792
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6780 2927 6783
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 2915 6752 3801 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 4120 6752 4165 6780
rect 4120 6740 4126 6752
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 4709 6783 4767 6789
rect 4709 6780 4721 6783
rect 4396 6752 4721 6780
rect 4396 6740 4402 6752
rect 4709 6749 4721 6752
rect 4755 6749 4767 6783
rect 4709 6743 4767 6749
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 1912 6684 1992 6712
rect 1912 6672 1918 6684
rect 2038 6672 2044 6724
rect 2096 6712 2102 6724
rect 3421 6715 3479 6721
rect 2096 6684 2141 6712
rect 2096 6672 2102 6684
rect 3421 6681 3433 6715
rect 3467 6712 3479 6715
rect 3510 6712 3516 6724
rect 3467 6684 3516 6712
rect 3467 6681 3479 6684
rect 3421 6675 3479 6681
rect 3510 6672 3516 6684
rect 3568 6672 3574 6724
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 3234 6644 3240 6656
rect 2832 6616 3240 6644
rect 2832 6604 2838 6616
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3326 6604 3332 6656
rect 3384 6644 3390 6656
rect 4080 6644 4108 6740
rect 5184 6712 5212 6743
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 6196 6780 6224 6820
rect 6917 6817 6929 6820
rect 6963 6817 6975 6851
rect 8588 6848 8616 6888
rect 6917 6811 6975 6817
rect 8496 6820 8616 6848
rect 5776 6752 6224 6780
rect 5776 6740 5782 6752
rect 7190 6740 7196 6792
rect 7248 6740 7254 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 8496 6780 8524 6820
rect 9030 6808 9036 6860
rect 9088 6848 9094 6860
rect 9876 6848 9904 6888
rect 10888 6857 10916 6956
rect 11146 6944 11152 6996
rect 11204 6944 11210 6996
rect 11790 6984 11796 6996
rect 11751 6956 11796 6984
rect 11790 6944 11796 6956
rect 11848 6944 11854 6996
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 12308 6956 15139 6984
rect 12308 6944 12314 6956
rect 11164 6916 11192 6944
rect 12526 6916 12532 6928
rect 11164 6888 12532 6916
rect 12526 6876 12532 6888
rect 12584 6876 12590 6928
rect 14734 6916 14740 6928
rect 12728 6888 14740 6916
rect 9088 6820 9904 6848
rect 10873 6851 10931 6857
rect 9088 6808 9094 6820
rect 10873 6817 10885 6851
rect 10919 6817 10931 6851
rect 10873 6811 10931 6817
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 11204 6820 11529 6848
rect 11204 6808 11210 6820
rect 11517 6817 11529 6820
rect 11563 6817 11575 6851
rect 11517 6811 11575 6817
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 12342 6848 12348 6860
rect 11940 6820 12348 6848
rect 11940 6808 11946 6820
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 12728 6857 12756 6888
rect 14734 6876 14740 6888
rect 14792 6916 14798 6928
rect 15111 6916 15139 6956
rect 15378 6944 15384 6996
rect 15436 6984 15442 6996
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 15436 6956 15669 6984
rect 15436 6944 15442 6956
rect 15657 6953 15669 6956
rect 15703 6953 15715 6987
rect 15657 6947 15715 6953
rect 16390 6944 16396 6996
rect 16448 6984 16454 6996
rect 17126 6984 17132 6996
rect 16448 6956 17132 6984
rect 16448 6944 16454 6956
rect 17126 6944 17132 6956
rect 17184 6944 17190 6996
rect 17494 6944 17500 6996
rect 17552 6984 17558 6996
rect 17552 6956 18828 6984
rect 17552 6944 17558 6956
rect 16022 6916 16028 6928
rect 14792 6888 15056 6916
rect 15111 6888 16028 6916
rect 14792 6876 14798 6888
rect 12713 6851 12771 6857
rect 12713 6817 12725 6851
rect 12759 6817 12771 6851
rect 13541 6851 13599 6857
rect 13541 6848 13553 6851
rect 12713 6811 12771 6817
rect 12820 6820 13553 6848
rect 7524 6752 8524 6780
rect 8573 6783 8631 6789
rect 7524 6740 7530 6752
rect 8573 6749 8585 6783
rect 8619 6780 8631 6783
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8619 6752 8953 6780
rect 8619 6749 8631 6752
rect 8573 6743 8631 6749
rect 8941 6749 8953 6752
rect 8987 6780 8999 6783
rect 9214 6780 9220 6792
rect 8987 6752 9220 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 9364 6752 9413 6780
rect 9364 6740 9370 6752
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 9732 6752 10732 6780
rect 9732 6740 9738 6752
rect 4724 6684 5212 6712
rect 4724 6656 4752 6684
rect 5258 6672 5264 6724
rect 5316 6712 5322 6724
rect 5316 6684 6408 6712
rect 5316 6672 5322 6684
rect 3384 6616 4108 6644
rect 3384 6604 3390 6616
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 4249 6647 4307 6653
rect 4249 6644 4261 6647
rect 4212 6616 4261 6644
rect 4212 6604 4218 6616
rect 4249 6613 4261 6616
rect 4295 6613 4307 6647
rect 4249 6607 4307 6613
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 4396 6616 4441 6644
rect 4396 6604 4402 6616
rect 4706 6604 4712 6656
rect 4764 6604 4770 6656
rect 4801 6647 4859 6653
rect 4801 6613 4813 6647
rect 4847 6644 4859 6647
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 4847 6616 5549 6644
rect 4847 6613 4859 6616
rect 4801 6607 4859 6613
rect 5537 6613 5549 6616
rect 5583 6613 5595 6647
rect 5902 6644 5908 6656
rect 5863 6616 5908 6644
rect 5537 6607 5595 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 5994 6604 6000 6656
rect 6052 6644 6058 6656
rect 6380 6653 6408 6684
rect 6638 6672 6644 6724
rect 6696 6712 6702 6724
rect 6825 6715 6883 6721
rect 6825 6712 6837 6715
rect 6696 6684 6837 6712
rect 6696 6672 6702 6684
rect 6825 6681 6837 6684
rect 6871 6681 6883 6715
rect 7208 6712 7236 6740
rect 8018 6712 8024 6724
rect 7208 6684 8024 6712
rect 6825 6675 6883 6681
rect 8018 6672 8024 6684
rect 8076 6672 8082 6724
rect 8328 6715 8386 6721
rect 8328 6681 8340 6715
rect 8374 6712 8386 6715
rect 8374 6684 9536 6712
rect 8374 6681 8386 6684
rect 8328 6675 8386 6681
rect 9508 6656 9536 6684
rect 10410 6672 10416 6724
rect 10468 6712 10474 6724
rect 10606 6715 10664 6721
rect 10606 6712 10618 6715
rect 10468 6684 10618 6712
rect 10468 6672 10474 6684
rect 10606 6681 10618 6684
rect 10652 6681 10664 6715
rect 10704 6712 10732 6752
rect 10778 6740 10784 6792
rect 10836 6780 10842 6792
rect 12158 6780 12164 6792
rect 10836 6752 12164 6780
rect 10836 6740 10842 6752
rect 12158 6740 12164 6752
rect 12216 6740 12222 6792
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12820 6780 12848 6820
rect 13541 6817 13553 6820
rect 13587 6848 13599 6851
rect 13630 6848 13636 6860
rect 13587 6820 13636 6848
rect 13587 6817 13599 6820
rect 13541 6811 13599 6817
rect 13630 6808 13636 6820
rect 13688 6808 13694 6860
rect 14182 6848 14188 6860
rect 14143 6820 14188 6848
rect 14182 6808 14188 6820
rect 14240 6808 14246 6860
rect 15028 6857 15056 6888
rect 16022 6876 16028 6888
rect 16080 6876 16086 6928
rect 18506 6916 18512 6928
rect 18432 6888 18512 6916
rect 15013 6851 15071 6857
rect 14292 6820 14596 6848
rect 12299 6752 12848 6780
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 12894 6740 12900 6792
rect 12952 6780 12958 6792
rect 13725 6783 13783 6789
rect 13725 6780 13737 6783
rect 12952 6752 13737 6780
rect 12952 6740 12958 6752
rect 13725 6749 13737 6752
rect 13771 6780 13783 6783
rect 14292 6780 14320 6820
rect 14458 6780 14464 6792
rect 13771 6752 14320 6780
rect 14419 6752 14464 6780
rect 13771 6749 13783 6752
rect 13725 6743 13783 6749
rect 14458 6740 14464 6752
rect 14516 6740 14522 6792
rect 14568 6780 14596 6820
rect 15013 6817 15025 6851
rect 15059 6817 15071 6851
rect 15194 6848 15200 6860
rect 15155 6820 15200 6848
rect 15013 6811 15071 6817
rect 15194 6808 15200 6820
rect 15252 6808 15258 6860
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 15562 6848 15568 6860
rect 15436 6820 15568 6848
rect 15436 6808 15442 6820
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 18049 6851 18107 6857
rect 18049 6817 18061 6851
rect 18095 6848 18107 6851
rect 18138 6848 18144 6860
rect 18095 6820 18144 6848
rect 18095 6817 18107 6820
rect 18049 6811 18107 6817
rect 18138 6808 18144 6820
rect 18196 6808 18202 6860
rect 18432 6857 18460 6888
rect 18506 6876 18512 6888
rect 18564 6876 18570 6928
rect 18800 6916 18828 6956
rect 18874 6944 18880 6996
rect 18932 6984 18938 6996
rect 18969 6987 19027 6993
rect 18969 6984 18981 6987
rect 18932 6956 18981 6984
rect 18932 6944 18938 6956
rect 18969 6953 18981 6956
rect 19015 6953 19027 6987
rect 21266 6984 21272 6996
rect 18969 6947 19027 6953
rect 19260 6956 21272 6984
rect 19260 6916 19288 6956
rect 21266 6944 21272 6956
rect 21324 6944 21330 6996
rect 18800 6888 19288 6916
rect 18417 6851 18475 6857
rect 18417 6817 18429 6851
rect 18463 6817 18475 6851
rect 20990 6848 20996 6860
rect 20951 6820 20996 6848
rect 18417 6811 18475 6817
rect 20990 6808 20996 6820
rect 21048 6808 21054 6860
rect 15841 6783 15899 6789
rect 14568 6752 15608 6780
rect 15580 6724 15608 6752
rect 15841 6749 15853 6783
rect 15887 6780 15899 6783
rect 16206 6780 16212 6792
rect 15887 6752 16212 6780
rect 15887 6749 15899 6752
rect 15841 6743 15899 6749
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 17046 6783 17104 6789
rect 17046 6780 17058 6783
rect 16724 6752 17058 6780
rect 16724 6740 16730 6752
rect 17046 6749 17058 6752
rect 17092 6749 17104 6783
rect 17046 6743 17104 6749
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17313 6783 17371 6789
rect 17313 6780 17325 6783
rect 17276 6752 17325 6780
rect 17276 6740 17282 6752
rect 17313 6749 17325 6752
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 17494 6740 17500 6792
rect 17552 6780 17558 6792
rect 18509 6783 18567 6789
rect 18509 6780 18521 6783
rect 17552 6752 18521 6780
rect 17552 6740 17558 6752
rect 18509 6749 18521 6752
rect 18555 6749 18567 6783
rect 18601 6783 18659 6789
rect 18601 6780 18613 6783
rect 18509 6743 18567 6749
rect 18596 6749 18613 6780
rect 18647 6749 18659 6783
rect 18596 6743 18659 6749
rect 12989 6715 13047 6721
rect 12989 6712 13001 6715
rect 10704 6684 13001 6712
rect 10606 6675 10664 6681
rect 12989 6681 13001 6684
rect 13035 6681 13047 6715
rect 14369 6715 14427 6721
rect 14369 6712 14381 6715
rect 12989 6675 13047 6681
rect 13372 6684 14381 6712
rect 6365 6647 6423 6653
rect 6052 6616 6097 6644
rect 6052 6604 6058 6616
rect 6365 6613 6377 6647
rect 6411 6613 6423 6647
rect 6730 6644 6736 6656
rect 6691 6616 6736 6644
rect 6365 6607 6423 6613
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6644 7251 6647
rect 7374 6644 7380 6656
rect 7239 6616 7380 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 7374 6604 7380 6616
rect 7432 6644 7438 6656
rect 8202 6644 8208 6656
rect 7432 6616 8208 6644
rect 7432 6604 7438 6616
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8754 6644 8760 6656
rect 8715 6616 8760 6644
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 8938 6604 8944 6656
rect 8996 6644 9002 6656
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 8996 6616 9137 6644
rect 8996 6604 9002 6616
rect 9125 6613 9137 6616
rect 9171 6613 9183 6647
rect 9125 6607 9183 6613
rect 9217 6647 9275 6653
rect 9217 6613 9229 6647
rect 9263 6644 9275 6647
rect 9306 6644 9312 6656
rect 9263 6616 9312 6644
rect 9263 6613 9275 6616
rect 9217 6607 9275 6613
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 9490 6644 9496 6656
rect 9451 6616 9496 6644
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 10226 6604 10232 6656
rect 10284 6644 10290 6656
rect 10965 6647 11023 6653
rect 10965 6644 10977 6647
rect 10284 6616 10977 6644
rect 10284 6604 10290 6616
rect 10965 6613 10977 6616
rect 11011 6613 11023 6647
rect 10965 6607 11023 6613
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11333 6647 11391 6653
rect 11333 6644 11345 6647
rect 11296 6616 11345 6644
rect 11296 6604 11302 6616
rect 11333 6613 11345 6616
rect 11379 6613 11391 6647
rect 11333 6607 11391 6613
rect 11425 6647 11483 6653
rect 11425 6613 11437 6647
rect 11471 6644 11483 6647
rect 11698 6644 11704 6656
rect 11471 6616 11704 6644
rect 11471 6613 11483 6616
rect 11425 6607 11483 6613
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 13372 6653 13400 6684
rect 14369 6681 14381 6684
rect 14415 6681 14427 6715
rect 14369 6675 14427 6681
rect 14550 6672 14556 6724
rect 14608 6712 14614 6724
rect 15289 6715 15347 6721
rect 15289 6712 15301 6715
rect 14608 6684 15301 6712
rect 14608 6672 14614 6684
rect 15289 6681 15301 6684
rect 15335 6681 15347 6715
rect 15289 6675 15347 6681
rect 15562 6672 15568 6724
rect 15620 6672 15626 6724
rect 17678 6672 17684 6724
rect 17736 6712 17742 6724
rect 18596 6712 18624 6743
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 18840 6752 19012 6780
rect 18840 6740 18846 6752
rect 17736 6684 18624 6712
rect 17736 6672 17742 6684
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 11848 6616 12909 6644
rect 11848 6604 11854 6616
rect 12897 6613 12909 6616
rect 12943 6613 12955 6647
rect 12897 6607 12955 6613
rect 13357 6647 13415 6653
rect 13357 6613 13369 6647
rect 13403 6613 13415 6647
rect 13814 6644 13820 6656
rect 13775 6616 13820 6644
rect 13357 6607 13415 6613
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 14826 6644 14832 6656
rect 14787 6616 14832 6644
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 15930 6644 15936 6656
rect 15891 6616 15936 6644
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 17405 6647 17463 6653
rect 17405 6644 17417 6647
rect 17000 6616 17417 6644
rect 17000 6604 17006 6616
rect 17405 6613 17417 6616
rect 17451 6613 17463 6647
rect 17770 6644 17776 6656
rect 17731 6616 17776 6644
rect 17405 6607 17463 6613
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 17862 6604 17868 6656
rect 17920 6644 17926 6656
rect 18984 6644 19012 6752
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 19116 6752 19257 6780
rect 19116 6740 19122 6752
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 19512 6783 19570 6789
rect 19512 6780 19524 6783
rect 19245 6743 19303 6749
rect 19352 6752 19524 6780
rect 19150 6672 19156 6724
rect 19208 6712 19214 6724
rect 19352 6712 19380 6752
rect 19512 6749 19524 6752
rect 19558 6780 19570 6783
rect 20254 6780 20260 6792
rect 19558 6752 20260 6780
rect 19558 6749 19570 6752
rect 19512 6743 19570 6749
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 20717 6783 20775 6789
rect 20717 6749 20729 6783
rect 20763 6780 20775 6783
rect 22094 6780 22100 6792
rect 20763 6752 22100 6780
rect 20763 6749 20775 6752
rect 20717 6743 20775 6749
rect 22094 6740 22100 6752
rect 22152 6740 22158 6792
rect 19208 6684 19380 6712
rect 19208 6672 19214 6684
rect 19426 6672 19432 6724
rect 19484 6712 19490 6724
rect 19794 6712 19800 6724
rect 19484 6684 19800 6712
rect 19484 6672 19490 6684
rect 19794 6672 19800 6684
rect 19852 6712 19858 6724
rect 22462 6712 22468 6724
rect 19852 6684 22468 6712
rect 19852 6672 19858 6684
rect 22462 6672 22468 6684
rect 22520 6672 22526 6724
rect 20254 6644 20260 6656
rect 17920 6616 17965 6644
rect 18984 6616 20260 6644
rect 17920 6604 17926 6616
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 20438 6604 20444 6656
rect 20496 6644 20502 6656
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 20496 6616 20637 6644
rect 20496 6604 20502 6616
rect 20625 6613 20637 6616
rect 20671 6613 20683 6647
rect 20625 6607 20683 6613
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1627 6412 3188 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 2590 6332 2596 6384
rect 2648 6372 2654 6384
rect 2694 6375 2752 6381
rect 2694 6372 2706 6375
rect 2648 6344 2706 6372
rect 2648 6332 2654 6344
rect 2694 6341 2706 6344
rect 2740 6341 2752 6375
rect 2694 6335 2752 6341
rect 2958 6332 2964 6384
rect 3016 6372 3022 6384
rect 3160 6372 3188 6412
rect 3234 6400 3240 6452
rect 3292 6440 3298 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 3292 6412 6009 6440
rect 3292 6400 3298 6412
rect 5997 6409 6009 6412
rect 6043 6409 6055 6443
rect 6454 6440 6460 6452
rect 5997 6403 6055 6409
rect 6104 6412 6460 6440
rect 3596 6375 3654 6381
rect 3596 6372 3608 6375
rect 3016 6344 3608 6372
rect 3016 6332 3022 6344
rect 3596 6341 3608 6344
rect 3642 6372 3654 6375
rect 3694 6372 3700 6384
rect 3642 6344 3700 6372
rect 3642 6341 3654 6344
rect 3596 6335 3654 6341
rect 3694 6332 3700 6344
rect 3752 6332 3758 6384
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 4982 6372 4988 6384
rect 4120 6344 4988 6372
rect 4120 6332 4126 6344
rect 4982 6332 4988 6344
rect 5040 6332 5046 6384
rect 6104 6316 6132 6412
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 6546 6400 6552 6452
rect 6604 6440 6610 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 6604 6412 6745 6440
rect 6604 6400 6610 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 6825 6443 6883 6449
rect 6825 6409 6837 6443
rect 6871 6440 6883 6443
rect 7193 6443 7251 6449
rect 7193 6440 7205 6443
rect 6871 6412 7205 6440
rect 6871 6409 6883 6412
rect 6825 6403 6883 6409
rect 7193 6409 7205 6412
rect 7239 6409 7251 6443
rect 7374 6440 7380 6452
rect 7193 6403 7251 6409
rect 7300 6412 7380 6440
rect 6270 6332 6276 6384
rect 6328 6372 6334 6384
rect 6328 6344 6776 6372
rect 6328 6332 6334 6344
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2924 6276 3065 6304
rect 2924 6264 2930 6276
rect 3053 6273 3065 6276
rect 3099 6273 3111 6307
rect 3326 6304 3332 6316
rect 3287 6276 3332 6304
rect 3053 6267 3111 6273
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 4154 6304 4160 6316
rect 3436 6276 4160 6304
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 3234 6236 3240 6248
rect 3007 6208 3240 6236
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 3234 6196 3240 6208
rect 3292 6236 3298 6248
rect 3436 6236 3464 6276
rect 4154 6264 4160 6276
rect 4212 6264 4218 6316
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6304 5779 6307
rect 6086 6304 6092 6316
rect 5767 6276 6092 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6748 6304 6776 6344
rect 7006 6332 7012 6384
rect 7064 6332 7070 6384
rect 7024 6304 7052 6332
rect 7300 6304 7328 6412
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 7650 6440 7656 6452
rect 7611 6412 7656 6440
rect 7650 6400 7656 6412
rect 7708 6400 7714 6452
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 8386 6440 8392 6452
rect 7800 6412 8156 6440
rect 8347 6412 8392 6440
rect 7800 6400 7806 6412
rect 7558 6372 7564 6384
rect 7519 6344 7564 6372
rect 7558 6332 7564 6344
rect 7616 6332 7622 6384
rect 8128 6372 8156 6412
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 8481 6443 8539 6449
rect 8481 6409 8493 6443
rect 8527 6440 8539 6443
rect 8662 6440 8668 6452
rect 8527 6412 8668 6440
rect 8527 6409 8539 6412
rect 8481 6403 8539 6409
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 9769 6443 9827 6449
rect 9769 6440 9781 6443
rect 9355 6412 9781 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 9769 6409 9781 6412
rect 9815 6409 9827 6443
rect 9769 6403 9827 6409
rect 10229 6443 10287 6449
rect 10229 6409 10241 6443
rect 10275 6440 10287 6443
rect 10597 6443 10655 6449
rect 10597 6440 10609 6443
rect 10275 6412 10609 6440
rect 10275 6409 10287 6412
rect 10229 6403 10287 6409
rect 10597 6409 10609 6412
rect 10643 6409 10655 6443
rect 10962 6440 10968 6452
rect 10923 6412 10968 6440
rect 10597 6403 10655 6409
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 11517 6443 11575 6449
rect 11112 6412 11157 6440
rect 11112 6400 11118 6412
rect 11517 6409 11529 6443
rect 11563 6409 11575 6443
rect 11517 6403 11575 6409
rect 11977 6443 12035 6449
rect 11977 6409 11989 6443
rect 12023 6440 12035 6443
rect 12618 6440 12624 6452
rect 12023 6412 12624 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 10137 6375 10195 6381
rect 8128 6344 9628 6372
rect 6236 6276 6281 6304
rect 6748 6276 7328 6304
rect 7392 6276 8616 6304
rect 6236 6264 6242 6276
rect 3292 6208 3464 6236
rect 3292 6196 3298 6208
rect 4706 6196 4712 6248
rect 4764 6236 4770 6248
rect 4801 6239 4859 6245
rect 4801 6236 4813 6239
rect 4764 6208 4813 6236
rect 4764 6196 4770 6208
rect 4801 6205 4813 6208
rect 4847 6205 4859 6239
rect 4801 6199 4859 6205
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6236 5135 6239
rect 5626 6236 5632 6248
rect 5123 6208 5632 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 5736 6208 6776 6236
rect 5258 6128 5264 6180
rect 5316 6168 5322 6180
rect 5736 6168 5764 6208
rect 6748 6168 6776 6208
rect 6822 6196 6828 6248
rect 6880 6236 6886 6248
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6880 6208 7021 6236
rect 6880 6196 6886 6208
rect 7009 6205 7021 6208
rect 7055 6236 7067 6239
rect 7392 6236 7420 6276
rect 7055 6208 7420 6236
rect 7055 6205 7067 6208
rect 7009 6199 7067 6205
rect 7558 6196 7564 6248
rect 7616 6236 7622 6248
rect 7745 6239 7803 6245
rect 7745 6236 7757 6239
rect 7616 6208 7757 6236
rect 7616 6196 7622 6208
rect 7745 6205 7757 6208
rect 7791 6236 7803 6239
rect 7834 6236 7840 6248
rect 7791 6208 7840 6236
rect 7791 6205 7803 6208
rect 7745 6199 7803 6205
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 8588 6245 8616 6276
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 8938 6304 8944 6316
rect 8720 6276 8944 6304
rect 8720 6264 8726 6276
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9490 6304 9496 6316
rect 9048 6276 9496 6304
rect 9048 6245 9076 6276
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 9600 6304 9628 6344
rect 10137 6341 10149 6375
rect 10183 6372 10195 6375
rect 11532 6372 11560 6403
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 13262 6440 13268 6452
rect 13223 6412 13268 6440
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 13541 6443 13599 6449
rect 13541 6440 13553 6443
rect 13412 6412 13553 6440
rect 13412 6400 13418 6412
rect 13541 6409 13553 6412
rect 13587 6440 13599 6443
rect 15565 6443 15623 6449
rect 13587 6412 14688 6440
rect 13587 6409 13599 6412
rect 13541 6403 13599 6409
rect 13814 6372 13820 6384
rect 10183 6344 11560 6372
rect 11624 6344 13820 6372
rect 10183 6341 10195 6344
rect 10137 6335 10195 6341
rect 11624 6304 11652 6344
rect 13814 6332 13820 6344
rect 13872 6332 13878 6384
rect 14084 6375 14142 6381
rect 14084 6341 14096 6375
rect 14130 6372 14142 6375
rect 14182 6372 14188 6384
rect 14130 6344 14188 6372
rect 14130 6341 14142 6344
rect 14084 6335 14142 6341
rect 14182 6332 14188 6344
rect 14240 6332 14246 6384
rect 9600 6276 11652 6304
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 12345 6307 12403 6313
rect 12345 6304 12357 6307
rect 11931 6276 12357 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 12345 6273 12357 6276
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 12710 6264 12716 6316
rect 12768 6304 12774 6316
rect 13354 6304 13360 6316
rect 12768 6276 13360 6304
rect 12768 6264 12774 6276
rect 13354 6264 13360 6276
rect 13412 6264 13418 6316
rect 13906 6264 13912 6316
rect 13964 6264 13970 6316
rect 14660 6304 14688 6412
rect 15565 6409 15577 6443
rect 15611 6440 15623 6443
rect 15746 6440 15752 6452
rect 15611 6412 15752 6440
rect 15611 6409 15623 6412
rect 15565 6403 15623 6409
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 16942 6440 16948 6452
rect 16903 6412 16948 6440
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 17497 6443 17555 6449
rect 17497 6440 17509 6443
rect 17083 6412 17509 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 17497 6409 17509 6412
rect 17543 6409 17555 6443
rect 17497 6403 17555 6409
rect 18506 6400 18512 6452
rect 18564 6440 18570 6452
rect 18693 6443 18751 6449
rect 18693 6440 18705 6443
rect 18564 6412 18705 6440
rect 18564 6400 18570 6412
rect 18693 6409 18705 6412
rect 18739 6409 18751 6443
rect 18966 6440 18972 6452
rect 18927 6412 18972 6440
rect 18693 6403 18751 6409
rect 18966 6400 18972 6412
rect 19024 6400 19030 6452
rect 19337 6443 19395 6449
rect 19337 6409 19349 6443
rect 19383 6440 19395 6443
rect 19518 6440 19524 6452
rect 19383 6412 19524 6440
rect 19383 6409 19395 6412
rect 19337 6403 19395 6409
rect 19518 6400 19524 6412
rect 19576 6400 19582 6452
rect 19797 6443 19855 6449
rect 19797 6409 19809 6443
rect 19843 6409 19855 6443
rect 20254 6440 20260 6452
rect 20215 6412 20260 6440
rect 19797 6403 19855 6409
rect 14826 6332 14832 6384
rect 14884 6372 14890 6384
rect 15657 6375 15715 6381
rect 15657 6372 15669 6375
rect 14884 6344 15669 6372
rect 14884 6332 14890 6344
rect 15657 6341 15669 6344
rect 15703 6341 15715 6375
rect 15657 6335 15715 6341
rect 16114 6332 16120 6384
rect 16172 6372 16178 6384
rect 19058 6372 19064 6384
rect 16172 6344 18184 6372
rect 16172 6332 16178 6344
rect 16209 6307 16267 6313
rect 14660 6276 15516 6304
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6205 9091 6239
rect 9214 6236 9220 6248
rect 9175 6208 9220 6236
rect 9033 6199 9091 6205
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 10410 6236 10416 6248
rect 10371 6208 10416 6236
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 11146 6236 11152 6248
rect 10520 6208 11152 6236
rect 5316 6140 5764 6168
rect 5920 6140 6684 6168
rect 6748 6140 7604 6168
rect 5316 6128 5322 6140
rect 1486 6100 1492 6112
rect 1447 6072 1492 6100
rect 1486 6060 1492 6072
rect 1544 6060 1550 6112
rect 2314 6060 2320 6112
rect 2372 6100 2378 6112
rect 3142 6100 3148 6112
rect 2372 6072 3148 6100
rect 2372 6060 2378 6072
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 4709 6103 4767 6109
rect 4709 6069 4721 6103
rect 4755 6100 4767 6103
rect 4982 6100 4988 6112
rect 4755 6072 4988 6100
rect 4755 6069 4767 6072
rect 4709 6063 4767 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5074 6060 5080 6112
rect 5132 6100 5138 6112
rect 5276 6100 5304 6128
rect 5920 6109 5948 6140
rect 5132 6072 5304 6100
rect 5905 6103 5963 6109
rect 5132 6060 5138 6072
rect 5905 6069 5917 6103
rect 5951 6069 5963 6103
rect 5905 6063 5963 6069
rect 6365 6103 6423 6109
rect 6365 6069 6377 6103
rect 6411 6100 6423 6103
rect 6546 6100 6552 6112
rect 6411 6072 6552 6100
rect 6411 6069 6423 6072
rect 6365 6063 6423 6069
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 6656 6100 6684 6140
rect 7466 6100 7472 6112
rect 6656 6072 7472 6100
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 7576 6100 7604 6140
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 9306 6168 9312 6180
rect 8812 6140 9312 6168
rect 8812 6128 8818 6140
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 10134 6128 10140 6180
rect 10192 6168 10198 6180
rect 10520 6168 10548 6208
rect 11146 6196 11152 6208
rect 11204 6236 11210 6248
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 11204 6208 12081 6236
rect 11204 6196 11210 6208
rect 12069 6205 12081 6208
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 13817 6239 13875 6245
rect 12492 6208 13676 6236
rect 12492 6196 12498 6208
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 10192 6140 10548 6168
rect 11072 6140 12817 6168
rect 10192 6128 10198 6140
rect 7834 6100 7840 6112
rect 7576 6072 7840 6100
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8021 6103 8079 6109
rect 8021 6069 8033 6103
rect 8067 6100 8079 6103
rect 8294 6100 8300 6112
rect 8067 6072 8300 6100
rect 8067 6069 8079 6072
rect 8021 6063 8079 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 10594 6100 10600 6112
rect 9723 6072 10600 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 10778 6060 10784 6112
rect 10836 6100 10842 6112
rect 11072 6100 11100 6140
rect 12805 6137 12817 6140
rect 12851 6137 12863 6171
rect 12805 6131 12863 6137
rect 10836 6072 11100 6100
rect 10836 6060 10842 6072
rect 12618 6060 12624 6112
rect 12676 6100 12682 6112
rect 12713 6103 12771 6109
rect 12713 6100 12725 6103
rect 12676 6072 12725 6100
rect 12676 6060 12682 6072
rect 12713 6069 12725 6072
rect 12759 6100 12771 6103
rect 12894 6100 12900 6112
rect 12759 6072 12900 6100
rect 12759 6069 12771 6072
rect 12713 6063 12771 6069
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13081 6103 13139 6109
rect 13081 6069 13093 6103
rect 13127 6100 13139 6103
rect 13354 6100 13360 6112
rect 13127 6072 13360 6100
rect 13127 6069 13139 6072
rect 13081 6063 13139 6069
rect 13354 6060 13360 6072
rect 13412 6060 13418 6112
rect 13648 6100 13676 6208
rect 13817 6205 13829 6239
rect 13863 6236 13875 6239
rect 13924 6236 13952 6264
rect 13863 6208 13952 6236
rect 15381 6239 15439 6245
rect 13863 6205 13875 6208
rect 13817 6199 13875 6205
rect 15381 6205 15393 6239
rect 15427 6205 15439 6239
rect 15488 6236 15516 6276
rect 16209 6273 16221 6307
rect 16255 6304 16267 6307
rect 16390 6304 16396 6316
rect 16255 6276 16396 6304
rect 16255 6273 16267 6276
rect 16209 6267 16267 6273
rect 16390 6264 16396 6276
rect 16448 6304 16454 6316
rect 17218 6304 17224 6316
rect 16448 6276 17224 6304
rect 16448 6264 16454 6276
rect 17218 6264 17224 6276
rect 17276 6304 17282 6316
rect 17678 6304 17684 6316
rect 17276 6276 17684 6304
rect 17276 6264 17282 6276
rect 17678 6264 17684 6276
rect 17736 6264 17742 6316
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 18046 6304 18052 6316
rect 17911 6276 18052 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 18156 6304 18184 6344
rect 18616 6344 19064 6372
rect 18517 6307 18575 6313
rect 18156 6276 18368 6304
rect 16482 6236 16488 6248
rect 15488 6208 16488 6236
rect 15381 6199 15439 6205
rect 15194 6168 15200 6180
rect 15107 6140 15200 6168
rect 15194 6128 15200 6140
rect 15252 6168 15258 6180
rect 15396 6168 15424 6199
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6236 16911 6239
rect 17310 6236 17316 6248
rect 16899 6208 17316 6236
rect 16899 6205 16911 6208
rect 16853 6199 16911 6205
rect 17310 6196 17316 6208
rect 17368 6196 17374 6248
rect 17494 6196 17500 6248
rect 17552 6236 17558 6248
rect 17957 6239 18015 6245
rect 17957 6236 17969 6239
rect 17552 6208 17969 6236
rect 17552 6196 17558 6208
rect 17957 6205 17969 6208
rect 18003 6205 18015 6239
rect 18138 6236 18144 6248
rect 18099 6208 18144 6236
rect 17957 6199 18015 6205
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 18340 6236 18368 6276
rect 18517 6273 18529 6307
rect 18563 6304 18575 6307
rect 18616 6304 18644 6344
rect 19058 6332 19064 6344
rect 19116 6332 19122 6384
rect 19812 6372 19840 6403
rect 20254 6400 20260 6412
rect 20312 6440 20318 6452
rect 20993 6443 21051 6449
rect 20993 6440 21005 6443
rect 20312 6412 21005 6440
rect 20312 6400 20318 6412
rect 20993 6409 21005 6412
rect 21039 6409 21051 6443
rect 20993 6403 21051 6409
rect 21174 6400 21180 6452
rect 21232 6440 21238 6452
rect 21361 6443 21419 6449
rect 21361 6440 21373 6443
rect 21232 6412 21373 6440
rect 21232 6400 21238 6412
rect 21361 6409 21373 6412
rect 21407 6409 21419 6443
rect 21361 6403 21419 6409
rect 19168 6344 19840 6372
rect 20165 6375 20223 6381
rect 18563 6276 18644 6304
rect 18563 6273 18575 6276
rect 18517 6267 18575 6273
rect 18782 6264 18788 6316
rect 18840 6304 18846 6316
rect 18840 6276 18885 6304
rect 18840 6264 18846 6276
rect 19168 6236 19196 6344
rect 20165 6341 20177 6375
rect 20211 6372 20223 6375
rect 20806 6372 20812 6384
rect 20211 6344 20812 6372
rect 20211 6341 20223 6344
rect 20165 6335 20223 6341
rect 20806 6332 20812 6344
rect 20864 6332 20870 6384
rect 19334 6264 19340 6316
rect 19392 6304 19398 6316
rect 20438 6304 20444 6316
rect 19392 6276 20444 6304
rect 19392 6264 19398 6276
rect 19426 6236 19432 6248
rect 18340 6208 18460 6236
rect 16206 6168 16212 6180
rect 15252 6140 15424 6168
rect 15488 6140 16212 6168
rect 15252 6128 15258 6140
rect 15488 6100 15516 6140
rect 16206 6128 16212 6140
rect 16264 6128 16270 6180
rect 18432 6168 18460 6208
rect 18708 6208 19196 6236
rect 19387 6208 19432 6236
rect 18708 6168 18736 6208
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 19628 6245 19656 6276
rect 20438 6264 20444 6276
rect 20496 6264 20502 6316
rect 20824 6276 21036 6304
rect 19613 6239 19671 6245
rect 19613 6205 19625 6239
rect 19659 6205 19671 6239
rect 19613 6199 19671 6205
rect 20349 6239 20407 6245
rect 20349 6205 20361 6239
rect 20395 6236 20407 6239
rect 20530 6236 20536 6248
rect 20395 6208 20536 6236
rect 20395 6205 20407 6208
rect 20349 6199 20407 6205
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 20714 6236 20720 6248
rect 20675 6208 20720 6236
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 18432 6140 18736 6168
rect 19058 6128 19064 6180
rect 19116 6168 19122 6180
rect 19886 6168 19892 6180
rect 19116 6140 19892 6168
rect 19116 6128 19122 6140
rect 19886 6128 19892 6140
rect 19944 6128 19950 6180
rect 20162 6128 20168 6180
rect 20220 6168 20226 6180
rect 20824 6168 20852 6276
rect 20901 6239 20959 6245
rect 20901 6205 20913 6239
rect 20947 6205 20959 6239
rect 21008 6236 21036 6276
rect 21453 6239 21511 6245
rect 21453 6236 21465 6239
rect 21008 6208 21465 6236
rect 20901 6199 20959 6205
rect 21453 6205 21465 6208
rect 21499 6205 21511 6239
rect 21453 6199 21511 6205
rect 20220 6140 20852 6168
rect 20220 6128 20226 6140
rect 16022 6100 16028 6112
rect 13648 6072 15516 6100
rect 15983 6072 16028 6100
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 16114 6060 16120 6112
rect 16172 6100 16178 6112
rect 17310 6100 17316 6112
rect 16172 6072 17316 6100
rect 16172 6060 16178 6072
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 17405 6103 17463 6109
rect 17405 6069 17417 6103
rect 17451 6100 17463 6103
rect 17678 6100 17684 6112
rect 17451 6072 17684 6100
rect 17451 6069 17463 6072
rect 17405 6063 17463 6069
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 18322 6060 18328 6112
rect 18380 6100 18386 6112
rect 18380 6072 18425 6100
rect 18380 6060 18386 6072
rect 18598 6060 18604 6112
rect 18656 6100 18662 6112
rect 20916 6100 20944 6199
rect 18656 6072 20944 6100
rect 18656 6060 18662 6072
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 1949 5899 2007 5905
rect 1949 5896 1961 5899
rect 1544 5868 1961 5896
rect 1544 5856 1550 5868
rect 1949 5865 1961 5868
rect 1995 5865 2007 5899
rect 1949 5859 2007 5865
rect 2985 5868 3464 5896
rect 934 5788 940 5840
rect 992 5828 998 5840
rect 992 5800 1532 5828
rect 992 5788 998 5800
rect 1394 5720 1400 5772
rect 1452 5720 1458 5772
rect 1412 5624 1440 5720
rect 1504 5692 1532 5800
rect 1670 5720 1676 5772
rect 1728 5760 1734 5772
rect 2133 5763 2191 5769
rect 2133 5760 2145 5763
rect 1728 5732 2145 5760
rect 1728 5720 1734 5732
rect 2133 5729 2145 5732
rect 2179 5760 2191 5763
rect 2590 5760 2596 5772
rect 2179 5732 2596 5760
rect 2179 5729 2191 5732
rect 2133 5723 2191 5729
rect 2590 5720 2596 5732
rect 2648 5760 2654 5772
rect 2985 5760 3013 5868
rect 3142 5788 3148 5840
rect 3200 5828 3206 5840
rect 3326 5828 3332 5840
rect 3200 5800 3332 5828
rect 3200 5788 3206 5800
rect 3326 5788 3332 5800
rect 3384 5788 3390 5840
rect 3436 5828 3464 5868
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 3605 5899 3663 5905
rect 3605 5896 3617 5899
rect 3568 5868 3617 5896
rect 3568 5856 3574 5868
rect 3605 5865 3617 5868
rect 3651 5865 3663 5899
rect 5810 5896 5816 5908
rect 3605 5859 3663 5865
rect 4080 5868 5816 5896
rect 4080 5828 4108 5868
rect 5810 5856 5816 5868
rect 5868 5856 5874 5908
rect 5902 5856 5908 5908
rect 5960 5896 5966 5908
rect 6365 5899 6423 5905
rect 6365 5896 6377 5899
rect 5960 5868 6377 5896
rect 5960 5856 5966 5868
rect 6365 5865 6377 5868
rect 6411 5865 6423 5899
rect 6365 5859 6423 5865
rect 6454 5856 6460 5908
rect 6512 5896 6518 5908
rect 10042 5896 10048 5908
rect 6512 5868 10048 5896
rect 6512 5856 6518 5868
rect 10042 5856 10048 5868
rect 10100 5896 10106 5908
rect 10321 5899 10379 5905
rect 10100 5868 10272 5896
rect 10100 5856 10106 5868
rect 3436 5800 4108 5828
rect 5994 5788 6000 5840
rect 6052 5828 6058 5840
rect 7193 5831 7251 5837
rect 7193 5828 7205 5831
rect 6052 5800 7205 5828
rect 6052 5788 6058 5800
rect 7193 5797 7205 5800
rect 7239 5797 7251 5831
rect 7193 5791 7251 5797
rect 7392 5800 7788 5828
rect 2648 5732 3013 5760
rect 3053 5763 3111 5769
rect 2648 5720 2654 5732
rect 3053 5729 3065 5763
rect 3099 5760 3111 5763
rect 4430 5760 4436 5772
rect 3099 5732 4292 5760
rect 4391 5732 4436 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 1765 5695 1823 5701
rect 1765 5692 1777 5695
rect 1504 5664 1777 5692
rect 1765 5661 1777 5664
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3237 5695 3295 5701
rect 3237 5692 3249 5695
rect 3200 5664 3249 5692
rect 3200 5652 3206 5664
rect 3237 5661 3249 5664
rect 3283 5661 3295 5695
rect 3786 5692 3792 5704
rect 3747 5664 3792 5692
rect 3237 5655 3295 5661
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4154 5692 4160 5704
rect 4115 5664 4160 5692
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4264 5692 4292 5732
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 5626 5720 5632 5772
rect 5684 5760 5690 5772
rect 6917 5763 6975 5769
rect 6917 5760 6929 5763
rect 5684 5732 6929 5760
rect 5684 5720 5690 5732
rect 6917 5729 6929 5732
rect 6963 5760 6975 5763
rect 7392 5760 7420 5800
rect 7760 5769 7788 5800
rect 7834 5788 7840 5840
rect 7892 5828 7898 5840
rect 10244 5828 10272 5868
rect 10321 5865 10333 5899
rect 10367 5896 10379 5899
rect 10410 5896 10416 5908
rect 10367 5868 10416 5896
rect 10367 5865 10379 5868
rect 10321 5859 10379 5865
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 10781 5899 10839 5905
rect 10781 5865 10793 5899
rect 10827 5896 10839 5899
rect 10962 5896 10968 5908
rect 10827 5868 10968 5896
rect 10827 5865 10839 5868
rect 10781 5859 10839 5865
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 11054 5856 11060 5908
rect 11112 5896 11118 5908
rect 11149 5899 11207 5905
rect 11149 5896 11161 5899
rect 11112 5868 11161 5896
rect 11112 5856 11118 5868
rect 11149 5865 11161 5868
rect 11195 5865 11207 5899
rect 11149 5859 11207 5865
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 12434 5896 12440 5908
rect 11388 5868 12440 5896
rect 11388 5856 11394 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 16485 5899 16543 5905
rect 12676 5868 15700 5896
rect 12676 5856 12682 5868
rect 11790 5828 11796 5840
rect 7892 5800 8331 5828
rect 10244 5800 11796 5828
rect 7892 5788 7898 5800
rect 6963 5732 7420 5760
rect 7745 5763 7803 5769
rect 6963 5729 6975 5732
rect 6917 5723 6975 5729
rect 7745 5729 7757 5763
rect 7791 5729 7803 5763
rect 7745 5723 7803 5729
rect 4706 5701 4712 5704
rect 4700 5692 4712 5701
rect 4264 5664 4568 5692
rect 4667 5664 4712 5692
rect 1489 5627 1547 5633
rect 1489 5624 1501 5627
rect 1412 5596 1501 5624
rect 1489 5593 1501 5596
rect 1535 5593 1547 5627
rect 1489 5587 1547 5593
rect 1673 5627 1731 5633
rect 1673 5593 1685 5627
rect 1719 5624 1731 5627
rect 2222 5624 2228 5636
rect 1719 5596 2228 5624
rect 1719 5593 1731 5596
rect 1673 5587 1731 5593
rect 2222 5584 2228 5596
rect 2280 5584 2286 5636
rect 2317 5627 2375 5633
rect 2317 5593 2329 5627
rect 2363 5624 2375 5627
rect 3050 5624 3056 5636
rect 2363 5596 3056 5624
rect 2363 5593 2375 5596
rect 2317 5587 2375 5593
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 4246 5624 4252 5636
rect 3160 5596 4252 5624
rect 2130 5516 2136 5568
rect 2188 5556 2194 5568
rect 2409 5559 2467 5565
rect 2409 5556 2421 5559
rect 2188 5528 2421 5556
rect 2188 5516 2194 5528
rect 2409 5525 2421 5528
rect 2455 5525 2467 5559
rect 2409 5519 2467 5525
rect 2774 5516 2780 5568
rect 2832 5556 2838 5568
rect 3160 5565 3188 5596
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 4540 5624 4568 5664
rect 4700 5655 4712 5664
rect 4706 5652 4712 5655
rect 4764 5652 4770 5704
rect 5718 5652 5724 5704
rect 5776 5692 5782 5704
rect 5905 5695 5963 5701
rect 5905 5692 5917 5695
rect 5776 5664 5917 5692
rect 5776 5652 5782 5664
rect 5905 5661 5917 5664
rect 5951 5661 5963 5695
rect 6454 5692 6460 5704
rect 5905 5655 5963 5661
rect 6012 5664 6460 5692
rect 4982 5624 4988 5636
rect 4540 5596 4988 5624
rect 4982 5584 4988 5596
rect 5040 5584 5046 5636
rect 3145 5559 3203 5565
rect 2832 5528 2877 5556
rect 2832 5516 2838 5528
rect 3145 5525 3157 5559
rect 3191 5525 3203 5559
rect 3145 5519 3203 5525
rect 3786 5516 3792 5568
rect 3844 5556 3850 5568
rect 3973 5559 4031 5565
rect 3973 5556 3985 5559
rect 3844 5528 3985 5556
rect 3844 5516 3850 5528
rect 3973 5525 3985 5528
rect 4019 5525 4031 5559
rect 3973 5519 4031 5525
rect 4341 5559 4399 5565
rect 4341 5525 4353 5559
rect 4387 5556 4399 5559
rect 6012 5556 6040 5664
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5692 6883 5695
rect 7190 5692 7196 5704
rect 6871 5664 7196 5692
rect 6871 5661 6883 5664
rect 6825 5655 6883 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 6914 5624 6920 5636
rect 6104 5596 6920 5624
rect 6104 5565 6132 5596
rect 6914 5584 6920 5596
rect 6972 5584 6978 5636
rect 7561 5627 7619 5633
rect 7561 5593 7573 5627
rect 7607 5624 7619 5627
rect 8110 5624 8116 5636
rect 7607 5596 8116 5624
rect 7607 5593 7619 5596
rect 7561 5587 7619 5593
rect 8110 5584 8116 5596
rect 8168 5584 8174 5636
rect 4387 5528 6040 5556
rect 6089 5559 6147 5565
rect 4387 5525 4399 5528
rect 4341 5519 4399 5525
rect 6089 5525 6101 5559
rect 6135 5525 6147 5559
rect 6270 5556 6276 5568
rect 6231 5528 6276 5556
rect 6089 5519 6147 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 6362 5516 6368 5568
rect 6420 5556 6426 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6420 5528 6745 5556
rect 6420 5516 6426 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 7006 5516 7012 5568
rect 7064 5556 7070 5568
rect 7653 5559 7711 5565
rect 7653 5556 7665 5559
rect 7064 5528 7665 5556
rect 7064 5516 7070 5528
rect 7653 5525 7665 5528
rect 7699 5556 7711 5559
rect 7834 5556 7840 5568
rect 7699 5528 7840 5556
rect 7699 5525 7711 5528
rect 7653 5519 7711 5525
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 8021 5559 8079 5565
rect 8021 5525 8033 5559
rect 8067 5556 8079 5559
rect 8202 5556 8208 5568
rect 8067 5528 8208 5556
rect 8067 5525 8079 5528
rect 8021 5519 8079 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 8303 5556 8331 5800
rect 8665 5763 8723 5769
rect 8665 5729 8677 5763
rect 8711 5729 8723 5763
rect 8938 5760 8944 5772
rect 8899 5732 8944 5760
rect 8665 5723 8723 5729
rect 8478 5692 8484 5704
rect 8439 5664 8484 5692
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 8680 5692 8708 5723
rect 8938 5720 8944 5732
rect 8996 5720 9002 5772
rect 10778 5720 10784 5772
rect 10836 5720 10842 5772
rect 9030 5692 9036 5704
rect 8680 5664 9036 5692
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9197 5695 9255 5701
rect 9197 5661 9209 5695
rect 9243 5692 9255 5695
rect 10134 5692 10140 5704
rect 9243 5664 10140 5692
rect 9243 5661 9255 5664
rect 9197 5655 9255 5661
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 10796 5692 10824 5720
rect 10643 5664 10824 5692
rect 10888 5692 10916 5800
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 13817 5831 13875 5837
rect 13817 5828 13829 5831
rect 13096 5800 13829 5828
rect 11146 5720 11152 5772
rect 11204 5760 11210 5772
rect 13096 5769 13124 5800
rect 13817 5797 13829 5800
rect 13863 5828 13875 5831
rect 14274 5828 14280 5840
rect 13863 5800 14280 5828
rect 13863 5797 13875 5800
rect 13817 5791 13875 5797
rect 14274 5788 14280 5800
rect 14332 5788 14338 5840
rect 15562 5828 15568 5840
rect 15523 5800 15568 5828
rect 15562 5788 15568 5800
rect 15620 5788 15626 5840
rect 11701 5763 11759 5769
rect 11701 5760 11713 5763
rect 11204 5732 11713 5760
rect 11204 5720 11210 5732
rect 11701 5729 11713 5732
rect 11747 5729 11759 5763
rect 11701 5723 11759 5729
rect 13081 5763 13139 5769
rect 13081 5729 13093 5763
rect 13127 5729 13139 5763
rect 13081 5723 13139 5729
rect 13265 5763 13323 5769
rect 13265 5729 13277 5763
rect 13311 5760 13323 5763
rect 13722 5760 13728 5772
rect 13311 5732 13728 5760
rect 13311 5729 13323 5732
rect 13265 5723 13323 5729
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 10888 5664 11621 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 11716 5692 11744 5723
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 11716 5664 12173 5692
rect 11609 5655 11667 5661
rect 12161 5661 12173 5664
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 8389 5627 8447 5633
rect 8389 5593 8401 5627
rect 8435 5624 8447 5627
rect 9582 5624 9588 5636
rect 8435 5596 9588 5624
rect 8435 5593 8447 5596
rect 8389 5587 8447 5593
rect 9582 5584 9588 5596
rect 9640 5584 9646 5636
rect 9858 5584 9864 5636
rect 9916 5624 9922 5636
rect 10612 5624 10640 5655
rect 12250 5652 12256 5704
rect 12308 5692 12314 5704
rect 12989 5695 13047 5701
rect 12989 5692 13001 5695
rect 12308 5664 13001 5692
rect 12308 5652 12314 5664
rect 12989 5661 13001 5664
rect 13035 5661 13047 5695
rect 12989 5655 13047 5661
rect 13633 5695 13691 5701
rect 13633 5661 13645 5695
rect 13679 5692 13691 5695
rect 13814 5692 13820 5704
rect 13679 5664 13820 5692
rect 13679 5661 13691 5664
rect 13633 5655 13691 5661
rect 13814 5652 13820 5664
rect 13872 5692 13878 5704
rect 14366 5692 14372 5704
rect 13872 5664 14372 5692
rect 13872 5652 13878 5664
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 15194 5652 15200 5704
rect 15252 5701 15258 5704
rect 15252 5692 15264 5701
rect 15473 5695 15531 5701
rect 15252 5664 15297 5692
rect 15252 5655 15264 5664
rect 15473 5661 15485 5695
rect 15519 5661 15531 5695
rect 15473 5655 15531 5661
rect 15252 5652 15258 5655
rect 9916 5596 10640 5624
rect 9916 5584 9922 5596
rect 10778 5584 10784 5636
rect 10836 5624 10842 5636
rect 11977 5627 12035 5633
rect 11977 5624 11989 5627
rect 10836 5596 11989 5624
rect 10836 5584 10842 5596
rect 11977 5593 11989 5596
rect 12023 5593 12035 5627
rect 14384 5624 14412 5652
rect 15488 5624 15516 5655
rect 14384 5596 15516 5624
rect 15672 5624 15700 5868
rect 16485 5865 16497 5899
rect 16531 5896 16543 5899
rect 16574 5896 16580 5908
rect 16531 5868 16580 5896
rect 16531 5865 16543 5868
rect 16485 5859 16543 5865
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 17678 5856 17684 5908
rect 17736 5896 17742 5908
rect 18693 5899 18751 5905
rect 17736 5868 18644 5896
rect 17736 5856 17742 5868
rect 18138 5828 18144 5840
rect 15948 5800 18144 5828
rect 15948 5769 15976 5800
rect 18138 5788 18144 5800
rect 18196 5788 18202 5840
rect 18322 5788 18328 5840
rect 18380 5788 18386 5840
rect 18616 5828 18644 5868
rect 18693 5865 18705 5899
rect 18739 5896 18751 5899
rect 18966 5896 18972 5908
rect 18739 5868 18972 5896
rect 18739 5865 18751 5868
rect 18693 5859 18751 5865
rect 18966 5856 18972 5868
rect 19024 5856 19030 5908
rect 20625 5899 20683 5905
rect 20625 5865 20637 5899
rect 20671 5896 20683 5899
rect 21082 5896 21088 5908
rect 20671 5868 21088 5896
rect 20671 5865 20683 5868
rect 20625 5859 20683 5865
rect 21082 5856 21088 5868
rect 21140 5856 21146 5908
rect 19058 5828 19064 5840
rect 18616 5800 19064 5828
rect 19058 5788 19064 5800
rect 19116 5788 19122 5840
rect 20806 5788 20812 5840
rect 20864 5828 20870 5840
rect 20864 5800 21036 5828
rect 20864 5788 20870 5800
rect 15933 5763 15991 5769
rect 15933 5729 15945 5763
rect 15979 5729 15991 5763
rect 15933 5723 15991 5729
rect 16025 5763 16083 5769
rect 16025 5729 16037 5763
rect 16071 5760 16083 5763
rect 16114 5760 16120 5772
rect 16071 5732 16120 5760
rect 16071 5729 16083 5732
rect 16025 5723 16083 5729
rect 15746 5652 15752 5704
rect 15804 5692 15810 5704
rect 16040 5692 16068 5723
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 16482 5720 16488 5772
rect 16540 5760 16546 5772
rect 17037 5763 17095 5769
rect 17037 5760 17049 5763
rect 16540 5732 17049 5760
rect 16540 5720 16546 5732
rect 17037 5729 17049 5732
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 17126 5720 17132 5772
rect 17184 5760 17190 5772
rect 17221 5763 17279 5769
rect 17221 5760 17233 5763
rect 17184 5732 17233 5760
rect 17184 5720 17190 5732
rect 17221 5729 17233 5732
rect 17267 5729 17279 5763
rect 17770 5760 17776 5772
rect 17221 5723 17279 5729
rect 17420 5732 17776 5760
rect 17420 5701 17448 5732
rect 17770 5720 17776 5732
rect 17828 5720 17834 5772
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5760 17923 5763
rect 17954 5760 17960 5772
rect 17911 5732 17960 5760
rect 17911 5729 17923 5732
rect 17865 5723 17923 5729
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 18340 5760 18368 5788
rect 18340 5732 19380 5760
rect 17405 5695 17463 5701
rect 17405 5692 17417 5695
rect 15804 5664 16068 5692
rect 16132 5688 16988 5692
rect 17052 5688 17417 5692
rect 16132 5664 17417 5688
rect 15804 5652 15810 5664
rect 16132 5624 16160 5664
rect 16960 5660 17080 5664
rect 17405 5661 17417 5664
rect 17451 5661 17463 5695
rect 17405 5655 17463 5661
rect 17678 5652 17684 5704
rect 17736 5692 17742 5704
rect 18046 5692 18052 5704
rect 17736 5664 18052 5692
rect 17736 5652 17742 5664
rect 18046 5652 18052 5664
rect 18104 5652 18110 5704
rect 18322 5652 18328 5704
rect 18380 5692 18386 5704
rect 18874 5692 18880 5704
rect 18380 5664 18880 5692
rect 18380 5652 18386 5664
rect 18874 5652 18880 5664
rect 18932 5692 18938 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 18932 5664 19257 5692
rect 18932 5652 18938 5664
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19352 5692 19380 5732
rect 21008 5704 21036 5800
rect 21100 5760 21128 5856
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 21100 5732 21281 5760
rect 21269 5729 21281 5732
rect 21315 5729 21327 5763
rect 21269 5723 21327 5729
rect 20806 5692 20812 5704
rect 19352 5664 20812 5692
rect 19245 5655 19303 5661
rect 20806 5652 20812 5664
rect 20864 5652 20870 5704
rect 20990 5652 20996 5704
rect 21048 5692 21054 5704
rect 21177 5695 21235 5701
rect 21177 5692 21189 5695
rect 21048 5664 21189 5692
rect 21048 5652 21054 5664
rect 21177 5661 21189 5664
rect 21223 5661 21235 5695
rect 21177 5655 21235 5661
rect 15672 5596 16160 5624
rect 11977 5587 12035 5593
rect 16298 5584 16304 5636
rect 16356 5624 16362 5636
rect 17494 5624 17500 5636
rect 16356 5596 17500 5624
rect 16356 5584 16362 5596
rect 17494 5584 17500 5596
rect 17552 5624 17558 5636
rect 17589 5627 17647 5633
rect 17589 5624 17601 5627
rect 17552 5596 17601 5624
rect 17552 5584 17558 5596
rect 17589 5593 17601 5596
rect 17635 5593 17647 5627
rect 18785 5627 18843 5633
rect 18785 5624 18797 5627
rect 17589 5587 17647 5593
rect 17696 5596 18797 5624
rect 10413 5559 10471 5565
rect 10413 5556 10425 5559
rect 8303 5528 10425 5556
rect 10413 5525 10425 5528
rect 10459 5525 10471 5559
rect 11054 5556 11060 5568
rect 10967 5528 11060 5556
rect 10413 5519 10471 5525
rect 11054 5516 11060 5528
rect 11112 5556 11118 5568
rect 11514 5556 11520 5568
rect 11112 5528 11520 5556
rect 11112 5516 11118 5528
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 12345 5559 12403 5565
rect 12345 5556 12357 5559
rect 11848 5528 12357 5556
rect 11848 5516 11854 5528
rect 12345 5525 12357 5528
rect 12391 5525 12403 5559
rect 12618 5556 12624 5568
rect 12579 5528 12624 5556
rect 12345 5519 12403 5525
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 13449 5559 13507 5565
rect 13449 5525 13461 5559
rect 13495 5556 13507 5559
rect 13630 5556 13636 5568
rect 13495 5528 13636 5556
rect 13495 5525 13507 5528
rect 13449 5519 13507 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 14090 5556 14096 5568
rect 14051 5528 14096 5556
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 16117 5559 16175 5565
rect 16117 5556 16129 5559
rect 15620 5528 16129 5556
rect 15620 5516 15626 5528
rect 16117 5525 16129 5528
rect 16163 5525 16175 5559
rect 16117 5519 16175 5525
rect 16574 5516 16580 5568
rect 16632 5556 16638 5568
rect 16942 5556 16948 5568
rect 16632 5528 16677 5556
rect 16903 5528 16948 5556
rect 16632 5516 16638 5528
rect 16942 5516 16948 5528
rect 17000 5516 17006 5568
rect 17310 5516 17316 5568
rect 17368 5556 17374 5568
rect 17696 5556 17724 5596
rect 18785 5593 18797 5596
rect 18831 5593 18843 5627
rect 18966 5624 18972 5636
rect 18927 5596 18972 5624
rect 18785 5587 18843 5593
rect 18966 5584 18972 5596
rect 19024 5584 19030 5636
rect 19512 5627 19570 5633
rect 19512 5593 19524 5627
rect 19558 5624 19570 5627
rect 19702 5624 19708 5636
rect 19558 5596 19708 5624
rect 19558 5593 19570 5596
rect 19512 5587 19570 5593
rect 19702 5584 19708 5596
rect 19760 5584 19766 5636
rect 22922 5624 22928 5636
rect 21100 5596 22928 5624
rect 21100 5568 21128 5596
rect 22922 5584 22928 5596
rect 22980 5584 22986 5636
rect 18046 5556 18052 5568
rect 17368 5528 17724 5556
rect 18007 5528 18052 5556
rect 17368 5516 17374 5528
rect 18046 5516 18052 5528
rect 18104 5516 18110 5568
rect 18141 5559 18199 5565
rect 18141 5525 18153 5559
rect 18187 5556 18199 5559
rect 18230 5556 18236 5568
rect 18187 5528 18236 5556
rect 18187 5525 18199 5528
rect 18141 5519 18199 5525
rect 18230 5516 18236 5528
rect 18288 5516 18294 5568
rect 18506 5556 18512 5568
rect 18467 5528 18512 5556
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 21082 5556 21088 5568
rect 20772 5528 20817 5556
rect 21043 5528 21088 5556
rect 20772 5516 20778 5528
rect 21082 5516 21088 5528
rect 21140 5516 21146 5568
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 4341 5355 4399 5361
rect 4341 5352 4353 5355
rect 3108 5324 4353 5352
rect 3108 5312 3114 5324
rect 4341 5321 4353 5324
rect 4387 5321 4399 5355
rect 4341 5315 4399 5321
rect 4709 5355 4767 5361
rect 4709 5321 4721 5355
rect 4755 5352 4767 5355
rect 5258 5352 5264 5364
rect 4755 5324 5264 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 5445 5355 5503 5361
rect 5445 5321 5457 5355
rect 5491 5352 5503 5355
rect 5718 5352 5724 5364
rect 5491 5324 5724 5352
rect 5491 5321 5503 5324
rect 5445 5315 5503 5321
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 5810 5312 5816 5364
rect 5868 5352 5874 5364
rect 5868 5324 6960 5352
rect 5868 5312 5874 5324
rect 1578 5244 1584 5296
rect 1636 5284 1642 5296
rect 2685 5287 2743 5293
rect 2685 5284 2697 5287
rect 1636 5256 2697 5284
rect 1636 5244 1642 5256
rect 2685 5253 2697 5256
rect 2731 5284 2743 5287
rect 3418 5284 3424 5296
rect 2731 5256 3424 5284
rect 2731 5253 2743 5256
rect 2685 5247 2743 5253
rect 3418 5244 3424 5256
rect 3476 5244 3482 5296
rect 3878 5244 3884 5296
rect 3936 5244 3942 5296
rect 4246 5244 4252 5296
rect 4304 5284 4310 5296
rect 4982 5284 4988 5296
rect 4304 5256 4988 5284
rect 4304 5244 4310 5256
rect 4982 5244 4988 5256
rect 5040 5284 5046 5296
rect 5905 5287 5963 5293
rect 5040 5256 5212 5284
rect 5040 5244 5046 5256
rect 1946 5216 1952 5228
rect 1907 5188 1952 5216
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 2406 5216 2412 5228
rect 2367 5188 2412 5216
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2590 5176 2596 5228
rect 2648 5216 2654 5228
rect 3125 5219 3183 5225
rect 3125 5216 3137 5219
rect 2648 5188 3137 5216
rect 2648 5176 2654 5188
rect 3125 5185 3137 5188
rect 3171 5185 3183 5219
rect 3896 5216 3924 5244
rect 5074 5216 5080 5228
rect 3896 5188 5080 5216
rect 3125 5179 3183 5185
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 5184 5225 5212 5256
rect 5905 5253 5917 5287
rect 5951 5284 5963 5287
rect 6932 5284 6960 5324
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 7193 5355 7251 5361
rect 7193 5352 7205 5355
rect 7064 5324 7205 5352
rect 7064 5312 7070 5324
rect 7193 5321 7205 5324
rect 7239 5321 7251 5355
rect 7558 5352 7564 5364
rect 7519 5324 7564 5352
rect 7193 5315 7251 5321
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 8202 5352 8208 5364
rect 8163 5324 8208 5352
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8665 5355 8723 5361
rect 8352 5324 8397 5352
rect 8352 5312 8358 5324
rect 8665 5321 8677 5355
rect 8711 5352 8723 5355
rect 9766 5352 9772 5364
rect 8711 5324 9772 5352
rect 8711 5321 8723 5324
rect 8665 5315 8723 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 10134 5352 10140 5364
rect 10095 5324 10140 5352
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10502 5312 10508 5364
rect 10560 5352 10566 5364
rect 11054 5352 11060 5364
rect 10560 5324 11060 5352
rect 10560 5312 10566 5324
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11330 5352 11336 5364
rect 11291 5324 11336 5352
rect 11330 5312 11336 5324
rect 11388 5312 11394 5364
rect 12069 5355 12127 5361
rect 12069 5321 12081 5355
rect 12115 5352 12127 5355
rect 12158 5352 12164 5364
rect 12115 5324 12164 5352
rect 12115 5321 12127 5324
rect 12069 5315 12127 5321
rect 12158 5312 12164 5324
rect 12216 5352 12222 5364
rect 12342 5352 12348 5364
rect 12216 5324 12348 5352
rect 12216 5312 12222 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 12618 5352 12624 5364
rect 12483 5324 12624 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 14553 5355 14611 5361
rect 12768 5324 14504 5352
rect 12768 5312 12774 5324
rect 7282 5284 7288 5296
rect 5951 5256 6868 5284
rect 6932 5256 7288 5284
rect 5951 5253 5963 5256
rect 5905 5247 5963 5253
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5185 5227 5219
rect 5813 5219 5871 5225
rect 5813 5216 5825 5219
rect 5169 5179 5227 5185
rect 5368 5188 5825 5216
rect 2222 5148 2228 5160
rect 2183 5120 2228 5148
rect 2222 5108 2228 5120
rect 2280 5108 2286 5160
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5117 2927 5151
rect 2869 5111 2927 5117
rect 1026 4972 1032 5024
rect 1084 5012 1090 5024
rect 2501 5015 2559 5021
rect 2501 5012 2513 5015
rect 1084 4984 2513 5012
rect 1084 4972 1090 4984
rect 2501 4981 2513 4984
rect 2547 4981 2559 5015
rect 2884 5012 2912 5111
rect 3878 5108 3884 5160
rect 3936 5148 3942 5160
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 3936 5120 4813 5148
rect 3936 5108 3942 5120
rect 4801 5117 4813 5120
rect 4847 5117 4859 5151
rect 4801 5111 4859 5117
rect 4893 5151 4951 5157
rect 4893 5117 4905 5151
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 4249 5083 4307 5089
rect 4249 5049 4261 5083
rect 4295 5080 4307 5083
rect 4706 5080 4712 5092
rect 4295 5052 4712 5080
rect 4295 5049 4307 5052
rect 4249 5043 4307 5049
rect 4706 5040 4712 5052
rect 4764 5080 4770 5092
rect 4908 5080 4936 5111
rect 5368 5089 5396 5188
rect 5813 5185 5825 5188
rect 5859 5216 5871 5219
rect 6086 5216 6092 5228
rect 5859 5188 6092 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 6086 5176 6092 5188
rect 6144 5176 6150 5228
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6733 5219 6791 5225
rect 6733 5216 6745 5219
rect 6328 5188 6745 5216
rect 6328 5176 6334 5188
rect 6733 5185 6745 5188
rect 6779 5185 6791 5219
rect 6840 5216 6868 5256
rect 7282 5244 7288 5256
rect 7340 5244 7346 5296
rect 8018 5284 8024 5296
rect 7852 5256 8024 5284
rect 7377 5219 7435 5225
rect 6840 5188 7328 5216
rect 6733 5179 6791 5185
rect 5626 5108 5632 5160
rect 5684 5148 5690 5160
rect 5997 5151 6055 5157
rect 5997 5148 6009 5151
rect 5684 5120 6009 5148
rect 5684 5108 5690 5120
rect 5997 5117 6009 5120
rect 6043 5117 6055 5151
rect 5997 5111 6055 5117
rect 4764 5052 4936 5080
rect 5353 5083 5411 5089
rect 4764 5040 4770 5052
rect 5353 5049 5365 5083
rect 5399 5049 5411 5083
rect 6012 5080 6040 5111
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6512 5120 6837 5148
rect 6512 5108 6518 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5117 6975 5151
rect 7300 5148 7328 5188
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 7558 5216 7564 5228
rect 7423 5188 7564 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 7558 5176 7564 5188
rect 7616 5216 7622 5228
rect 7742 5216 7748 5228
rect 7616 5188 7748 5216
rect 7616 5176 7622 5188
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 7852 5225 7880 5256
rect 8018 5244 8024 5256
rect 8076 5284 8082 5296
rect 10152 5284 10180 5312
rect 8076 5256 8708 5284
rect 8076 5244 8082 5256
rect 8680 5228 8708 5256
rect 8956 5256 10180 5284
rect 7837 5219 7895 5225
rect 7837 5185 7849 5219
rect 7883 5185 7895 5219
rect 8478 5216 8484 5228
rect 7837 5179 7895 5185
rect 8036 5188 8484 5216
rect 8036 5148 8064 5188
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 8662 5176 8668 5228
rect 8720 5216 8726 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8720 5188 8769 5216
rect 8720 5176 8726 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8956 5216 8984 5256
rect 9030 5225 9036 5228
rect 8757 5179 8815 5185
rect 8864 5188 8984 5216
rect 7300 5120 8064 5148
rect 8113 5151 8171 5157
rect 6917 5111 6975 5117
rect 8113 5117 8125 5151
rect 8159 5148 8171 5151
rect 8864 5148 8892 5188
rect 9024 5179 9036 5225
rect 9088 5216 9094 5228
rect 9306 5216 9312 5228
rect 9088 5188 9312 5216
rect 9030 5176 9036 5179
rect 9088 5176 9094 5188
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 9490 5176 9496 5228
rect 9548 5216 9554 5228
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 9548 5188 10241 5216
rect 9548 5176 9554 5188
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10962 5216 10968 5228
rect 10923 5188 10968 5216
rect 10229 5179 10287 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5216 11759 5219
rect 11790 5216 11796 5228
rect 11747 5188 11796 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 12529 5219 12587 5225
rect 12529 5185 12541 5219
rect 12575 5216 12587 5219
rect 12894 5216 12900 5228
rect 12575 5188 12900 5216
rect 12575 5185 12587 5188
rect 12529 5179 12587 5185
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 14102 5219 14160 5225
rect 14102 5216 14114 5219
rect 13872 5188 14114 5216
rect 13872 5176 13878 5188
rect 14102 5185 14114 5188
rect 14148 5185 14160 5219
rect 14366 5216 14372 5228
rect 14327 5188 14372 5216
rect 14102 5179 14160 5185
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 14476 5216 14504 5324
rect 14553 5321 14565 5355
rect 14599 5352 14611 5355
rect 14737 5355 14795 5361
rect 14737 5352 14749 5355
rect 14599 5324 14749 5352
rect 14599 5321 14611 5324
rect 14553 5315 14611 5321
rect 14737 5321 14749 5324
rect 14783 5352 14795 5355
rect 14918 5352 14924 5364
rect 14783 5324 14924 5352
rect 14783 5321 14795 5324
rect 14737 5315 14795 5321
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 15010 5312 15016 5364
rect 15068 5352 15074 5364
rect 15194 5352 15200 5364
rect 15068 5324 15113 5352
rect 15155 5324 15200 5352
rect 15068 5312 15074 5324
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 15654 5352 15660 5364
rect 15488 5324 15660 5352
rect 15488 5293 15516 5324
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 16025 5355 16083 5361
rect 16025 5321 16037 5355
rect 16071 5352 16083 5355
rect 16669 5355 16727 5361
rect 16669 5352 16681 5355
rect 16071 5324 16681 5352
rect 16071 5321 16083 5324
rect 16025 5315 16083 5321
rect 16669 5321 16681 5324
rect 16715 5321 16727 5355
rect 16669 5315 16727 5321
rect 17586 5312 17592 5364
rect 17644 5352 17650 5364
rect 20165 5355 20223 5361
rect 17644 5324 19196 5352
rect 17644 5312 17650 5324
rect 15473 5287 15531 5293
rect 15473 5253 15485 5287
rect 15519 5253 15531 5287
rect 15838 5284 15844 5296
rect 15473 5247 15531 5253
rect 15580 5256 15844 5284
rect 15580 5216 15608 5256
rect 15838 5244 15844 5256
rect 15896 5244 15902 5296
rect 16117 5287 16175 5293
rect 16117 5253 16129 5287
rect 16163 5284 16175 5287
rect 16390 5284 16396 5296
rect 16163 5256 16396 5284
rect 16163 5253 16175 5256
rect 16117 5247 16175 5253
rect 16390 5244 16396 5256
rect 16448 5244 16454 5296
rect 16574 5244 16580 5296
rect 16632 5284 16638 5296
rect 17037 5287 17095 5293
rect 17037 5284 17049 5287
rect 16632 5256 17049 5284
rect 16632 5244 16638 5256
rect 17037 5253 17049 5256
rect 17083 5253 17095 5287
rect 17037 5247 17095 5253
rect 17126 5244 17132 5296
rect 17184 5244 17190 5296
rect 17954 5284 17960 5296
rect 17696 5256 17960 5284
rect 14476 5188 15608 5216
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5216 15715 5219
rect 17144 5216 17172 5244
rect 15703 5188 17264 5216
rect 15703 5185 15715 5188
rect 15657 5179 15715 5185
rect 10778 5148 10784 5160
rect 8159 5120 8892 5148
rect 10739 5120 10784 5148
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 6932 5080 6960 5111
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 10873 5151 10931 5157
rect 10873 5117 10885 5151
rect 10919 5148 10931 5151
rect 11606 5148 11612 5160
rect 10919 5120 11612 5148
rect 10919 5117 10931 5120
rect 10873 5111 10931 5117
rect 6012 5052 6960 5080
rect 5353 5043 5411 5049
rect 7282 5040 7288 5092
rect 7340 5080 7346 5092
rect 8754 5080 8760 5092
rect 7340 5052 8760 5080
rect 7340 5040 7346 5052
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 10686 5040 10692 5092
rect 10744 5080 10750 5092
rect 10888 5080 10916 5111
rect 11606 5108 11612 5120
rect 11664 5108 11670 5160
rect 12345 5151 12403 5157
rect 12345 5117 12357 5151
rect 12391 5148 12403 5151
rect 12391 5120 12848 5148
rect 12391 5117 12403 5120
rect 12345 5111 12403 5117
rect 10744 5052 10916 5080
rect 10744 5040 10750 5052
rect 11054 5040 11060 5092
rect 11112 5080 11118 5092
rect 11517 5083 11575 5089
rect 11517 5080 11529 5083
rect 11112 5052 11529 5080
rect 11112 5040 11118 5052
rect 11517 5049 11529 5052
rect 11563 5080 11575 5083
rect 12250 5080 12256 5092
rect 11563 5052 12256 5080
rect 11563 5049 11575 5052
rect 11517 5043 11575 5049
rect 12250 5040 12256 5052
rect 12308 5040 12314 5092
rect 3234 5012 3240 5024
rect 2884 4984 3240 5012
rect 2501 4975 2559 4981
rect 3234 4972 3240 4984
rect 3292 5012 3298 5024
rect 4154 5012 4160 5024
rect 3292 4984 4160 5012
rect 3292 4972 3298 4984
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 5626 5012 5632 5024
rect 4672 4984 5632 5012
rect 4672 4972 4678 4984
rect 5626 4972 5632 4984
rect 5684 5012 5690 5024
rect 6178 5012 6184 5024
rect 5684 4984 6184 5012
rect 5684 4972 5690 4984
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 6362 5012 6368 5024
rect 6323 4984 6368 5012
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 7650 5012 7656 5024
rect 7611 4984 7656 5012
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 10134 5012 10140 5024
rect 7892 4984 10140 5012
rect 7892 4972 7898 4984
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 10413 5015 10471 5021
rect 10413 4981 10425 5015
rect 10459 5012 10471 5015
rect 11422 5012 11428 5024
rect 10459 4984 11428 5012
rect 10459 4981 10471 4984
rect 10413 4975 10471 4981
rect 11422 4972 11428 4984
rect 11480 4972 11486 5024
rect 11606 4972 11612 5024
rect 11664 5012 11670 5024
rect 11885 5015 11943 5021
rect 11885 5012 11897 5015
rect 11664 4984 11897 5012
rect 11664 4972 11670 4984
rect 11885 4981 11897 4984
rect 11931 5012 11943 5015
rect 12710 5012 12716 5024
rect 11931 4984 12716 5012
rect 11931 4981 11943 4984
rect 11885 4975 11943 4981
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 12820 5012 12848 5120
rect 14458 5108 14464 5160
rect 14516 5148 14522 5160
rect 15838 5148 15844 5160
rect 14516 5120 15844 5148
rect 14516 5108 14522 5120
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5148 15991 5151
rect 16758 5148 16764 5160
rect 15979 5120 16764 5148
rect 15979 5117 15991 5120
rect 15933 5111 15991 5117
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 16942 5108 16948 5160
rect 17000 5148 17006 5160
rect 17236 5157 17264 5188
rect 17696 5157 17724 5256
rect 17954 5244 17960 5256
rect 18012 5284 18018 5296
rect 19168 5284 19196 5324
rect 20165 5321 20177 5355
rect 20211 5352 20223 5355
rect 20714 5352 20720 5364
rect 20211 5324 20720 5352
rect 20211 5321 20223 5324
rect 20165 5315 20223 5321
rect 20714 5312 20720 5324
rect 20772 5312 20778 5364
rect 20257 5287 20315 5293
rect 20257 5284 20269 5287
rect 18012 5256 18460 5284
rect 19168 5256 20269 5284
rect 18012 5244 18018 5256
rect 18432 5228 18460 5256
rect 20257 5253 20269 5256
rect 20303 5253 20315 5287
rect 20257 5247 20315 5253
rect 17862 5216 17868 5228
rect 17823 5188 17868 5216
rect 17862 5176 17868 5188
rect 17920 5176 17926 5228
rect 18414 5176 18420 5228
rect 18472 5216 18478 5228
rect 18581 5219 18639 5225
rect 18581 5216 18593 5219
rect 18472 5188 18593 5216
rect 18472 5176 18478 5188
rect 18581 5185 18593 5188
rect 18627 5185 18639 5219
rect 21542 5216 21548 5228
rect 21503 5188 21548 5216
rect 18581 5179 18639 5185
rect 21542 5176 21548 5188
rect 21600 5176 21606 5228
rect 17129 5151 17187 5157
rect 17129 5148 17141 5151
rect 17000 5120 17141 5148
rect 17000 5108 17006 5120
rect 17129 5117 17141 5120
rect 17175 5117 17187 5151
rect 17129 5111 17187 5117
rect 17221 5151 17279 5157
rect 17221 5117 17233 5151
rect 17267 5117 17279 5151
rect 17221 5111 17279 5117
rect 17681 5151 17739 5157
rect 17681 5117 17693 5151
rect 17727 5117 17739 5151
rect 17681 5111 17739 5117
rect 17773 5151 17831 5157
rect 17773 5117 17785 5151
rect 17819 5117 17831 5151
rect 18322 5148 18328 5160
rect 17773 5111 17831 5117
rect 17880 5120 18328 5148
rect 12897 5083 12955 5089
rect 12897 5049 12909 5083
rect 12943 5080 12955 5083
rect 13262 5080 13268 5092
rect 12943 5052 13268 5080
rect 12943 5049 12955 5052
rect 12897 5043 12955 5049
rect 13262 5040 13268 5052
rect 13320 5040 13326 5092
rect 14366 5040 14372 5092
rect 14424 5080 14430 5092
rect 14829 5083 14887 5089
rect 14829 5080 14841 5083
rect 14424 5052 14841 5080
rect 14424 5040 14430 5052
rect 14829 5049 14841 5052
rect 14875 5049 14887 5083
rect 14829 5043 14887 5049
rect 16485 5083 16543 5089
rect 16485 5049 16497 5083
rect 16531 5080 16543 5083
rect 17788 5080 17816 5111
rect 16531 5052 17816 5080
rect 16531 5049 16543 5052
rect 16485 5043 16543 5049
rect 12986 5012 12992 5024
rect 12820 4984 12992 5012
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 15010 4972 15016 5024
rect 15068 5012 15074 5024
rect 16390 5012 16396 5024
rect 15068 4984 16396 5012
rect 15068 4972 15074 4984
rect 16390 4972 16396 4984
rect 16448 5012 16454 5024
rect 16574 5012 16580 5024
rect 16448 4984 16580 5012
rect 16448 4972 16454 4984
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 16850 4972 16856 5024
rect 16908 5012 16914 5024
rect 17880 5012 17908 5120
rect 18322 5108 18328 5120
rect 18380 5108 18386 5160
rect 20438 5148 20444 5160
rect 20399 5120 20444 5148
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 21269 5151 21327 5157
rect 21269 5117 21281 5151
rect 21315 5148 21327 5151
rect 22094 5148 22100 5160
rect 21315 5120 22100 5148
rect 21315 5117 21327 5120
rect 21269 5111 21327 5117
rect 22094 5108 22100 5120
rect 22152 5108 22158 5160
rect 19797 5083 19855 5089
rect 19797 5049 19809 5083
rect 19843 5080 19855 5083
rect 20346 5080 20352 5092
rect 19843 5052 20352 5080
rect 19843 5049 19855 5052
rect 19797 5043 19855 5049
rect 20346 5040 20352 5052
rect 20404 5040 20410 5092
rect 16908 4984 17908 5012
rect 18233 5015 18291 5021
rect 16908 4972 16914 4984
rect 18233 4981 18245 5015
rect 18279 5012 18291 5015
rect 19518 5012 19524 5024
rect 18279 4984 19524 5012
rect 18279 4981 18291 4984
rect 18233 4975 18291 4981
rect 19518 4972 19524 4984
rect 19576 4972 19582 5024
rect 19702 5012 19708 5024
rect 19663 4984 19708 5012
rect 19702 4972 19708 4984
rect 19760 4972 19766 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 1578 4808 1584 4820
rect 1539 4780 1584 4808
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2590 4808 2596 4820
rect 1995 4780 2596 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2590 4768 2596 4780
rect 2648 4768 2654 4820
rect 3326 4768 3332 4820
rect 3384 4808 3390 4820
rect 3421 4811 3479 4817
rect 3421 4808 3433 4811
rect 3384 4780 3433 4808
rect 3384 4768 3390 4780
rect 3421 4777 3433 4780
rect 3467 4777 3479 4811
rect 3421 4771 3479 4777
rect 4430 4768 4436 4820
rect 4488 4808 4494 4820
rect 4890 4808 4896 4820
rect 4488 4780 4896 4808
rect 4488 4768 4494 4780
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 5353 4811 5411 4817
rect 5353 4808 5365 4811
rect 5316 4780 5365 4808
rect 5316 4768 5322 4780
rect 5353 4777 5365 4780
rect 5399 4777 5411 4811
rect 5353 4771 5411 4777
rect 5460 4780 6408 4808
rect 1857 4743 1915 4749
rect 1857 4709 1869 4743
rect 1903 4740 1915 4743
rect 2038 4740 2044 4752
rect 1903 4712 2044 4740
rect 1903 4709 1915 4712
rect 1857 4703 1915 4709
rect 2038 4700 2044 4712
rect 2096 4700 2102 4752
rect 3878 4672 3884 4684
rect 3252 4644 3884 4672
rect 1118 4564 1124 4616
rect 1176 4604 1182 4616
rect 1489 4607 1547 4613
rect 1489 4604 1501 4607
rect 1176 4576 1501 4604
rect 1176 4564 1182 4576
rect 1489 4573 1501 4576
rect 1535 4573 1547 4607
rect 1489 4567 1547 4573
rect 1946 4564 1952 4616
rect 2004 4604 2010 4616
rect 3252 4604 3280 4644
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 4157 4675 4215 4681
rect 4157 4641 4169 4675
rect 4203 4672 4215 4675
rect 4709 4675 4767 4681
rect 4203 4644 4568 4672
rect 4203 4641 4215 4644
rect 4157 4635 4215 4641
rect 2004 4576 3280 4604
rect 3329 4607 3387 4613
rect 2004 4564 2010 4576
rect 3329 4573 3341 4607
rect 3375 4573 3387 4607
rect 3329 4567 3387 4573
rect 3050 4496 3056 4548
rect 3108 4545 3114 4548
rect 3108 4536 3120 4545
rect 3344 4536 3372 4567
rect 3602 4564 3608 4616
rect 3660 4604 3666 4616
rect 3660 4576 3705 4604
rect 3660 4564 3666 4576
rect 3786 4564 3792 4616
rect 3844 4604 3850 4616
rect 4172 4604 4200 4635
rect 4430 4604 4436 4616
rect 3844 4576 4200 4604
rect 4391 4576 4436 4604
rect 3844 4564 3850 4576
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 4540 4604 4568 4644
rect 4709 4641 4721 4675
rect 4755 4672 4767 4675
rect 5074 4672 5080 4684
rect 4755 4644 5080 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 5074 4632 5080 4644
rect 5132 4672 5138 4684
rect 5460 4672 5488 4780
rect 5718 4700 5724 4752
rect 5776 4740 5782 4752
rect 6270 4740 6276 4752
rect 5776 4712 6276 4740
rect 5776 4700 5782 4712
rect 6270 4700 6276 4712
rect 6328 4700 6334 4752
rect 6380 4740 6408 4780
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 6880 4780 7420 4808
rect 6880 4768 6886 4780
rect 6380 4712 6960 4740
rect 5810 4672 5816 4684
rect 5132 4644 5488 4672
rect 5771 4644 5816 4672
rect 5132 4632 5138 4644
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 5960 4644 6005 4672
rect 5960 4632 5966 4644
rect 6178 4632 6184 4684
rect 6236 4632 6242 4684
rect 6454 4632 6460 4684
rect 6512 4672 6518 4684
rect 6932 4681 6960 4712
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6512 4644 6653 4672
rect 6512 4632 6518 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4641 6975 4675
rect 7392 4672 7420 4780
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 8941 4811 8999 4817
rect 8941 4808 8953 4811
rect 8352 4780 8953 4808
rect 8352 4768 8358 4780
rect 8941 4777 8953 4780
rect 8987 4777 8999 4811
rect 8941 4771 8999 4777
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9769 4811 9827 4817
rect 9769 4808 9781 4811
rect 9272 4780 9781 4808
rect 9272 4768 9278 4780
rect 9769 4777 9781 4780
rect 9815 4777 9827 4811
rect 11698 4808 11704 4820
rect 11659 4780 11704 4808
rect 9769 4771 9827 4777
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 12894 4808 12900 4820
rect 12855 4780 12900 4808
rect 12894 4768 12900 4780
rect 12952 4768 12958 4820
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 15286 4808 15292 4820
rect 13136 4780 15292 4808
rect 13136 4768 13142 4780
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 16758 4808 16764 4820
rect 16719 4780 16764 4808
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 18325 4811 18383 4817
rect 18325 4808 18337 4811
rect 17920 4780 18337 4808
rect 17920 4768 17926 4780
rect 18325 4777 18337 4780
rect 18371 4777 18383 4811
rect 18325 4771 18383 4777
rect 20625 4811 20683 4817
rect 20625 4777 20637 4811
rect 20671 4808 20683 4811
rect 21634 4808 21640 4820
rect 20671 4780 21640 4808
rect 20671 4777 20683 4780
rect 20625 4771 20683 4777
rect 21634 4768 21640 4780
rect 21692 4768 21698 4820
rect 8570 4700 8576 4752
rect 8628 4740 8634 4752
rect 8665 4743 8723 4749
rect 8665 4740 8677 4743
rect 8628 4712 8677 4740
rect 8628 4700 8634 4712
rect 8665 4709 8677 4712
rect 8711 4709 8723 4743
rect 8665 4703 8723 4709
rect 9306 4700 9312 4752
rect 9364 4740 9370 4752
rect 10778 4740 10784 4752
rect 9364 4712 10784 4740
rect 9364 4700 9370 4712
rect 8110 4672 8116 4684
rect 7392 4644 8116 4672
rect 6917 4635 6975 4641
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 9600 4681 9628 4712
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 10962 4700 10968 4752
rect 11020 4740 11026 4752
rect 12618 4740 12624 4752
rect 11020 4712 12624 4740
rect 11020 4700 11026 4712
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 13814 4740 13820 4752
rect 13648 4712 13820 4740
rect 9401 4675 9459 4681
rect 9401 4672 9413 4675
rect 9180 4644 9413 4672
rect 9180 4632 9186 4644
rect 9401 4641 9413 4644
rect 9447 4641 9459 4675
rect 9401 4635 9459 4641
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4641 9643 4675
rect 10226 4672 10232 4684
rect 10187 4644 10232 4672
rect 9585 4635 9643 4641
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 10410 4672 10416 4684
rect 10371 4644 10416 4672
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 11149 4675 11207 4681
rect 11149 4641 11161 4675
rect 11195 4672 11207 4675
rect 11238 4672 11244 4684
rect 11195 4644 11244 4672
rect 11195 4641 11207 4644
rect 11149 4635 11207 4641
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 13648 4681 13676 4712
rect 13814 4700 13820 4712
rect 13872 4740 13878 4752
rect 14734 4740 14740 4752
rect 13872 4712 14740 4740
rect 13872 4700 13878 4712
rect 14734 4700 14740 4712
rect 14792 4700 14798 4752
rect 12345 4675 12403 4681
rect 12345 4641 12357 4675
rect 12391 4672 12403 4675
rect 13633 4675 13691 4681
rect 13633 4672 13645 4675
rect 12391 4644 13645 4672
rect 12391 4641 12403 4644
rect 12345 4635 12403 4641
rect 13633 4641 13645 4644
rect 13679 4641 13691 4675
rect 13633 4635 13691 4641
rect 13722 4632 13728 4684
rect 13780 4672 13786 4684
rect 13909 4675 13967 4681
rect 13909 4672 13921 4675
rect 13780 4644 13921 4672
rect 13780 4632 13786 4644
rect 13909 4641 13921 4644
rect 13955 4672 13967 4675
rect 14366 4672 14372 4684
rect 13955 4644 14372 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 14366 4632 14372 4644
rect 14424 4632 14430 4684
rect 14645 4675 14703 4681
rect 14645 4641 14657 4675
rect 14691 4672 14703 4675
rect 16776 4672 16804 4768
rect 18233 4743 18291 4749
rect 18233 4709 18245 4743
rect 18279 4740 18291 4743
rect 18414 4740 18420 4752
rect 18279 4712 18420 4740
rect 18279 4709 18291 4712
rect 18233 4703 18291 4709
rect 18414 4700 18420 4712
rect 18472 4700 18478 4752
rect 19981 4743 20039 4749
rect 19981 4709 19993 4743
rect 20027 4709 20039 4743
rect 19981 4703 20039 4709
rect 18877 4675 18935 4681
rect 18877 4672 18889 4675
rect 14691 4644 15332 4672
rect 16776 4644 16988 4672
rect 14691 4641 14703 4644
rect 14645 4635 14703 4641
rect 5442 4604 5448 4616
rect 4540 4576 5448 4604
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 6086 4604 6092 4616
rect 5767 4576 6092 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 6196 4604 6224 4632
rect 6273 4607 6331 4613
rect 6273 4604 6285 4607
rect 6196 4576 6285 4604
rect 6273 4573 6285 4576
rect 6319 4573 6331 4607
rect 7742 4604 7748 4616
rect 6273 4567 6331 4573
rect 6472 4576 7748 4604
rect 4154 4536 4160 4548
rect 3108 4508 3153 4536
rect 3344 4508 4160 4536
rect 3108 4499 3120 4508
rect 3108 4496 3114 4499
rect 4154 4496 4160 4508
rect 4212 4536 4218 4548
rect 4614 4536 4620 4548
rect 4212 4508 4620 4536
rect 4212 4496 4218 4508
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 5810 4536 5816 4548
rect 5276 4508 5816 4536
rect 2038 4428 2044 4480
rect 2096 4468 2102 4480
rect 3602 4468 3608 4480
rect 2096 4440 3608 4468
rect 2096 4428 2102 4440
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 3970 4468 3976 4480
rect 3931 4440 3976 4468
rect 3970 4428 3976 4440
rect 4028 4428 4034 4480
rect 4246 4468 4252 4480
rect 4207 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4798 4468 4804 4480
rect 4759 4440 4804 4468
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 4890 4428 4896 4480
rect 4948 4468 4954 4480
rect 5276 4477 5304 4508
rect 5810 4496 5816 4508
rect 5868 4496 5874 4548
rect 6472 4536 6500 4576
rect 7742 4564 7748 4576
rect 7800 4604 7806 4616
rect 8481 4607 8539 4613
rect 8481 4604 8493 4607
rect 7800 4576 8493 4604
rect 7800 4564 7806 4576
rect 8481 4573 8493 4576
rect 8527 4573 8539 4607
rect 8481 4567 8539 4573
rect 8570 4564 8576 4616
rect 8628 4604 8634 4616
rect 9309 4607 9367 4613
rect 9309 4604 9321 4607
rect 8628 4576 9321 4604
rect 8628 4564 8634 4576
rect 9309 4573 9321 4576
rect 9355 4604 9367 4607
rect 9355 4576 9674 4604
rect 9355 4573 9367 4576
rect 9309 4567 9367 4573
rect 7282 4536 7288 4548
rect 5920 4508 6500 4536
rect 6748 4508 7288 4536
rect 5261 4471 5319 4477
rect 4948 4440 4993 4468
rect 4948 4428 4954 4440
rect 5261 4437 5273 4471
rect 5307 4437 5319 4471
rect 5261 4431 5319 4437
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 5920 4468 5948 4508
rect 5500 4440 5948 4468
rect 6365 4471 6423 4477
rect 5500 4428 5506 4440
rect 6365 4437 6377 4471
rect 6411 4468 6423 4471
rect 6748 4468 6776 4508
rect 7282 4496 7288 4508
rect 7340 4496 7346 4548
rect 7929 4539 7987 4545
rect 7929 4505 7941 4539
rect 7975 4536 7987 4539
rect 9646 4536 9674 4576
rect 9766 4564 9772 4616
rect 9824 4604 9830 4616
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 9824 4576 10149 4604
rect 9824 4564 9830 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10594 4604 10600 4616
rect 10555 4576 10600 4604
rect 10137 4567 10195 4573
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 11422 4564 11428 4616
rect 11480 4604 11486 4616
rect 11793 4607 11851 4613
rect 11793 4604 11805 4607
rect 11480 4576 11805 4604
rect 11480 4564 11486 4576
rect 11793 4573 11805 4576
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 12250 4564 12256 4616
rect 12308 4604 12314 4616
rect 14829 4607 14887 4613
rect 14829 4604 14841 4607
rect 12308 4576 14841 4604
rect 12308 4564 12314 4576
rect 14829 4573 14841 4576
rect 14875 4573 14887 4607
rect 14829 4567 14887 4573
rect 9950 4536 9956 4548
rect 7975 4508 8371 4536
rect 9646 4508 9956 4536
rect 7975 4505 7987 4508
rect 7929 4499 7987 4505
rect 6411 4440 6776 4468
rect 6411 4437 6423 4440
rect 6365 4431 6423 4437
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 7561 4471 7619 4477
rect 7561 4468 7573 4471
rect 7064 4440 7573 4468
rect 7064 4428 7070 4440
rect 7561 4437 7573 4440
rect 7607 4437 7619 4471
rect 7561 4431 7619 4437
rect 8018 4428 8024 4480
rect 8076 4468 8082 4480
rect 8343 4468 8371 4508
rect 9950 4496 9956 4508
rect 10008 4496 10014 4548
rect 10226 4496 10232 4548
rect 10284 4536 10290 4548
rect 11241 4539 11299 4545
rect 11241 4536 11253 4539
rect 10284 4508 11253 4536
rect 10284 4496 10290 4508
rect 11241 4505 11253 4508
rect 11287 4505 11299 4539
rect 11241 4499 11299 4505
rect 9214 4468 9220 4480
rect 8076 4440 8121 4468
rect 8343 4440 9220 4468
rect 8076 4428 8082 4440
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 10778 4468 10784 4480
rect 10739 4440 10784 4468
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11256 4468 11284 4499
rect 11330 4496 11336 4548
rect 11388 4536 11394 4548
rect 12342 4536 12348 4548
rect 11388 4508 12348 4536
rect 11388 4496 11394 4508
rect 12342 4496 12348 4508
rect 12400 4496 12406 4548
rect 12526 4536 12532 4548
rect 12487 4508 12532 4536
rect 12526 4496 12532 4508
rect 12584 4496 12590 4548
rect 13170 4496 13176 4548
rect 13228 4536 13234 4548
rect 13449 4539 13507 4545
rect 13449 4536 13461 4539
rect 13228 4508 13461 4536
rect 13228 4496 13234 4508
rect 13449 4505 13461 4508
rect 13495 4505 13507 4539
rect 13449 4499 13507 4505
rect 14458 4496 14464 4548
rect 14516 4536 14522 4548
rect 14737 4539 14795 4545
rect 14737 4536 14749 4539
rect 14516 4508 14749 4536
rect 14516 4496 14522 4508
rect 14737 4505 14749 4508
rect 14783 4536 14795 4539
rect 14918 4536 14924 4548
rect 14783 4508 14924 4536
rect 14783 4505 14795 4508
rect 14737 4499 14795 4505
rect 14918 4496 14924 4508
rect 14976 4496 14982 4548
rect 15304 4536 15332 4644
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 16850 4604 16856 4616
rect 15427 4576 16856 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 16960 4604 16988 4644
rect 17972 4644 18889 4672
rect 17972 4616 18000 4644
rect 18877 4641 18889 4644
rect 18923 4641 18935 4675
rect 18877 4635 18935 4641
rect 19429 4675 19487 4681
rect 19429 4641 19441 4675
rect 19475 4672 19487 4675
rect 19702 4672 19708 4684
rect 19475 4644 19708 4672
rect 19475 4641 19487 4644
rect 19429 4635 19487 4641
rect 19702 4632 19708 4644
rect 19760 4632 19766 4684
rect 17109 4607 17167 4613
rect 17109 4604 17121 4607
rect 16960 4576 17121 4604
rect 17109 4573 17121 4576
rect 17155 4604 17167 4607
rect 17954 4604 17960 4616
rect 17155 4576 17960 4604
rect 17155 4573 17167 4576
rect 17109 4567 17167 4573
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 18322 4564 18328 4616
rect 18380 4604 18386 4616
rect 18690 4604 18696 4616
rect 18380 4576 18696 4604
rect 18380 4564 18386 4576
rect 18690 4564 18696 4576
rect 18748 4564 18754 4616
rect 19518 4604 19524 4616
rect 19479 4576 19524 4604
rect 19518 4564 19524 4576
rect 19576 4564 19582 4616
rect 19996 4604 20024 4703
rect 20717 4675 20775 4681
rect 20717 4641 20729 4675
rect 20763 4672 20775 4675
rect 22554 4672 22560 4684
rect 20763 4644 22560 4672
rect 20763 4641 20775 4644
rect 20717 4635 20775 4641
rect 22554 4632 22560 4644
rect 22612 4632 22618 4684
rect 20073 4607 20131 4613
rect 20073 4604 20085 4607
rect 19996 4576 20085 4604
rect 20073 4573 20085 4576
rect 20119 4573 20131 4607
rect 20441 4607 20499 4613
rect 20441 4604 20453 4607
rect 20073 4567 20131 4573
rect 20272 4576 20453 4604
rect 15654 4545 15660 4548
rect 15648 4536 15660 4545
rect 15304 4508 15660 4536
rect 15648 4499 15660 4508
rect 15654 4496 15660 4499
rect 15712 4496 15718 4548
rect 18506 4496 18512 4548
rect 18564 4536 18570 4548
rect 19613 4539 19671 4545
rect 19613 4536 19625 4539
rect 18564 4508 19625 4536
rect 18564 4496 18570 4508
rect 19613 4505 19625 4508
rect 19659 4505 19671 4539
rect 19613 4499 19671 4505
rect 11882 4468 11888 4480
rect 11256 4440 11888 4468
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 11977 4471 12035 4477
rect 11977 4437 11989 4471
rect 12023 4468 12035 4471
rect 12250 4468 12256 4480
rect 12023 4440 12256 4468
rect 12023 4437 12035 4440
rect 11977 4431 12035 4437
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 12437 4471 12495 4477
rect 12437 4437 12449 4471
rect 12483 4468 12495 4471
rect 12618 4468 12624 4480
rect 12483 4440 12624 4468
rect 12483 4437 12495 4440
rect 12437 4431 12495 4437
rect 12618 4428 12624 4440
rect 12676 4428 12682 4480
rect 12989 4471 13047 4477
rect 12989 4437 13001 4471
rect 13035 4468 13047 4471
rect 13078 4468 13084 4480
rect 13035 4440 13084 4468
rect 13035 4437 13047 4440
rect 12989 4431 13047 4437
rect 13078 4428 13084 4440
rect 13136 4428 13142 4480
rect 13354 4468 13360 4480
rect 13315 4440 13360 4468
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 14366 4468 14372 4480
rect 14327 4440 14372 4468
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 15197 4471 15255 4477
rect 15197 4437 15209 4471
rect 15243 4468 15255 4471
rect 16942 4468 16948 4480
rect 15243 4440 16948 4468
rect 15243 4437 15255 4440
rect 15197 4431 15255 4437
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 18690 4468 18696 4480
rect 18651 4440 18696 4468
rect 18690 4428 18696 4440
rect 18748 4428 18754 4480
rect 18782 4428 18788 4480
rect 18840 4468 18846 4480
rect 20272 4477 20300 4576
rect 20441 4573 20453 4576
rect 20487 4573 20499 4607
rect 20441 4567 20499 4573
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4604 21051 4607
rect 21358 4604 21364 4616
rect 21039 4576 21364 4604
rect 21039 4573 21051 4576
rect 20993 4567 21051 4573
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 20257 4471 20315 4477
rect 18840 4440 18885 4468
rect 18840 4428 18846 4440
rect 20257 4437 20269 4471
rect 20303 4437 20315 4471
rect 20257 4431 20315 4437
rect 20714 4428 20720 4480
rect 20772 4468 20778 4480
rect 21266 4468 21272 4480
rect 20772 4440 21272 4468
rect 20772 4428 20778 4440
rect 21266 4428 21272 4440
rect 21324 4428 21330 4480
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 1854 4264 1860 4276
rect 1815 4236 1860 4264
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 2317 4267 2375 4273
rect 2317 4233 2329 4267
rect 2363 4264 2375 4267
rect 2685 4267 2743 4273
rect 2363 4236 2636 4264
rect 2363 4233 2375 4236
rect 2317 4227 2375 4233
rect 2608 4196 2636 4236
rect 2685 4233 2697 4267
rect 2731 4264 2743 4267
rect 2774 4264 2780 4276
rect 2731 4236 2780 4264
rect 2731 4233 2743 4236
rect 2685 4227 2743 4233
rect 2774 4224 2780 4236
rect 2832 4224 2838 4276
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3237 4267 3295 4273
rect 3237 4264 3249 4267
rect 3108 4236 3249 4264
rect 3108 4224 3114 4236
rect 3237 4233 3249 4236
rect 3283 4264 3295 4267
rect 3878 4264 3884 4276
rect 3283 4236 3884 4264
rect 3283 4233 3295 4236
rect 3237 4227 3295 4233
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 5534 4264 5540 4276
rect 4764 4236 5540 4264
rect 4764 4224 4770 4236
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 5902 4264 5908 4276
rect 5736 4236 5908 4264
rect 2608 4168 2820 4196
rect 2792 4137 2820 4168
rect 3142 4156 3148 4208
rect 3200 4196 3206 4208
rect 5736 4196 5764 4236
rect 5902 4224 5908 4236
rect 5960 4224 5966 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 9125 4267 9183 4273
rect 9125 4264 9137 4267
rect 8352 4236 9137 4264
rect 8352 4224 8358 4236
rect 9125 4233 9137 4236
rect 9171 4233 9183 4267
rect 9490 4264 9496 4276
rect 9451 4236 9496 4264
rect 9125 4227 9183 4233
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 11333 4267 11391 4273
rect 11333 4233 11345 4267
rect 11379 4264 11391 4267
rect 11698 4264 11704 4276
rect 11379 4236 11704 4264
rect 11379 4233 11391 4236
rect 11333 4227 11391 4233
rect 11698 4224 11704 4236
rect 11756 4224 11762 4276
rect 11790 4224 11796 4276
rect 11848 4264 11854 4276
rect 12158 4264 12164 4276
rect 11848 4236 12164 4264
rect 11848 4224 11854 4236
rect 12158 4224 12164 4236
rect 12216 4264 12222 4276
rect 12618 4264 12624 4276
rect 12216 4236 12624 4264
rect 12216 4224 12222 4236
rect 12618 4224 12624 4236
rect 12676 4224 12682 4276
rect 12986 4224 12992 4276
rect 13044 4264 13050 4276
rect 13173 4267 13231 4273
rect 13173 4264 13185 4267
rect 13044 4236 13185 4264
rect 13044 4224 13050 4236
rect 13173 4233 13185 4236
rect 13219 4264 13231 4267
rect 13722 4264 13728 4276
rect 13219 4236 13728 4264
rect 13219 4233 13231 4236
rect 13173 4227 13231 4233
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 14829 4267 14887 4273
rect 14829 4233 14841 4267
rect 14875 4264 14887 4267
rect 15289 4267 15347 4273
rect 15289 4264 15301 4267
rect 14875 4236 15301 4264
rect 14875 4233 14887 4236
rect 14829 4227 14887 4233
rect 15289 4233 15301 4236
rect 15335 4233 15347 4267
rect 15289 4227 15347 4233
rect 16298 4224 16304 4276
rect 16356 4264 16362 4276
rect 16850 4264 16856 4276
rect 16356 4236 16856 4264
rect 16356 4224 16362 4236
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 16942 4224 16948 4276
rect 17000 4264 17006 4276
rect 17000 4236 17448 4264
rect 17000 4224 17006 4236
rect 3200 4168 5764 4196
rect 5813 4199 5871 4205
rect 3200 4156 3206 4168
rect 5813 4165 5825 4199
rect 5859 4196 5871 4199
rect 6270 4196 6276 4208
rect 5859 4168 6276 4196
rect 5859 4165 5871 4168
rect 5813 4159 5871 4165
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 6454 4156 6460 4208
rect 6512 4196 6518 4208
rect 6641 4199 6699 4205
rect 6641 4196 6653 4199
rect 6512 4168 6653 4196
rect 6512 4156 6518 4168
rect 6641 4165 6653 4168
rect 6687 4165 6699 4199
rect 6641 4159 6699 4165
rect 6825 4199 6883 4205
rect 6825 4165 6837 4199
rect 6871 4196 6883 4199
rect 7098 4196 7104 4208
rect 6871 4168 7104 4196
rect 6871 4165 6883 4168
rect 6825 4159 6883 4165
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 9677 4199 9735 4205
rect 9048 4168 9260 4196
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4128 2007 4131
rect 2777 4131 2835 4137
rect 1995 4100 2452 4128
rect 1995 4097 2007 4100
rect 1949 4091 2007 4097
rect 1670 4060 1676 4072
rect 1631 4032 1676 4060
rect 1670 4020 1676 4032
rect 1728 4020 1734 4072
rect 2424 3992 2452 4100
rect 2777 4097 2789 4131
rect 2823 4097 2835 4131
rect 2777 4091 2835 4097
rect 4361 4131 4419 4137
rect 4361 4097 4373 4131
rect 4407 4128 4419 4131
rect 4890 4128 4896 4140
rect 4407 4100 4896 4128
rect 4407 4097 4419 4100
rect 4361 4091 4419 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5166 4128 5172 4140
rect 5127 4100 5172 4128
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 7184 4131 7242 4137
rect 5592 4100 6500 4128
rect 5592 4088 5598 4100
rect 2593 4063 2651 4069
rect 2593 4029 2605 4063
rect 2639 4060 2651 4063
rect 2958 4060 2964 4072
rect 2639 4032 2964 4060
rect 2639 4029 2651 4032
rect 2593 4023 2651 4029
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 4614 4060 4620 4072
rect 4575 4032 4620 4060
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 4706 4020 4712 4072
rect 4764 4060 4770 4072
rect 5442 4060 5448 4072
rect 4764 4032 4809 4060
rect 5276 4032 5448 4060
rect 4764 4020 4770 4032
rect 2866 3992 2872 4004
rect 2424 3964 2872 3992
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 3145 3995 3203 4001
rect 3145 3961 3157 3995
rect 3191 3992 3203 3995
rect 3326 3992 3332 4004
rect 3191 3964 3332 3992
rect 3191 3961 3203 3964
rect 3145 3955 3203 3961
rect 3326 3952 3332 3964
rect 3384 3952 3390 4004
rect 5276 3992 5304 4032
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5905 4063 5963 4069
rect 5905 4029 5917 4063
rect 5951 4060 5963 4063
rect 5994 4060 6000 4072
rect 5951 4032 6000 4060
rect 5951 4029 5963 4032
rect 5905 4023 5963 4029
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4060 6147 4063
rect 6178 4060 6184 4072
rect 6135 4032 6184 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 6362 4060 6368 4072
rect 6323 4032 6368 4060
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 6472 4060 6500 4100
rect 7184 4097 7196 4131
rect 7230 4128 7242 4131
rect 8110 4128 8116 4140
rect 7230 4100 8116 4128
rect 7230 4097 7242 4100
rect 7184 4091 7242 4097
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8478 4128 8484 4140
rect 8439 4100 8484 4128
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 9048 4128 9076 4168
rect 8956 4100 9076 4128
rect 8956 4069 8984 4100
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 6472 4032 6929 4060
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 8941 4063 8999 4069
rect 8941 4029 8953 4063
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 9033 4063 9091 4069
rect 9033 4029 9045 4063
rect 9079 4029 9091 4063
rect 9232 4060 9260 4168
rect 9677 4165 9689 4199
rect 9723 4165 9735 4199
rect 13538 4196 13544 4208
rect 9677 4159 9735 4165
rect 12728 4168 13544 4196
rect 9306 4088 9312 4140
rect 9364 4128 9370 4140
rect 9692 4128 9720 4159
rect 10209 4131 10267 4137
rect 10209 4128 10221 4131
rect 9364 4100 9720 4128
rect 9784 4100 10221 4128
rect 9364 4088 9370 4100
rect 9582 4060 9588 4072
rect 9232 4032 9588 4060
rect 9033 4023 9091 4029
rect 4724 3964 5304 3992
rect 5353 3995 5411 4001
rect 1489 3927 1547 3933
rect 1489 3893 1501 3927
rect 1535 3924 1547 3927
rect 4724 3924 4752 3964
rect 5353 3961 5365 3995
rect 5399 3992 5411 3995
rect 5399 3964 6868 3992
rect 5399 3961 5411 3964
rect 5353 3955 5411 3961
rect 1535 3896 4752 3924
rect 1535 3893 1547 3896
rect 1489 3887 1547 3893
rect 4798 3884 4804 3936
rect 4856 3924 4862 3936
rect 4985 3927 5043 3933
rect 4985 3924 4997 3927
rect 4856 3896 4997 3924
rect 4856 3884 4862 3896
rect 4985 3893 4997 3896
rect 5031 3893 5043 3927
rect 4985 3887 5043 3893
rect 5445 3927 5503 3933
rect 5445 3893 5457 3927
rect 5491 3924 5503 3927
rect 5718 3924 5724 3936
rect 5491 3896 5724 3924
rect 5491 3893 5503 3896
rect 5445 3887 5503 3893
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6840 3924 6868 3964
rect 8036 3964 8708 3992
rect 8036 3924 8064 3964
rect 6840 3896 8064 3924
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8297 3927 8355 3933
rect 8297 3924 8309 3927
rect 8168 3896 8309 3924
rect 8168 3884 8174 3896
rect 8297 3893 8309 3896
rect 8343 3893 8355 3927
rect 8570 3924 8576 3936
rect 8531 3896 8576 3924
rect 8297 3887 8355 3893
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 8680 3924 8708 3964
rect 8754 3952 8760 4004
rect 8812 3992 8818 4004
rect 9048 3992 9076 4023
rect 9582 4020 9588 4032
rect 9640 4060 9646 4072
rect 9784 4060 9812 4100
rect 10209 4097 10221 4100
rect 10255 4097 10267 4131
rect 10209 4091 10267 4097
rect 10778 4088 10784 4140
rect 10836 4128 10842 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 10836 4100 11529 4128
rect 10836 4088 10842 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 12161 4131 12219 4137
rect 12161 4128 12173 4131
rect 11793 4091 11851 4097
rect 11992 4100 12173 4128
rect 9950 4060 9956 4072
rect 9640 4032 9812 4060
rect 9911 4032 9956 4060
rect 9640 4020 9646 4032
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 10962 4020 10968 4072
rect 11020 4060 11026 4072
rect 11808 4060 11836 4091
rect 11020 4032 11836 4060
rect 11020 4020 11026 4032
rect 11992 4001 12020 4100
rect 12161 4097 12173 4100
rect 12207 4097 12219 4131
rect 12618 4128 12624 4140
rect 12579 4100 12624 4128
rect 12161 4091 12219 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 12728 4060 12756 4168
rect 13538 4156 13544 4168
rect 13596 4156 13602 4208
rect 15657 4199 15715 4205
rect 15657 4165 15669 4199
rect 15703 4196 15715 4199
rect 16114 4196 16120 4208
rect 15703 4168 16120 4196
rect 15703 4165 15715 4168
rect 15657 4159 15715 4165
rect 16114 4156 16120 4168
rect 16172 4196 16178 4208
rect 16172 4168 17356 4196
rect 16172 4156 16178 4168
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 12860 4100 12940 4128
rect 12860 4088 12866 4100
rect 12912 4069 12940 4100
rect 13078 4088 13084 4140
rect 13136 4128 13142 4140
rect 13136 4100 13181 4128
rect 13136 4088 13142 4100
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13872 4100 14013 4128
rect 13872 4088 13878 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 12084 4032 12756 4060
rect 12897 4063 12955 4069
rect 11977 3995 12035 4001
rect 8812 3964 9076 3992
rect 11532 3964 11928 3992
rect 8812 3952 8818 3964
rect 9674 3924 9680 3936
rect 8680 3896 9680 3924
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 9769 3927 9827 3933
rect 9769 3893 9781 3927
rect 9815 3924 9827 3927
rect 11532 3924 11560 3964
rect 11698 3924 11704 3936
rect 9815 3896 11560 3924
rect 11659 3896 11704 3924
rect 9815 3893 9827 3896
rect 9769 3887 9827 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 11900 3924 11928 3964
rect 11977 3961 11989 3995
rect 12023 3961 12035 3995
rect 11977 3955 12035 3961
rect 12084 3924 12112 4032
rect 12897 4029 12909 4063
rect 12943 4029 12955 4063
rect 14093 4063 14151 4069
rect 14093 4060 14105 4063
rect 12897 4023 12955 4029
rect 13556 4032 14105 4060
rect 12526 3952 12532 4004
rect 12584 3992 12590 4004
rect 13446 3992 13452 4004
rect 12584 3964 13452 3992
rect 12584 3952 12590 3964
rect 13446 3952 13452 3964
rect 13504 3952 13510 4004
rect 13556 4001 13584 4032
rect 14093 4029 14105 4032
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4029 14243 4063
rect 14918 4060 14924 4072
rect 14879 4032 14924 4060
rect 14185 4023 14243 4029
rect 13541 3995 13599 4001
rect 13541 3961 13553 3995
rect 13587 3961 13599 3995
rect 13541 3955 13599 3961
rect 13722 3952 13728 4004
rect 13780 3992 13786 4004
rect 14200 3992 14228 4023
rect 14918 4020 14924 4032
rect 14976 4020 14982 4072
rect 15010 4020 15016 4072
rect 15068 4060 15074 4072
rect 15068 4032 15113 4060
rect 15068 4020 15074 4032
rect 15562 4020 15568 4072
rect 15620 4060 15626 4072
rect 15749 4063 15807 4069
rect 15749 4060 15761 4063
rect 15620 4032 15761 4060
rect 15620 4020 15626 4032
rect 15749 4029 15761 4032
rect 15795 4029 15807 4063
rect 15930 4060 15936 4072
rect 15891 4032 15936 4060
rect 15749 4023 15807 4029
rect 15930 4020 15936 4032
rect 15988 4060 15994 4072
rect 16316 4060 16344 4091
rect 16390 4088 16396 4140
rect 16448 4128 16454 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16448 4100 16681 4128
rect 16448 4088 16454 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 16942 4088 16948 4140
rect 17000 4128 17006 4140
rect 17037 4131 17095 4137
rect 17037 4128 17049 4131
rect 17000 4100 17049 4128
rect 17000 4088 17006 4100
rect 17037 4097 17049 4100
rect 17083 4128 17095 4131
rect 17218 4128 17224 4140
rect 17083 4100 17224 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 15988 4032 16344 4060
rect 15988 4020 15994 4032
rect 13780 3964 14228 3992
rect 13780 3952 13786 3964
rect 15654 3952 15660 4004
rect 15712 3992 15718 4004
rect 16408 3992 16436 4088
rect 16942 3992 16948 4004
rect 15712 3964 16948 3992
rect 15712 3952 15718 3964
rect 16942 3952 16948 3964
rect 17000 3952 17006 4004
rect 17328 4001 17356 4168
rect 17420 4128 17448 4236
rect 17586 4224 17592 4276
rect 17644 4264 17650 4276
rect 17773 4267 17831 4273
rect 17773 4264 17785 4267
rect 17644 4236 17785 4264
rect 17644 4224 17650 4236
rect 17773 4233 17785 4236
rect 17819 4233 17831 4267
rect 17773 4227 17831 4233
rect 18138 4224 18144 4276
rect 18196 4264 18202 4276
rect 20438 4264 20444 4276
rect 18196 4236 20444 4264
rect 18196 4224 18202 4236
rect 20438 4224 20444 4236
rect 20496 4224 20502 4276
rect 20533 4267 20591 4273
rect 20533 4233 20545 4267
rect 20579 4233 20591 4267
rect 20533 4227 20591 4233
rect 18601 4199 18659 4205
rect 18601 4165 18613 4199
rect 18647 4196 18659 4199
rect 19061 4199 19119 4205
rect 19061 4196 19073 4199
rect 18647 4168 19073 4196
rect 18647 4165 18659 4168
rect 18601 4159 18659 4165
rect 19061 4165 19073 4168
rect 19107 4165 19119 4199
rect 20548 4196 20576 4227
rect 20990 4196 20996 4208
rect 19061 4159 19119 4165
rect 19628 4168 20208 4196
rect 20548 4168 20996 4196
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 17420 4100 17693 4128
rect 17681 4097 17693 4100
rect 17727 4097 17739 4131
rect 17681 4091 17739 4097
rect 17972 4100 18828 4128
rect 17972 4072 18000 4100
rect 17589 4063 17647 4069
rect 17589 4029 17601 4063
rect 17635 4060 17647 4063
rect 17954 4060 17960 4072
rect 17635 4032 17960 4060
rect 17635 4029 17647 4032
rect 17589 4023 17647 4029
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 18800 4069 18828 4100
rect 18966 4088 18972 4140
rect 19024 4128 19030 4140
rect 19628 4128 19656 4168
rect 19794 4128 19800 4140
rect 19024 4100 19656 4128
rect 19755 4100 19800 4128
rect 19024 4088 19030 4100
rect 19794 4088 19800 4100
rect 19852 4088 19858 4140
rect 19978 4088 19984 4140
rect 20036 4128 20042 4140
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 20036 4100 20085 4128
rect 20036 4088 20042 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20180 4128 20208 4168
rect 20990 4156 20996 4168
rect 21048 4156 21054 4208
rect 21082 4156 21088 4208
rect 21140 4196 21146 4208
rect 21450 4196 21456 4208
rect 21140 4168 21185 4196
rect 21411 4168 21456 4196
rect 21140 4156 21146 4168
rect 21450 4156 21456 4168
rect 21508 4156 21514 4208
rect 22002 4156 22008 4208
rect 22060 4196 22066 4208
rect 22554 4196 22560 4208
rect 22060 4168 22560 4196
rect 22060 4156 22066 4168
rect 22554 4156 22560 4168
rect 22612 4156 22618 4208
rect 20349 4131 20407 4137
rect 20349 4128 20361 4131
rect 20180 4100 20361 4128
rect 20073 4091 20131 4097
rect 20349 4097 20361 4100
rect 20395 4097 20407 4131
rect 20714 4128 20720 4140
rect 20349 4091 20407 4097
rect 20456 4100 20720 4128
rect 18693 4063 18751 4069
rect 18693 4029 18705 4063
rect 18739 4029 18751 4063
rect 18693 4023 18751 4029
rect 18785 4063 18843 4069
rect 18785 4029 18797 4063
rect 18831 4029 18843 4063
rect 18785 4023 18843 4029
rect 17313 3995 17371 4001
rect 17313 3961 17325 3995
rect 17359 3992 17371 3995
rect 17770 3992 17776 4004
rect 17359 3964 17776 3992
rect 17359 3961 17371 3964
rect 17313 3955 17371 3961
rect 17770 3952 17776 3964
rect 17828 3952 17834 4004
rect 18046 3952 18052 4004
rect 18104 3992 18110 4004
rect 18141 3995 18199 4001
rect 18141 3992 18153 3995
rect 18104 3964 18153 3992
rect 18104 3952 18110 3964
rect 18141 3961 18153 3964
rect 18187 3961 18199 3995
rect 18141 3955 18199 3961
rect 18230 3952 18236 4004
rect 18288 3992 18294 4004
rect 18288 3964 18333 3992
rect 18288 3952 18294 3964
rect 12342 3924 12348 3936
rect 11900 3896 12112 3924
rect 12303 3896 12348 3924
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12492 3896 12537 3924
rect 12492 3884 12498 3896
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 13633 3927 13691 3933
rect 13633 3924 13645 3927
rect 12952 3896 13645 3924
rect 12952 3884 12958 3896
rect 13633 3893 13645 3896
rect 13679 3893 13691 3927
rect 13633 3887 13691 3893
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3924 14519 3927
rect 14550 3924 14556 3936
rect 14507 3896 14556 3924
rect 14507 3893 14519 3896
rect 14461 3887 14519 3893
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 16209 3927 16267 3933
rect 16209 3924 16221 3927
rect 14792 3896 16221 3924
rect 14792 3884 14798 3896
rect 16209 3893 16221 3896
rect 16255 3893 16267 3927
rect 16209 3887 16267 3893
rect 17218 3884 17224 3936
rect 17276 3924 17282 3936
rect 18708 3924 18736 4023
rect 19613 3995 19671 4001
rect 19613 3961 19625 3995
rect 19659 3992 19671 3995
rect 19702 3992 19708 4004
rect 19659 3964 19708 3992
rect 19659 3961 19671 3964
rect 19613 3955 19671 3961
rect 19702 3952 19708 3964
rect 19760 3952 19766 4004
rect 19981 3995 20039 4001
rect 19981 3961 19993 3995
rect 20027 3992 20039 3995
rect 20162 3992 20168 4004
rect 20027 3964 20168 3992
rect 20027 3961 20039 3964
rect 19981 3955 20039 3961
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 20257 3995 20315 4001
rect 20257 3961 20269 3995
rect 20303 3992 20315 3995
rect 20456 3992 20484 4100
rect 20714 4088 20720 4100
rect 20772 4088 20778 4140
rect 20809 4131 20867 4137
rect 20809 4097 20821 4131
rect 20855 4128 20867 4131
rect 20855 4100 21036 4128
rect 20855 4097 20867 4100
rect 20809 4091 20867 4097
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 20901 4063 20959 4069
rect 20901 4060 20913 4063
rect 20588 4032 20913 4060
rect 20588 4020 20594 4032
rect 20901 4029 20913 4032
rect 20947 4029 20959 4063
rect 21008 4060 21036 4100
rect 22002 4060 22008 4072
rect 21008 4032 22008 4060
rect 20901 4023 20959 4029
rect 22002 4020 22008 4032
rect 22060 4020 22066 4072
rect 22186 3992 22192 4004
rect 20303 3964 20484 3992
rect 21284 3964 22192 3992
rect 20303 3961 20315 3964
rect 20257 3955 20315 3961
rect 19426 3924 19432 3936
rect 17276 3896 18736 3924
rect 19339 3896 19432 3924
rect 17276 3884 17282 3896
rect 19426 3884 19432 3896
rect 19484 3924 19490 3936
rect 20438 3924 20444 3936
rect 19484 3896 20444 3924
rect 19484 3884 19490 3896
rect 20438 3884 20444 3896
rect 20496 3884 20502 3936
rect 20625 3927 20683 3933
rect 20625 3893 20637 3927
rect 20671 3924 20683 3927
rect 21284 3924 21312 3964
rect 22186 3952 22192 3964
rect 22244 3952 22250 4004
rect 20671 3896 21312 3924
rect 20671 3893 20683 3896
rect 20625 3887 20683 3893
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 21416 3896 21461 3924
rect 21416 3884 21422 3896
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 1949 3723 2007 3729
rect 1949 3689 1961 3723
rect 1995 3720 2007 3723
rect 2038 3720 2044 3732
rect 1995 3692 2044 3720
rect 1995 3689 2007 3692
rect 1949 3683 2007 3689
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 3881 3723 3939 3729
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 5534 3720 5540 3732
rect 3927 3692 5540 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 5902 3680 5908 3732
rect 5960 3720 5966 3732
rect 6181 3723 6239 3729
rect 6181 3720 6193 3723
rect 5960 3692 6193 3720
rect 5960 3680 5966 3692
rect 6181 3689 6193 3692
rect 6227 3689 6239 3723
rect 6181 3683 6239 3689
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 8294 3720 8300 3732
rect 7147 3692 8300 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 8662 3680 8668 3732
rect 8720 3720 8726 3732
rect 8757 3723 8815 3729
rect 8757 3720 8769 3723
rect 8720 3692 8769 3720
rect 8720 3680 8726 3692
rect 8757 3689 8769 3692
rect 8803 3689 8815 3723
rect 10134 3720 10140 3732
rect 10095 3692 10140 3720
rect 8757 3683 8815 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10686 3720 10692 3732
rect 10336 3692 10692 3720
rect 1670 3652 1676 3664
rect 1583 3624 1676 3652
rect 1670 3612 1676 3624
rect 1728 3652 1734 3664
rect 2314 3652 2320 3664
rect 1728 3624 2320 3652
rect 1728 3612 1734 3624
rect 2314 3612 2320 3624
rect 2372 3612 2378 3664
rect 4706 3652 4712 3664
rect 2424 3624 4712 3652
rect 1854 3544 1860 3596
rect 1912 3584 1918 3596
rect 2424 3584 2452 3624
rect 4706 3612 4712 3624
rect 4764 3612 4770 3664
rect 8110 3652 8116 3664
rect 6472 3624 8116 3652
rect 2590 3584 2596 3596
rect 1912 3556 2452 3584
rect 2551 3556 2596 3584
rect 1912 3544 1918 3556
rect 2590 3544 2596 3556
rect 2648 3544 2654 3596
rect 3050 3544 3056 3596
rect 3108 3584 3114 3596
rect 3421 3587 3479 3593
rect 3421 3584 3433 3587
rect 3108 3556 3433 3584
rect 3108 3544 3114 3556
rect 3421 3553 3433 3556
rect 3467 3553 3479 3587
rect 3421 3547 3479 3553
rect 3510 3544 3516 3596
rect 3568 3584 3574 3596
rect 6472 3593 6500 3624
rect 8110 3612 8116 3624
rect 8168 3652 8174 3664
rect 9306 3652 9312 3664
rect 8168 3624 8248 3652
rect 8168 3612 8174 3624
rect 4157 3587 4215 3593
rect 4157 3584 4169 3587
rect 3568 3556 4169 3584
rect 3568 3544 3574 3556
rect 4157 3553 4169 3556
rect 4203 3584 4215 3587
rect 6457 3587 6515 3593
rect 4203 3556 4936 3584
rect 4203 3553 4215 3556
rect 4157 3547 4215 3553
rect 1486 3516 1492 3528
rect 1447 3488 1492 3516
rect 1486 3476 1492 3488
rect 1544 3476 1550 3528
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3516 1823 3519
rect 2409 3519 2467 3525
rect 1811 3488 2084 3516
rect 1811 3485 1823 3488
rect 1765 3479 1823 3485
rect 2056 3389 2084 3488
rect 2409 3485 2421 3519
rect 2455 3516 2467 3519
rect 2498 3516 2504 3528
rect 2455 3488 2504 3516
rect 2455 3485 2467 3488
rect 2409 3479 2467 3485
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 4614 3516 4620 3528
rect 4295 3488 4620 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3485 4859 3519
rect 4908 3516 4936 3556
rect 6457 3553 6469 3587
rect 6503 3553 6515 3587
rect 6457 3547 6515 3553
rect 6641 3587 6699 3593
rect 6641 3553 6653 3587
rect 6687 3584 6699 3587
rect 7006 3584 7012 3596
rect 6687 3556 7012 3584
rect 6687 3553 6699 3556
rect 6641 3547 6699 3553
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 8220 3593 8248 3624
rect 8680 3624 9312 3652
rect 8680 3596 8708 3624
rect 9306 3612 9312 3624
rect 9364 3612 9370 3664
rect 10042 3612 10048 3664
rect 10100 3652 10106 3664
rect 10336 3652 10364 3692
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 11238 3680 11244 3732
rect 11296 3720 11302 3732
rect 11701 3723 11759 3729
rect 11701 3720 11713 3723
rect 11296 3692 11713 3720
rect 11296 3680 11302 3692
rect 11701 3689 11713 3692
rect 11747 3689 11759 3723
rect 11882 3720 11888 3732
rect 11843 3692 11888 3720
rect 11701 3683 11759 3689
rect 11882 3680 11888 3692
rect 11940 3680 11946 3732
rect 12342 3680 12348 3732
rect 12400 3720 12406 3732
rect 13170 3720 13176 3732
rect 12400 3692 13176 3720
rect 12400 3680 12406 3692
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 14458 3720 14464 3732
rect 13320 3692 14464 3720
rect 13320 3680 13326 3692
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 14918 3680 14924 3732
rect 14976 3720 14982 3732
rect 15105 3723 15163 3729
rect 15105 3720 15117 3723
rect 14976 3692 15117 3720
rect 14976 3680 14982 3692
rect 15105 3689 15117 3692
rect 15151 3689 15163 3723
rect 16485 3723 16543 3729
rect 16485 3720 16497 3723
rect 15105 3683 15163 3689
rect 15212 3692 16497 3720
rect 10100 3624 10364 3652
rect 10100 3612 10106 3624
rect 13906 3612 13912 3664
rect 13964 3652 13970 3664
rect 15212 3652 15240 3692
rect 16485 3689 16497 3692
rect 16531 3689 16543 3723
rect 16850 3720 16856 3732
rect 16811 3692 16856 3720
rect 16485 3683 16543 3689
rect 16850 3680 16856 3692
rect 16908 3680 16914 3732
rect 18141 3723 18199 3729
rect 18141 3689 18153 3723
rect 18187 3720 18199 3723
rect 18690 3720 18696 3732
rect 18187 3692 18696 3720
rect 18187 3689 18199 3692
rect 18141 3683 18199 3689
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 18782 3680 18788 3732
rect 18840 3720 18846 3732
rect 18969 3723 19027 3729
rect 18969 3720 18981 3723
rect 18840 3692 18981 3720
rect 18840 3680 18846 3692
rect 18969 3689 18981 3692
rect 19015 3689 19027 3723
rect 18969 3683 19027 3689
rect 19886 3680 19892 3732
rect 19944 3720 19950 3732
rect 19981 3723 20039 3729
rect 19981 3720 19993 3723
rect 19944 3692 19993 3720
rect 19944 3680 19950 3692
rect 19981 3689 19993 3692
rect 20027 3689 20039 3723
rect 19981 3683 20039 3689
rect 20162 3680 20168 3732
rect 20220 3720 20226 3732
rect 20530 3720 20536 3732
rect 20220 3692 20536 3720
rect 20220 3680 20226 3692
rect 20530 3680 20536 3692
rect 20588 3680 20594 3732
rect 20714 3680 20720 3732
rect 20772 3720 20778 3732
rect 22646 3720 22652 3732
rect 20772 3692 22652 3720
rect 20772 3680 20778 3692
rect 22646 3680 22652 3692
rect 22704 3680 22710 3732
rect 15930 3652 15936 3664
rect 13964 3624 15240 3652
rect 15764 3624 15936 3652
rect 13964 3612 13970 3624
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3553 7343 3587
rect 7285 3547 7343 3553
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3553 8263 3587
rect 8205 3547 8263 3553
rect 8297 3587 8355 3593
rect 8297 3553 8309 3587
rect 8343 3584 8355 3587
rect 8386 3584 8392 3596
rect 8343 3556 8392 3584
rect 8343 3553 8355 3556
rect 8297 3547 8355 3553
rect 5074 3525 5080 3528
rect 5068 3516 5080 3525
rect 4908 3488 5080 3516
rect 4801 3479 4859 3485
rect 5068 3479 5080 3488
rect 3878 3408 3884 3460
rect 3936 3448 3942 3460
rect 4816 3448 4844 3479
rect 5074 3476 5080 3479
rect 5132 3476 5138 3528
rect 5442 3476 5448 3528
rect 5500 3476 5506 3528
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6604 3488 6745 3516
rect 6604 3476 6610 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 6822 3476 6828 3528
rect 6880 3516 6886 3528
rect 7300 3516 7328 3547
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 8662 3544 8668 3596
rect 8720 3544 8726 3596
rect 12526 3584 12532 3596
rect 11348 3556 12532 3584
rect 6880 3488 7328 3516
rect 7469 3519 7527 3525
rect 6880 3476 6886 3488
rect 7469 3485 7481 3519
rect 7515 3516 7527 3519
rect 8754 3516 8760 3528
rect 7515 3512 8156 3516
rect 8220 3512 8760 3516
rect 7515 3488 8760 3512
rect 7515 3485 7527 3488
rect 7469 3479 7527 3485
rect 8128 3484 8248 3488
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 5460 3448 5488 3476
rect 5994 3448 6000 3460
rect 3936 3420 6000 3448
rect 3936 3408 3942 3420
rect 5994 3408 6000 3420
rect 6052 3408 6058 3460
rect 6178 3408 6184 3460
rect 6236 3448 6242 3460
rect 7006 3448 7012 3460
rect 6236 3420 7012 3448
rect 6236 3408 6242 3420
rect 7006 3408 7012 3420
rect 7064 3408 7070 3460
rect 8389 3451 8447 3457
rect 8389 3448 8401 3451
rect 7944 3420 8401 3448
rect 2041 3383 2099 3389
rect 2041 3349 2053 3383
rect 2087 3349 2099 3383
rect 2041 3343 2099 3349
rect 2501 3383 2559 3389
rect 2501 3349 2513 3383
rect 2547 3380 2559 3383
rect 2869 3383 2927 3389
rect 2869 3380 2881 3383
rect 2547 3352 2881 3380
rect 2547 3349 2559 3352
rect 2501 3343 2559 3349
rect 2869 3349 2881 3352
rect 2915 3349 2927 3383
rect 3234 3380 3240 3392
rect 3195 3352 3240 3380
rect 2869 3343 2927 3349
rect 3234 3340 3240 3352
rect 3292 3340 3298 3392
rect 3326 3340 3332 3392
rect 3384 3380 3390 3392
rect 4338 3380 4344 3392
rect 3384 3352 3429 3380
rect 4299 3352 4344 3380
rect 3384 3340 3390 3352
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 4709 3383 4767 3389
rect 4709 3349 4721 3383
rect 4755 3380 4767 3383
rect 5442 3380 5448 3392
rect 4755 3352 5448 3380
rect 4755 3349 4767 3352
rect 4709 3343 4767 3349
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 7282 3380 7288 3392
rect 5592 3352 7288 3380
rect 5592 3340 5598 3352
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7561 3383 7619 3389
rect 7561 3349 7573 3383
rect 7607 3380 7619 3383
rect 7834 3380 7840 3392
rect 7607 3352 7840 3380
rect 7607 3349 7619 3352
rect 7561 3343 7619 3349
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 7944 3389 7972 3420
rect 8389 3417 8401 3420
rect 8435 3417 8447 3451
rect 8389 3411 8447 3417
rect 7929 3383 7987 3389
rect 7929 3349 7941 3383
rect 7975 3349 7987 3383
rect 7929 3343 7987 3349
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 8956 3380 8984 3479
rect 9122 3476 9128 3528
rect 9180 3476 9186 3528
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9306 3516 9312 3528
rect 9263 3488 9312 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10321 3519 10379 3525
rect 10321 3516 10333 3519
rect 10008 3488 10333 3516
rect 10008 3476 10014 3488
rect 10321 3485 10333 3488
rect 10367 3516 10379 3519
rect 11348 3516 11376 3556
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 14550 3584 14556 3596
rect 14511 3556 14556 3584
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 15764 3593 15792 3624
rect 15930 3612 15936 3624
rect 15988 3612 15994 3664
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 17184 3624 17540 3652
rect 17184 3612 17190 3624
rect 14737 3587 14795 3593
rect 14737 3553 14749 3587
rect 14783 3584 14795 3587
rect 15749 3587 15807 3593
rect 14783 3556 15056 3584
rect 14783 3553 14795 3556
rect 14737 3547 14795 3553
rect 10367 3488 11376 3516
rect 12253 3519 12311 3525
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 12434 3516 12440 3528
rect 12299 3488 12440 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 12434 3476 12440 3488
rect 12492 3476 12498 3528
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 12636 3488 14933 3516
rect 9140 3448 9168 3476
rect 9490 3448 9496 3460
rect 9140 3420 9496 3448
rect 9490 3408 9496 3420
rect 9548 3408 9554 3460
rect 9674 3408 9680 3460
rect 9732 3448 9738 3460
rect 10045 3451 10103 3457
rect 10045 3448 10057 3451
rect 9732 3420 10057 3448
rect 9732 3408 9738 3420
rect 9968 3392 9996 3420
rect 10045 3417 10057 3420
rect 10091 3417 10103 3451
rect 10045 3411 10103 3417
rect 10588 3451 10646 3457
rect 10588 3417 10600 3451
rect 10634 3448 10646 3451
rect 11238 3448 11244 3460
rect 10634 3420 11244 3448
rect 10634 3417 10646 3420
rect 10588 3411 10646 3417
rect 11238 3408 11244 3420
rect 11296 3408 11302 3460
rect 11977 3451 12035 3457
rect 11977 3417 11989 3451
rect 12023 3448 12035 3451
rect 12636 3448 12664 3488
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 14921 3479 14979 3485
rect 12802 3457 12808 3460
rect 12023 3420 12664 3448
rect 12023 3417 12035 3420
rect 11977 3411 12035 3417
rect 12796 3411 12808 3457
rect 12860 3448 12866 3460
rect 15028 3448 15056 3556
rect 15749 3553 15761 3587
rect 15795 3553 15807 3587
rect 15749 3547 15807 3553
rect 16761 3587 16819 3593
rect 16761 3553 16773 3587
rect 16807 3584 16819 3587
rect 17218 3584 17224 3596
rect 16807 3556 17224 3584
rect 16807 3553 16819 3556
rect 16761 3547 16819 3553
rect 17218 3544 17224 3556
rect 17276 3544 17282 3596
rect 17512 3593 17540 3624
rect 18598 3612 18604 3664
rect 18656 3612 18662 3664
rect 18874 3612 18880 3664
rect 18932 3652 18938 3664
rect 19337 3655 19395 3661
rect 19337 3652 19349 3655
rect 18932 3624 19349 3652
rect 18932 3612 18938 3624
rect 19337 3621 19349 3624
rect 19383 3621 19395 3655
rect 19337 3615 19395 3621
rect 19613 3655 19671 3661
rect 19613 3621 19625 3655
rect 19659 3652 19671 3655
rect 20990 3652 20996 3664
rect 19659 3624 20996 3652
rect 19659 3621 19671 3624
rect 19613 3615 19671 3621
rect 20990 3612 20996 3624
rect 21048 3612 21054 3664
rect 17497 3587 17555 3593
rect 17497 3553 17509 3587
rect 17543 3584 17555 3587
rect 18325 3587 18383 3593
rect 18325 3584 18337 3587
rect 17543 3556 18337 3584
rect 17543 3553 17555 3556
rect 17497 3547 17555 3553
rect 18325 3553 18337 3556
rect 18371 3553 18383 3587
rect 18325 3547 18383 3553
rect 18509 3587 18567 3593
rect 18509 3553 18521 3587
rect 18555 3584 18567 3587
rect 18616 3584 18644 3612
rect 19242 3584 19248 3596
rect 18555 3556 19248 3584
rect 18555 3553 18567 3556
rect 18509 3547 18567 3553
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 20898 3584 20904 3596
rect 19444 3556 20904 3584
rect 15473 3519 15531 3525
rect 15473 3485 15485 3519
rect 15519 3516 15531 3519
rect 15654 3516 15660 3528
rect 15519 3488 15660 3516
rect 15519 3485 15531 3488
rect 15473 3479 15531 3485
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 15838 3476 15844 3528
rect 15896 3516 15902 3528
rect 15933 3519 15991 3525
rect 15933 3516 15945 3519
rect 15896 3488 15945 3516
rect 15896 3476 15902 3488
rect 15933 3485 15945 3488
rect 15979 3485 15991 3519
rect 15933 3479 15991 3485
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 16209 3519 16267 3525
rect 16209 3516 16221 3519
rect 16080 3488 16221 3516
rect 16080 3476 16086 3488
rect 16209 3485 16221 3488
rect 16255 3485 16267 3519
rect 16209 3479 16267 3485
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17129 3519 17187 3525
rect 17129 3516 17141 3519
rect 17092 3488 17141 3516
rect 17092 3476 17098 3488
rect 17129 3485 17141 3488
rect 17175 3485 17187 3519
rect 17129 3479 17187 3485
rect 17310 3476 17316 3528
rect 17368 3516 17374 3528
rect 19444 3525 19472 3556
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 17773 3519 17831 3525
rect 17773 3516 17785 3519
rect 17368 3488 17785 3516
rect 17368 3476 17374 3488
rect 17773 3485 17785 3488
rect 17819 3485 17831 3519
rect 17773 3479 17831 3485
rect 18601 3519 18659 3525
rect 18601 3485 18613 3519
rect 18647 3516 18659 3519
rect 19429 3519 19487 3525
rect 18647 3488 19380 3516
rect 18647 3485 18659 3488
rect 18601 3479 18659 3485
rect 15565 3451 15623 3457
rect 15565 3448 15577 3451
rect 12860 3420 12896 3448
rect 13924 3420 15056 3448
rect 15120 3420 15577 3448
rect 8352 3352 8984 3380
rect 8352 3340 8358 3352
rect 9950 3340 9956 3392
rect 10008 3340 10014 3392
rect 10962 3340 10968 3392
rect 11020 3380 11026 3392
rect 11992 3380 12020 3411
rect 12802 3408 12808 3411
rect 12860 3408 12866 3420
rect 11020 3352 12020 3380
rect 12437 3383 12495 3389
rect 11020 3340 11026 3352
rect 12437 3349 12449 3383
rect 12483 3380 12495 3383
rect 13354 3380 13360 3392
rect 12483 3352 13360 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 13722 3340 13728 3392
rect 13780 3380 13786 3392
rect 13924 3389 13952 3420
rect 13909 3383 13967 3389
rect 13909 3380 13921 3383
rect 13780 3352 13921 3380
rect 13780 3340 13786 3352
rect 13909 3349 13921 3352
rect 13955 3349 13967 3383
rect 13909 3343 13967 3349
rect 14093 3383 14151 3389
rect 14093 3349 14105 3383
rect 14139 3380 14151 3383
rect 14274 3380 14280 3392
rect 14139 3352 14280 3380
rect 14139 3349 14151 3352
rect 14093 3343 14151 3349
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 14458 3380 14464 3392
rect 14419 3352 14464 3380
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 14918 3340 14924 3392
rect 14976 3380 14982 3392
rect 15120 3380 15148 3420
rect 15565 3417 15577 3420
rect 15611 3448 15623 3451
rect 16850 3448 16856 3460
rect 15611 3420 16856 3448
rect 15611 3417 15623 3420
rect 15565 3411 15623 3417
rect 16850 3408 16856 3420
rect 16908 3408 16914 3460
rect 19150 3448 19156 3460
rect 17328 3420 19156 3448
rect 14976 3352 15148 3380
rect 14976 3340 14982 3352
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 16117 3383 16175 3389
rect 16117 3380 16129 3383
rect 15988 3352 16129 3380
rect 15988 3340 15994 3352
rect 16117 3349 16129 3352
rect 16163 3349 16175 3383
rect 16390 3380 16396 3392
rect 16351 3352 16396 3380
rect 16117 3343 16175 3349
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 17328 3389 17356 3420
rect 19150 3408 19156 3420
rect 19208 3408 19214 3460
rect 19352 3448 19380 3488
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 19610 3476 19616 3528
rect 19668 3516 19674 3528
rect 19705 3519 19763 3525
rect 19705 3516 19717 3519
rect 19668 3488 19717 3516
rect 19668 3476 19674 3488
rect 19705 3485 19717 3488
rect 19751 3485 19763 3519
rect 19705 3479 19763 3485
rect 19886 3476 19892 3528
rect 19944 3516 19950 3528
rect 20070 3516 20076 3528
rect 19944 3488 20076 3516
rect 19944 3476 19950 3488
rect 20070 3476 20076 3488
rect 20128 3516 20134 3528
rect 20165 3519 20223 3525
rect 20165 3516 20177 3519
rect 20128 3488 20177 3516
rect 20128 3476 20134 3488
rect 20165 3485 20177 3488
rect 20211 3485 20223 3519
rect 20622 3516 20628 3528
rect 20583 3488 20628 3516
rect 20165 3479 20223 3485
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 20993 3519 21051 3525
rect 20772 3488 20817 3516
rect 20772 3476 20778 3488
rect 20993 3485 21005 3519
rect 21039 3516 21051 3519
rect 21082 3516 21088 3528
rect 21039 3488 21088 3516
rect 21039 3485 21051 3488
rect 20993 3479 21051 3485
rect 21082 3476 21088 3488
rect 21140 3476 21146 3528
rect 20898 3448 20904 3460
rect 19352 3420 20904 3448
rect 20898 3408 20904 3420
rect 20956 3408 20962 3460
rect 17313 3383 17371 3389
rect 17313 3349 17325 3383
rect 17359 3349 17371 3383
rect 17313 3343 17371 3349
rect 17681 3383 17739 3389
rect 17681 3349 17693 3383
rect 17727 3380 17739 3383
rect 19889 3383 19947 3389
rect 19889 3380 19901 3383
rect 17727 3352 19901 3380
rect 17727 3349 17739 3352
rect 17681 3343 17739 3349
rect 19889 3349 19901 3352
rect 19935 3380 19947 3383
rect 20162 3380 20168 3392
rect 19935 3352 20168 3380
rect 19935 3349 19947 3352
rect 19889 3343 19947 3349
rect 20162 3340 20168 3352
rect 20220 3340 20226 3392
rect 20441 3383 20499 3389
rect 20441 3349 20453 3383
rect 20487 3380 20499 3383
rect 21358 3380 21364 3392
rect 20487 3352 21364 3380
rect 20487 3349 20499 3352
rect 20441 3343 20499 3349
rect 21358 3340 21364 3352
rect 21416 3340 21422 3392
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 2406 3176 2412 3188
rect 2367 3148 2412 3176
rect 2406 3136 2412 3148
rect 2464 3136 2470 3188
rect 2682 3176 2688 3188
rect 2643 3148 2688 3176
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 3142 3176 3148 3188
rect 3007 3148 3148 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 5353 3179 5411 3185
rect 5353 3176 5365 3179
rect 3384 3148 5365 3176
rect 3384 3136 3390 3148
rect 5353 3145 5365 3148
rect 5399 3145 5411 3179
rect 5718 3176 5724 3188
rect 5679 3148 5724 3176
rect 5353 3139 5411 3145
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 6365 3179 6423 3185
rect 5868 3148 5913 3176
rect 5868 3136 5874 3148
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 6822 3176 6828 3188
rect 6411 3148 6828 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7006 3136 7012 3188
rect 7064 3176 7070 3188
rect 7064 3148 8616 3176
rect 7064 3136 7070 3148
rect 3418 3108 3424 3120
rect 3379 3080 3424 3108
rect 3418 3068 3424 3080
rect 3476 3068 3482 3120
rect 7190 3108 7196 3120
rect 3804 3080 7196 3108
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3040 2007 3043
rect 2130 3040 2136 3052
rect 1995 3012 2136 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 2498 3040 2504 3052
rect 2459 3012 2504 3040
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 3510 3040 3516 3052
rect 2777 3003 2835 3009
rect 3252 3012 3516 3040
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2682 2972 2688 2984
rect 2271 2944 2688 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 842 2864 848 2916
rect 900 2904 906 2916
rect 2792 2904 2820 3003
rect 3252 2981 3280 3012
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2941 3295 2975
rect 3237 2935 3295 2941
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2972 3387 2975
rect 3804 2972 3832 3080
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 7374 3068 7380 3120
rect 7432 3108 7438 3120
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 7432 3080 7849 3108
rect 7432 3068 7438 3080
rect 7837 3077 7849 3080
rect 7883 3077 7895 3111
rect 7837 3071 7895 3077
rect 7926 3068 7932 3120
rect 7984 3108 7990 3120
rect 8021 3111 8079 3117
rect 8021 3108 8033 3111
rect 7984 3080 8033 3108
rect 7984 3068 7990 3080
rect 8021 3077 8033 3080
rect 8067 3077 8079 3111
rect 8021 3071 8079 3077
rect 8110 3068 8116 3120
rect 8168 3108 8174 3120
rect 8450 3111 8508 3117
rect 8450 3108 8462 3111
rect 8168 3080 8462 3108
rect 8168 3068 8174 3080
rect 8450 3077 8462 3080
rect 8496 3077 8508 3111
rect 8450 3071 8508 3077
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 4154 3049 4160 3052
rect 4148 3040 4160 3049
rect 3936 3012 3981 3040
rect 4115 3012 4160 3040
rect 3936 3000 3942 3012
rect 4148 3003 4160 3012
rect 4154 3000 4160 3003
rect 4212 3000 4218 3052
rect 7489 3043 7547 3049
rect 7489 3009 7501 3043
rect 7535 3040 7547 3043
rect 8202 3040 8208 3052
rect 7535 3012 7972 3040
rect 8163 3012 8208 3040
rect 7535 3009 7547 3012
rect 7489 3003 7547 3009
rect 3375 2944 3832 2972
rect 3375 2941 3387 2944
rect 3329 2935 3387 2941
rect 4890 2932 4896 2984
rect 4948 2972 4954 2984
rect 5902 2972 5908 2984
rect 4948 2944 5908 2972
rect 4948 2932 4954 2944
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 7742 2972 7748 2984
rect 7703 2944 7748 2972
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 5810 2904 5816 2916
rect 900 2876 3924 2904
rect 900 2864 906 2876
rect 3142 2796 3148 2848
rect 3200 2836 3206 2848
rect 3789 2839 3847 2845
rect 3789 2836 3801 2839
rect 3200 2808 3801 2836
rect 3200 2796 3206 2808
rect 3789 2805 3801 2808
rect 3835 2805 3847 2839
rect 3896 2836 3924 2876
rect 4816 2876 5816 2904
rect 4816 2836 4844 2876
rect 5810 2864 5816 2876
rect 5868 2864 5874 2916
rect 3896 2808 4844 2836
rect 5261 2839 5319 2845
rect 3789 2799 3847 2805
rect 5261 2805 5273 2839
rect 5307 2836 5319 2839
rect 5350 2836 5356 2848
rect 5307 2808 5356 2836
rect 5307 2805 5319 2808
rect 5261 2799 5319 2805
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 5994 2796 6000 2848
rect 6052 2836 6058 2848
rect 7760 2836 7788 2932
rect 6052 2808 7788 2836
rect 7944 2836 7972 3012
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8588 3040 8616 3148
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 9677 3179 9735 3185
rect 9677 3176 9689 3179
rect 8812 3148 9689 3176
rect 8812 3136 8818 3148
rect 9677 3145 9689 3148
rect 9723 3145 9735 3179
rect 9677 3139 9735 3145
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 9824 3148 10057 3176
rect 9824 3136 9830 3148
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 10045 3139 10103 3145
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 10505 3179 10563 3185
rect 10192 3148 10237 3176
rect 10192 3136 10198 3148
rect 10505 3145 10517 3179
rect 10551 3145 10563 3179
rect 10505 3139 10563 3145
rect 9214 3068 9220 3120
rect 9272 3108 9278 3120
rect 10520 3108 10548 3139
rect 10870 3136 10876 3188
rect 10928 3176 10934 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 10928 3148 10977 3176
rect 10928 3136 10934 3148
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 10965 3139 11023 3145
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 12066 3176 12072 3188
rect 11940 3148 12072 3176
rect 11940 3136 11946 3148
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 13446 3176 13452 3188
rect 12860 3148 13452 3176
rect 12860 3136 12866 3148
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 13722 3176 13728 3188
rect 13565 3148 13728 3176
rect 9272 3080 10548 3108
rect 10621 3080 11008 3108
rect 9272 3068 9278 3080
rect 10621 3040 10649 3080
rect 8588 3012 10649 3040
rect 10686 3000 10692 3052
rect 10744 3040 10750 3052
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 10744 3012 10885 3040
rect 10744 3000 10750 3012
rect 10873 3009 10885 3012
rect 10919 3009 10931 3043
rect 10980 3040 11008 3080
rect 11146 3068 11152 3120
rect 11204 3108 11210 3120
rect 11977 3111 12035 3117
rect 11977 3108 11989 3111
rect 11204 3080 11989 3108
rect 11204 3068 11210 3080
rect 11977 3077 11989 3080
rect 12023 3108 12035 3111
rect 12158 3108 12164 3120
rect 12023 3080 12164 3108
rect 12023 3077 12035 3080
rect 11977 3071 12035 3077
rect 12158 3068 12164 3080
rect 12216 3068 12222 3120
rect 13565 3117 13593 3148
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 13909 3179 13967 3185
rect 13909 3176 13921 3179
rect 13872 3148 13921 3176
rect 13872 3136 13878 3148
rect 13909 3145 13921 3148
rect 13955 3145 13967 3179
rect 13909 3139 13967 3145
rect 14277 3179 14335 3185
rect 14277 3145 14289 3179
rect 14323 3176 14335 3179
rect 14366 3176 14372 3188
rect 14323 3148 14372 3176
rect 14323 3145 14335 3148
rect 14277 3139 14335 3145
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 15010 3176 15016 3188
rect 14752 3148 15016 3176
rect 13550 3111 13608 3117
rect 13550 3077 13562 3111
rect 13596 3077 13608 3111
rect 13550 3071 13608 3077
rect 10980 3012 12020 3040
rect 10873 3003 10931 3009
rect 11992 2984 12020 3012
rect 13170 3000 13176 3052
rect 13228 3040 13234 3052
rect 14642 3040 14648 3052
rect 13228 3012 14648 3040
rect 13228 3000 13234 3012
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 10321 2975 10379 2981
rect 10321 2972 10333 2975
rect 9364 2944 10333 2972
rect 9364 2932 9370 2944
rect 10321 2941 10333 2944
rect 10367 2972 10379 2975
rect 11057 2975 11115 2981
rect 11057 2972 11069 2975
rect 10367 2944 11069 2972
rect 10367 2941 10379 2944
rect 10321 2935 10379 2941
rect 11057 2941 11069 2944
rect 11103 2941 11115 2975
rect 11057 2935 11115 2941
rect 11974 2932 11980 2984
rect 12032 2972 12038 2984
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 12032 2944 12081 2972
rect 12032 2932 12038 2944
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 13814 2972 13820 2984
rect 13775 2944 13820 2972
rect 12069 2935 12127 2941
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 14366 2972 14372 2984
rect 14327 2944 14372 2972
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 14553 2975 14611 2981
rect 14553 2941 14565 2975
rect 14599 2972 14611 2975
rect 14752 2972 14780 3148
rect 15010 3136 15016 3148
rect 15068 3136 15074 3188
rect 15286 3136 15292 3188
rect 15344 3176 15350 3188
rect 15473 3179 15531 3185
rect 15344 3148 15424 3176
rect 15344 3136 15350 3148
rect 15194 3108 15200 3120
rect 15028 3080 15200 3108
rect 14918 3040 14924 3052
rect 14879 3012 14924 3040
rect 14918 3000 14924 3012
rect 14976 3000 14982 3052
rect 15028 3049 15056 3080
rect 15194 3068 15200 3080
rect 15252 3068 15258 3120
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3009 15071 3043
rect 15286 3040 15292 3052
rect 15247 3012 15292 3040
rect 15013 3003 15071 3009
rect 15286 3000 15292 3012
rect 15344 3000 15350 3052
rect 14599 2944 14780 2972
rect 15396 2972 15424 3148
rect 15473 3145 15485 3179
rect 15519 3145 15531 3179
rect 15473 3139 15531 3145
rect 15488 3040 15516 3139
rect 16390 3136 16396 3188
rect 16448 3176 16454 3188
rect 17405 3179 17463 3185
rect 16448 3148 17356 3176
rect 16448 3136 16454 3148
rect 15930 3068 15936 3120
rect 15988 3108 15994 3120
rect 15988 3080 16988 3108
rect 15988 3068 15994 3080
rect 15565 3043 15623 3049
rect 15565 3040 15577 3043
rect 15488 3012 15577 3040
rect 15565 3009 15577 3012
rect 15611 3009 15623 3043
rect 15565 3003 15623 3009
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 16132 2972 16160 3003
rect 16206 3000 16212 3052
rect 16264 3040 16270 3052
rect 16264 3012 16309 3040
rect 16264 3000 16270 3012
rect 16482 3000 16488 3052
rect 16540 3040 16546 3052
rect 16960 3049 16988 3080
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16540 3012 16681 3040
rect 16540 3000 16546 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3009 17003 3043
rect 16945 3003 17003 3009
rect 17034 3000 17040 3052
rect 17092 3040 17098 3052
rect 17221 3043 17279 3049
rect 17221 3040 17233 3043
rect 17092 3012 17233 3040
rect 17092 3000 17098 3012
rect 17221 3009 17233 3012
rect 17267 3009 17279 3043
rect 17328 3040 17356 3148
rect 17405 3145 17417 3179
rect 17451 3176 17463 3179
rect 18138 3176 18144 3188
rect 17451 3148 18144 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 18693 3179 18751 3185
rect 18693 3145 18705 3179
rect 18739 3145 18751 3179
rect 18693 3139 18751 3145
rect 17497 3043 17555 3049
rect 17497 3040 17509 3043
rect 17328 3012 17509 3040
rect 17221 3003 17279 3009
rect 17497 3009 17509 3012
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 17586 3000 17592 3052
rect 17644 3040 17650 3052
rect 17773 3043 17831 3049
rect 17773 3040 17785 3043
rect 17644 3012 17785 3040
rect 17644 3000 17650 3012
rect 17773 3009 17785 3012
rect 17819 3009 17831 3043
rect 17773 3003 17831 3009
rect 18046 3000 18052 3052
rect 18104 3040 18110 3052
rect 18141 3043 18199 3049
rect 18141 3040 18153 3043
rect 18104 3012 18153 3040
rect 18104 3000 18110 3012
rect 18141 3009 18153 3012
rect 18187 3009 18199 3043
rect 18506 3040 18512 3052
rect 18467 3012 18512 3040
rect 18141 3003 18199 3009
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 18708 3040 18736 3139
rect 19242 3136 19248 3188
rect 19300 3176 19306 3188
rect 21082 3176 21088 3188
rect 19300 3148 21088 3176
rect 19300 3136 19306 3148
rect 21082 3136 21088 3148
rect 21140 3136 21146 3188
rect 18877 3043 18935 3049
rect 18877 3040 18889 3043
rect 18708 3012 18889 3040
rect 18877 3009 18889 3012
rect 18923 3009 18935 3043
rect 18877 3003 18935 3009
rect 19150 3000 19156 3052
rect 19208 3040 19214 3052
rect 19245 3043 19303 3049
rect 19245 3040 19257 3043
rect 19208 3012 19257 3040
rect 19208 3000 19214 3012
rect 19245 3009 19257 3012
rect 19291 3009 19303 3043
rect 19610 3040 19616 3052
rect 19571 3012 19616 3040
rect 19245 3003 19303 3009
rect 19610 3000 19616 3012
rect 19668 3000 19674 3052
rect 20254 3040 20260 3052
rect 20215 3012 20260 3040
rect 20254 3000 20260 3012
rect 20312 3000 20318 3052
rect 20346 3000 20352 3052
rect 20404 3040 20410 3052
rect 20717 3043 20775 3049
rect 20404 3012 20449 3040
rect 20404 3000 20410 3012
rect 20717 3009 20729 3043
rect 20763 3040 20775 3043
rect 21634 3040 21640 3052
rect 20763 3012 21640 3040
rect 20763 3009 20775 3012
rect 20717 3003 20775 3009
rect 21634 3000 21640 3012
rect 21692 3040 21698 3052
rect 22738 3040 22744 3052
rect 21692 3012 22744 3040
rect 21692 3000 21698 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 17402 2972 17408 2984
rect 15396 2944 17408 2972
rect 14599 2941 14611 2944
rect 14553 2935 14611 2941
rect 8570 2836 8576 2848
rect 7944 2808 8576 2836
rect 6052 2796 6058 2808
rect 8570 2796 8576 2808
rect 8628 2836 8634 2848
rect 9324 2836 9352 2932
rect 9582 2904 9588 2916
rect 9543 2876 9588 2904
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 11238 2864 11244 2916
rect 11296 2904 11302 2916
rect 12437 2907 12495 2913
rect 12437 2904 12449 2907
rect 11296 2876 12449 2904
rect 11296 2864 11302 2876
rect 12437 2873 12449 2876
rect 12483 2873 12495 2907
rect 12437 2867 12495 2873
rect 8628 2808 9352 2836
rect 8628 2796 8634 2808
rect 11146 2796 11152 2848
rect 11204 2836 11210 2848
rect 11517 2839 11575 2845
rect 11517 2836 11529 2839
rect 11204 2808 11529 2836
rect 11204 2796 11210 2808
rect 11517 2805 11529 2808
rect 11563 2805 11575 2839
rect 11517 2799 11575 2805
rect 11698 2796 11704 2848
rect 11756 2836 11762 2848
rect 12158 2836 12164 2848
rect 11756 2808 12164 2836
rect 11756 2796 11762 2808
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 12452 2836 12480 2867
rect 13078 2836 13084 2848
rect 12452 2808 13084 2836
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 13446 2796 13452 2848
rect 13504 2836 13510 2848
rect 14568 2836 14596 2935
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 18966 2972 18972 2984
rect 17696 2944 18972 2972
rect 15562 2864 15568 2916
rect 15620 2904 15626 2916
rect 16482 2904 16488 2916
rect 15620 2876 16488 2904
rect 15620 2864 15626 2876
rect 16482 2864 16488 2876
rect 16540 2864 16546 2916
rect 16853 2907 16911 2913
rect 16853 2873 16865 2907
rect 16899 2904 16911 2907
rect 17310 2904 17316 2916
rect 16899 2876 17316 2904
rect 16899 2873 16911 2876
rect 16853 2867 16911 2873
rect 17310 2864 17316 2876
rect 17368 2864 17374 2916
rect 17696 2913 17724 2944
rect 18966 2932 18972 2944
rect 19024 2932 19030 2984
rect 20806 2932 20812 2984
rect 20864 2972 20870 2984
rect 20993 2975 21051 2981
rect 20993 2972 21005 2975
rect 20864 2944 21005 2972
rect 20864 2932 20870 2944
rect 20993 2941 21005 2944
rect 21039 2941 21051 2975
rect 20993 2935 21051 2941
rect 17681 2907 17739 2913
rect 17681 2873 17693 2907
rect 17727 2873 17739 2907
rect 17681 2867 17739 2873
rect 18046 2864 18052 2916
rect 18104 2904 18110 2916
rect 18325 2907 18383 2913
rect 18325 2904 18337 2907
rect 18104 2876 18337 2904
rect 18104 2864 18110 2876
rect 18325 2873 18337 2876
rect 18371 2873 18383 2907
rect 18325 2867 18383 2873
rect 20073 2907 20131 2913
rect 20073 2873 20085 2907
rect 20119 2904 20131 2907
rect 20622 2904 20628 2916
rect 20119 2876 20628 2904
rect 20119 2873 20131 2876
rect 20073 2867 20131 2873
rect 20622 2864 20628 2876
rect 20680 2864 20686 2916
rect 14734 2836 14740 2848
rect 13504 2808 14596 2836
rect 14695 2808 14740 2836
rect 13504 2796 13510 2808
rect 14734 2796 14740 2808
rect 14792 2796 14798 2848
rect 15194 2836 15200 2848
rect 15155 2808 15200 2836
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 15470 2796 15476 2848
rect 15528 2836 15534 2848
rect 15749 2839 15807 2845
rect 15749 2836 15761 2839
rect 15528 2808 15761 2836
rect 15528 2796 15534 2808
rect 15749 2805 15761 2808
rect 15795 2805 15807 2839
rect 15930 2836 15936 2848
rect 15891 2808 15936 2836
rect 15749 2799 15807 2805
rect 15930 2796 15936 2808
rect 15988 2796 15994 2848
rect 16390 2836 16396 2848
rect 16351 2808 16396 2836
rect 16390 2796 16396 2808
rect 16448 2796 16454 2848
rect 17126 2836 17132 2848
rect 17087 2808 17132 2836
rect 17126 2796 17132 2808
rect 17184 2796 17190 2848
rect 17957 2839 18015 2845
rect 17957 2805 17969 2839
rect 18003 2836 18015 2839
rect 18230 2836 18236 2848
rect 18003 2808 18236 2836
rect 18003 2805 18015 2808
rect 17957 2799 18015 2805
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 18782 2796 18788 2848
rect 18840 2836 18846 2848
rect 19061 2839 19119 2845
rect 19061 2836 19073 2839
rect 18840 2808 19073 2836
rect 18840 2796 18846 2808
rect 19061 2805 19073 2808
rect 19107 2805 19119 2839
rect 19061 2799 19119 2805
rect 19150 2796 19156 2848
rect 19208 2836 19214 2848
rect 19429 2839 19487 2845
rect 19429 2836 19441 2839
rect 19208 2808 19441 2836
rect 19208 2796 19214 2808
rect 19429 2805 19441 2808
rect 19475 2805 19487 2839
rect 19429 2799 19487 2805
rect 19518 2796 19524 2848
rect 19576 2836 19582 2848
rect 19797 2839 19855 2845
rect 19797 2836 19809 2839
rect 19576 2808 19809 2836
rect 19576 2796 19582 2808
rect 19797 2805 19809 2808
rect 19843 2805 19855 2839
rect 19797 2799 19855 2805
rect 20254 2796 20260 2848
rect 20312 2836 20318 2848
rect 20533 2839 20591 2845
rect 20533 2836 20545 2839
rect 20312 2808 20545 2836
rect 20312 2796 20318 2808
rect 20533 2805 20545 2808
rect 20579 2805 20591 2839
rect 20533 2799 20591 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 3142 2592 3148 2644
rect 3200 2632 3206 2644
rect 3200 2604 4936 2632
rect 3200 2592 3206 2604
rect 3605 2567 3663 2573
rect 3605 2533 3617 2567
rect 3651 2564 3663 2567
rect 4706 2564 4712 2576
rect 3651 2536 4712 2564
rect 3651 2533 3663 2536
rect 3605 2527 3663 2533
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 4908 2564 4936 2604
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 5040 2604 5089 2632
rect 5040 2592 5046 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 5077 2595 5135 2601
rect 6546 2592 6552 2644
rect 6604 2632 6610 2644
rect 7101 2635 7159 2641
rect 7101 2632 7113 2635
rect 6604 2604 7113 2632
rect 6604 2592 6610 2604
rect 7101 2601 7113 2604
rect 7147 2601 7159 2635
rect 7101 2595 7159 2601
rect 7929 2635 7987 2641
rect 7929 2601 7941 2635
rect 7975 2632 7987 2635
rect 8018 2632 8024 2644
rect 7975 2604 8024 2632
rect 7975 2601 7987 2604
rect 7929 2595 7987 2601
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 8202 2592 8208 2644
rect 8260 2632 8266 2644
rect 9033 2635 9091 2641
rect 9033 2632 9045 2635
rect 8260 2604 9045 2632
rect 8260 2592 8266 2604
rect 9033 2601 9045 2604
rect 9079 2601 9091 2635
rect 9033 2595 9091 2601
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 11882 2632 11888 2644
rect 11747 2604 11888 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12529 2635 12587 2641
rect 12529 2601 12541 2635
rect 12575 2632 12587 2635
rect 12618 2632 12624 2644
rect 12575 2604 12624 2632
rect 12575 2601 12587 2604
rect 12529 2595 12587 2601
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 13906 2632 13912 2644
rect 13565 2604 13912 2632
rect 5258 2564 5264 2576
rect 4908 2536 5264 2564
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 8478 2564 8484 2576
rect 5368 2536 8484 2564
rect 1946 2496 1952 2508
rect 1907 2468 1952 2496
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 3142 2496 3148 2508
rect 3103 2468 3148 2496
rect 3142 2456 3148 2468
rect 3200 2456 3206 2508
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 3752 2468 4629 2496
rect 3752 2456 3758 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 4801 2499 4859 2505
rect 4801 2465 4813 2499
rect 4847 2496 4859 2499
rect 5368 2496 5396 2536
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 9398 2524 9404 2576
rect 9456 2564 9462 2576
rect 11146 2564 11152 2576
rect 9456 2536 11152 2564
rect 9456 2524 9462 2536
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 12250 2524 12256 2576
rect 12308 2564 12314 2576
rect 13565 2564 13593 2604
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 15013 2635 15071 2641
rect 15013 2632 15025 2635
rect 14056 2604 15025 2632
rect 14056 2592 14062 2604
rect 15013 2601 15025 2604
rect 15059 2601 15071 2635
rect 15013 2595 15071 2601
rect 15838 2592 15844 2644
rect 15896 2632 15902 2644
rect 16758 2632 16764 2644
rect 15896 2604 16764 2632
rect 15896 2592 15902 2604
rect 16758 2592 16764 2604
rect 16816 2592 16822 2644
rect 17221 2635 17279 2641
rect 17221 2632 17233 2635
rect 16868 2604 17233 2632
rect 12308 2536 13593 2564
rect 12308 2524 12314 2536
rect 13630 2524 13636 2576
rect 13688 2564 13694 2576
rect 14553 2567 14611 2573
rect 14553 2564 14565 2567
rect 13688 2536 14565 2564
rect 13688 2524 13694 2536
rect 14553 2533 14565 2536
rect 14599 2533 14611 2567
rect 14553 2527 14611 2533
rect 15102 2524 15108 2576
rect 15160 2564 15166 2576
rect 15160 2536 15608 2564
rect 15160 2524 15166 2536
rect 4847 2468 5396 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 5442 2456 5448 2508
rect 5500 2496 5506 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5500 2468 5733 2496
rect 5500 2456 5506 2468
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 5902 2456 5908 2508
rect 5960 2496 5966 2508
rect 6546 2496 6552 2508
rect 5960 2468 6552 2496
rect 5960 2456 5966 2468
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 7374 2496 7380 2508
rect 7287 2468 7380 2496
rect 7374 2456 7380 2468
rect 7432 2496 7438 2508
rect 8294 2496 8300 2508
rect 7432 2468 8300 2496
rect 7432 2456 7438 2468
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 8570 2496 8576 2508
rect 8531 2468 8576 2496
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 10318 2496 10324 2508
rect 9232 2468 10324 2496
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2774 2428 2780 2440
rect 2271 2400 2780 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 2866 2388 2872 2440
rect 2924 2428 2930 2440
rect 2924 2400 2969 2428
rect 2924 2388 2930 2400
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3292 2400 4292 2428
rect 3292 2388 3298 2400
rect 3421 2363 3479 2369
rect 3421 2329 3433 2363
rect 3467 2360 3479 2363
rect 3510 2360 3516 2372
rect 3467 2332 3516 2360
rect 3467 2329 3479 2332
rect 3421 2323 3479 2329
rect 3510 2320 3516 2332
rect 3568 2320 3574 2372
rect 4264 2360 4292 2400
rect 4338 2388 4344 2440
rect 4396 2428 4402 2440
rect 4396 2400 4441 2428
rect 4396 2388 4402 2400
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 5224 2400 6745 2428
rect 5224 2388 5230 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7248 2400 7481 2428
rect 7248 2388 7254 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 9232 2437 9260 2468
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 10778 2496 10784 2508
rect 10739 2468 10784 2496
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 13078 2496 13084 2508
rect 13039 2468 13084 2496
rect 13078 2456 13084 2468
rect 13136 2456 13142 2508
rect 14274 2496 14280 2508
rect 13188 2468 14280 2496
rect 9217 2431 9275 2437
rect 7616 2400 7661 2428
rect 7616 2388 7622 2400
rect 9217 2397 9229 2431
rect 9263 2397 9275 2431
rect 9858 2428 9864 2440
rect 9819 2400 9864 2428
rect 9217 2391 9275 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 10134 2428 10140 2440
rect 10095 2400 10140 2428
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 10686 2428 10692 2440
rect 10647 2400 10692 2428
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2428 11575 2431
rect 11698 2428 11704 2440
rect 11563 2400 11704 2428
rect 11563 2397 11575 2400
rect 11517 2391 11575 2397
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 12066 2428 12072 2440
rect 12027 2400 12072 2428
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 12894 2428 12900 2440
rect 12216 2400 12261 2428
rect 12855 2400 12900 2428
rect 12216 2388 12222 2400
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 12989 2431 13047 2437
rect 12989 2397 13001 2431
rect 13035 2428 13047 2431
rect 13188 2428 13216 2468
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 15286 2496 15292 2508
rect 14568 2468 15292 2496
rect 13354 2428 13360 2440
rect 13035 2400 13216 2428
rect 13315 2400 13360 2428
rect 13035 2397 13047 2400
rect 12989 2391 13047 2397
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 13722 2428 13728 2440
rect 13683 2400 13728 2428
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13964 2400 14105 2428
rect 13964 2388 13970 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 4982 2360 4988 2372
rect 4264 2332 4844 2360
rect 4943 2332 4988 2360
rect 4816 2292 4844 2332
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 5350 2320 5356 2372
rect 5408 2360 5414 2372
rect 6641 2363 6699 2369
rect 6641 2360 6653 2363
rect 5408 2332 6653 2360
rect 5408 2320 5414 2332
rect 6641 2329 6653 2332
rect 6687 2329 6699 2363
rect 6641 2323 6699 2329
rect 8389 2363 8447 2369
rect 8389 2329 8401 2363
rect 8435 2360 8447 2363
rect 9582 2360 9588 2372
rect 8435 2332 9588 2360
rect 8435 2329 8447 2332
rect 8389 2323 8447 2329
rect 9582 2320 9588 2332
rect 9640 2320 9646 2372
rect 5261 2295 5319 2301
rect 5261 2292 5273 2295
rect 4816 2264 5273 2292
rect 5261 2261 5273 2264
rect 5307 2261 5319 2295
rect 5626 2292 5632 2304
rect 5587 2264 5632 2292
rect 5261 2255 5319 2261
rect 5626 2252 5632 2264
rect 5684 2252 5690 2304
rect 6181 2295 6239 2301
rect 6181 2261 6193 2295
rect 6227 2292 6239 2295
rect 7742 2292 7748 2304
rect 6227 2264 7748 2292
rect 6227 2261 6239 2264
rect 6181 2255 6239 2261
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 7834 2252 7840 2304
rect 7892 2292 7898 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7892 2264 8033 2292
rect 7892 2252 7898 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 8202 2252 8208 2304
rect 8260 2292 8266 2304
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8260 2264 8493 2292
rect 8260 2252 8266 2264
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 8481 2255 8539 2261
rect 9214 2252 9220 2304
rect 9272 2292 9278 2304
rect 10152 2292 10180 2388
rect 11238 2360 11244 2372
rect 11151 2332 11244 2360
rect 11238 2320 11244 2332
rect 11296 2360 11302 2372
rect 12434 2360 12440 2372
rect 11296 2332 12440 2360
rect 11296 2320 11302 2332
rect 12434 2320 12440 2332
rect 12492 2320 12498 2372
rect 12526 2320 12532 2372
rect 12584 2360 12590 2372
rect 14568 2360 14596 2468
rect 15286 2456 15292 2468
rect 15344 2456 15350 2508
rect 14734 2428 14740 2440
rect 14695 2400 14740 2428
rect 14734 2388 14740 2400
rect 14792 2388 14798 2440
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2397 14887 2431
rect 15194 2428 15200 2440
rect 15155 2400 15200 2428
rect 14829 2391 14887 2397
rect 12584 2332 13124 2360
rect 12584 2320 12590 2332
rect 9272 2264 10180 2292
rect 9272 2252 9278 2264
rect 10226 2252 10232 2304
rect 10284 2292 10290 2304
rect 10594 2292 10600 2304
rect 10284 2264 10329 2292
rect 10555 2264 10600 2292
rect 10284 2252 10290 2264
rect 10594 2252 10600 2264
rect 10652 2252 10658 2304
rect 11146 2292 11152 2304
rect 11107 2264 11152 2292
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 11882 2292 11888 2304
rect 11843 2264 11888 2292
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 12345 2295 12403 2301
rect 12345 2261 12357 2295
rect 12391 2292 12403 2295
rect 12802 2292 12808 2304
rect 12391 2264 12808 2292
rect 12391 2261 12403 2264
rect 12345 2255 12403 2261
rect 12802 2252 12808 2264
rect 12860 2252 12866 2304
rect 13096 2292 13124 2332
rect 13924 2332 14596 2360
rect 13924 2301 13952 2332
rect 14642 2320 14648 2372
rect 14700 2360 14706 2372
rect 14844 2360 14872 2391
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 15580 2437 15608 2536
rect 16206 2524 16212 2576
rect 16264 2564 16270 2576
rect 16868 2564 16896 2604
rect 17221 2601 17233 2604
rect 17267 2601 17279 2635
rect 17221 2595 17279 2601
rect 17770 2592 17776 2644
rect 17828 2632 17834 2644
rect 18693 2635 18751 2641
rect 18693 2632 18705 2635
rect 17828 2604 18705 2632
rect 17828 2592 17834 2604
rect 18693 2601 18705 2604
rect 18739 2601 18751 2635
rect 18693 2595 18751 2601
rect 19061 2635 19119 2641
rect 19061 2601 19073 2635
rect 19107 2632 19119 2635
rect 19610 2632 19616 2644
rect 19107 2604 19616 2632
rect 19107 2601 19119 2604
rect 19061 2595 19119 2601
rect 19610 2592 19616 2604
rect 19668 2592 19674 2644
rect 19702 2592 19708 2644
rect 19760 2632 19766 2644
rect 19760 2604 19805 2632
rect 19760 2592 19766 2604
rect 16264 2536 16896 2564
rect 16264 2524 16270 2536
rect 16942 2524 16948 2576
rect 17000 2564 17006 2576
rect 17957 2567 18015 2573
rect 17957 2564 17969 2567
rect 17000 2536 17969 2564
rect 17000 2524 17006 2536
rect 17957 2533 17969 2536
rect 18003 2533 18015 2567
rect 17957 2527 18015 2533
rect 18414 2524 18420 2576
rect 18472 2564 18478 2576
rect 19429 2567 19487 2573
rect 19429 2564 19441 2567
rect 18472 2536 19441 2564
rect 18472 2524 18478 2536
rect 19429 2533 19441 2536
rect 19475 2533 19487 2567
rect 19429 2527 19487 2533
rect 17126 2456 17132 2508
rect 17184 2496 17190 2508
rect 17184 2468 17816 2496
rect 17184 2456 17190 2468
rect 15565 2431 15623 2437
rect 15565 2397 15577 2431
rect 15611 2397 15623 2431
rect 15930 2428 15936 2440
rect 15891 2400 15936 2428
rect 15565 2391 15623 2397
rect 15930 2388 15936 2400
rect 15988 2388 15994 2440
rect 16298 2428 16304 2440
rect 16259 2400 16304 2428
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 16390 2388 16396 2440
rect 16448 2428 16454 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16448 2400 16681 2428
rect 16448 2388 16454 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 14700 2332 14872 2360
rect 14700 2320 14706 2332
rect 15102 2320 15108 2372
rect 15160 2360 15166 2372
rect 17052 2360 17080 2391
rect 17310 2388 17316 2440
rect 17368 2428 17374 2440
rect 17405 2431 17463 2437
rect 17405 2428 17417 2431
rect 17368 2400 17417 2428
rect 17368 2388 17374 2400
rect 17405 2397 17417 2400
rect 17451 2397 17463 2431
rect 17405 2391 17463 2397
rect 17678 2388 17684 2440
rect 17736 2388 17742 2440
rect 17788 2437 17816 2468
rect 18322 2456 18328 2508
rect 18380 2496 18386 2508
rect 18380 2468 18920 2496
rect 18380 2456 18386 2468
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2397 17831 2431
rect 18138 2428 18144 2440
rect 18099 2400 18144 2428
rect 17773 2391 17831 2397
rect 18138 2388 18144 2400
rect 18196 2388 18202 2440
rect 18230 2388 18236 2440
rect 18288 2428 18294 2440
rect 18892 2437 18920 2468
rect 19150 2456 19156 2508
rect 19208 2496 19214 2508
rect 20714 2496 20720 2508
rect 19208 2468 20720 2496
rect 19208 2456 19214 2468
rect 20714 2456 20720 2468
rect 20772 2456 20778 2508
rect 20898 2456 20904 2508
rect 20956 2496 20962 2508
rect 20993 2499 21051 2505
rect 20993 2496 21005 2499
rect 20956 2468 21005 2496
rect 20956 2456 20962 2468
rect 20993 2465 21005 2468
rect 21039 2496 21051 2499
rect 22830 2496 22836 2508
rect 21039 2468 22836 2496
rect 21039 2465 21051 2468
rect 20993 2459 21051 2465
rect 22830 2456 22836 2468
rect 22888 2456 22894 2508
rect 18509 2431 18567 2437
rect 18509 2428 18521 2431
rect 18288 2400 18521 2428
rect 18288 2388 18294 2400
rect 18509 2397 18521 2400
rect 18555 2397 18567 2431
rect 18509 2391 18567 2397
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 18966 2388 18972 2440
rect 19024 2428 19030 2440
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 19024 2400 19257 2428
rect 19024 2388 19030 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2397 20407 2431
rect 20349 2391 20407 2397
rect 15160 2332 16160 2360
rect 15160 2320 15166 2332
rect 13541 2295 13599 2301
rect 13541 2292 13553 2295
rect 13096 2264 13553 2292
rect 13541 2261 13553 2264
rect 13587 2261 13599 2295
rect 13541 2255 13599 2261
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2261 13967 2295
rect 13909 2255 13967 2261
rect 14274 2252 14280 2304
rect 14332 2292 14338 2304
rect 14332 2264 14377 2292
rect 14332 2252 14338 2264
rect 14550 2252 14556 2304
rect 14608 2292 14614 2304
rect 15381 2295 15439 2301
rect 15381 2292 15393 2295
rect 14608 2264 15393 2292
rect 14608 2252 14614 2264
rect 15381 2261 15393 2264
rect 15427 2261 15439 2295
rect 15381 2255 15439 2261
rect 15654 2252 15660 2304
rect 15712 2292 15718 2304
rect 16132 2301 16160 2332
rect 16500 2332 17080 2360
rect 17696 2360 17724 2388
rect 20364 2360 20392 2391
rect 20530 2388 20536 2440
rect 20588 2428 20594 2440
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 20588 2400 20637 2428
rect 20588 2388 20594 2400
rect 20625 2397 20637 2400
rect 20671 2397 20683 2431
rect 20625 2391 20683 2397
rect 17696 2332 20392 2360
rect 16500 2301 16528 2332
rect 15749 2295 15807 2301
rect 15749 2292 15761 2295
rect 15712 2264 15761 2292
rect 15712 2252 15718 2264
rect 15749 2261 15761 2264
rect 15795 2261 15807 2295
rect 15749 2255 15807 2261
rect 16117 2295 16175 2301
rect 16117 2261 16129 2295
rect 16163 2261 16175 2295
rect 16117 2255 16175 2261
rect 16485 2295 16543 2301
rect 16485 2261 16497 2295
rect 16531 2261 16543 2295
rect 16485 2255 16543 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16816 2264 16865 2292
rect 16816 2252 16822 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 17586 2292 17592 2304
rect 17547 2264 17592 2292
rect 16853 2255 16911 2261
rect 17586 2252 17592 2264
rect 17644 2252 17650 2304
rect 17678 2252 17684 2304
rect 17736 2292 17742 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 17736 2264 18337 2292
rect 17736 2252 17742 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 6546 2048 6552 2100
rect 6604 2088 6610 2100
rect 10778 2088 10784 2100
rect 6604 2060 10784 2088
rect 6604 2048 6610 2060
rect 10778 2048 10784 2060
rect 10836 2048 10842 2100
rect 11882 2048 11888 2100
rect 11940 2088 11946 2100
rect 14918 2088 14924 2100
rect 11940 2060 14924 2088
rect 11940 2048 11946 2060
rect 14918 2048 14924 2060
rect 14976 2048 14982 2100
rect 16298 2088 16304 2100
rect 15028 2060 16304 2088
rect 3510 1980 3516 2032
rect 3568 2020 3574 2032
rect 6638 2020 6644 2032
rect 3568 1992 6644 2020
rect 3568 1980 3574 1992
rect 6638 1980 6644 1992
rect 6696 1980 6702 2032
rect 6730 1980 6736 2032
rect 6788 2020 6794 2032
rect 10226 2020 10232 2032
rect 6788 1992 10232 2020
rect 6788 1980 6794 1992
rect 10226 1980 10232 1992
rect 10284 1980 10290 2032
rect 13538 1980 13544 2032
rect 13596 2020 13602 2032
rect 15028 2020 15056 2060
rect 16298 2048 16304 2060
rect 16356 2048 16362 2100
rect 13596 1992 15056 2020
rect 13596 1980 13602 1992
rect 15378 1980 15384 2032
rect 15436 2020 15442 2032
rect 19150 2020 19156 2032
rect 15436 1992 19156 2020
rect 15436 1980 15442 1992
rect 19150 1980 19156 1992
rect 19208 1980 19214 2032
rect 4982 1912 4988 1964
rect 5040 1952 5046 1964
rect 7374 1952 7380 1964
rect 5040 1924 7380 1952
rect 5040 1912 5046 1924
rect 7374 1912 7380 1924
rect 7432 1912 7438 1964
rect 7742 1912 7748 1964
rect 7800 1952 7806 1964
rect 11698 1952 11704 1964
rect 7800 1924 11704 1952
rect 7800 1912 7806 1924
rect 11698 1912 11704 1924
rect 11756 1952 11762 1964
rect 12158 1952 12164 1964
rect 11756 1924 12164 1952
rect 11756 1912 11762 1924
rect 12158 1912 12164 1924
rect 12216 1912 12222 1964
rect 13262 1912 13268 1964
rect 13320 1952 13326 1964
rect 14274 1952 14280 1964
rect 13320 1924 14280 1952
rect 13320 1912 13326 1924
rect 14274 1912 14280 1924
rect 14332 1912 14338 1964
rect 14458 1912 14464 1964
rect 14516 1952 14522 1964
rect 19794 1952 19800 1964
rect 14516 1924 19800 1952
rect 14516 1912 14522 1924
rect 19794 1912 19800 1924
rect 19852 1912 19858 1964
rect 5626 1844 5632 1896
rect 5684 1884 5690 1896
rect 9398 1884 9404 1896
rect 5684 1856 9404 1884
rect 5684 1844 5690 1856
rect 9398 1844 9404 1856
rect 9456 1844 9462 1896
rect 9858 1844 9864 1896
rect 9916 1884 9922 1896
rect 15746 1884 15752 1896
rect 9916 1856 15752 1884
rect 9916 1844 9922 1856
rect 15746 1844 15752 1856
rect 15804 1844 15810 1896
rect 4338 1776 4344 1828
rect 4396 1816 4402 1828
rect 10870 1816 10876 1828
rect 4396 1788 10876 1816
rect 4396 1776 4402 1788
rect 10870 1776 10876 1788
rect 10928 1776 10934 1828
rect 14734 1776 14740 1828
rect 14792 1816 14798 1828
rect 15654 1816 15660 1828
rect 14792 1788 15660 1816
rect 14792 1776 14798 1788
rect 15654 1776 15660 1788
rect 15712 1776 15718 1828
rect 3786 1708 3792 1760
rect 3844 1748 3850 1760
rect 9766 1748 9772 1760
rect 3844 1720 9772 1748
rect 3844 1708 3850 1720
rect 9766 1708 9772 1720
rect 9824 1708 9830 1760
rect 2866 1640 2872 1692
rect 2924 1680 2930 1692
rect 8202 1680 8208 1692
rect 2924 1652 8208 1680
rect 2924 1640 2930 1652
rect 8202 1640 8208 1652
rect 8260 1680 8266 1692
rect 11790 1680 11796 1692
rect 8260 1652 11796 1680
rect 8260 1640 8266 1652
rect 11790 1640 11796 1652
rect 11848 1640 11854 1692
rect 7926 1572 7932 1624
rect 7984 1612 7990 1624
rect 9582 1612 9588 1624
rect 7984 1584 9588 1612
rect 7984 1572 7990 1584
rect 9582 1572 9588 1584
rect 9640 1572 9646 1624
rect 5810 1368 5816 1420
rect 5868 1408 5874 1420
rect 6270 1408 6276 1420
rect 5868 1380 6276 1408
rect 5868 1368 5874 1380
rect 6270 1368 6276 1380
rect 6328 1368 6334 1420
rect 16574 1368 16580 1420
rect 16632 1408 16638 1420
rect 17586 1408 17592 1420
rect 16632 1380 17592 1408
rect 16632 1368 16638 1380
rect 17586 1368 17592 1380
rect 17644 1368 17650 1420
rect 4614 1232 4620 1284
rect 4672 1272 4678 1284
rect 15562 1272 15568 1284
rect 4672 1244 15568 1272
rect 4672 1232 4678 1244
rect 15562 1232 15568 1244
rect 15620 1232 15626 1284
rect 842 1164 848 1216
rect 900 1204 906 1216
rect 11146 1204 11152 1216
rect 900 1176 11152 1204
rect 900 1164 906 1176
rect 11146 1164 11152 1176
rect 11204 1164 11210 1216
rect 1670 1096 1676 1148
rect 1728 1136 1734 1148
rect 13170 1136 13176 1148
rect 1728 1108 13176 1136
rect 1728 1096 1734 1108
rect 13170 1096 13176 1108
rect 13228 1096 13234 1148
<< via1 >>
rect 1032 21088 1084 21140
rect 11060 21088 11112 21140
rect 1676 21020 1728 21072
rect 17776 21020 17828 21072
rect 4528 20884 4580 20936
rect 11152 20884 11204 20936
rect 2136 20816 2188 20868
rect 17224 20816 17276 20868
rect 3976 20748 4028 20800
rect 6736 20748 6788 20800
rect 10048 20748 10100 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 1860 20587 1912 20596
rect 1860 20553 1869 20587
rect 1869 20553 1903 20587
rect 1903 20553 1912 20587
rect 1860 20544 1912 20553
rect 2228 20587 2280 20596
rect 2228 20553 2237 20587
rect 2237 20553 2271 20587
rect 2271 20553 2280 20587
rect 2228 20544 2280 20553
rect 3976 20476 4028 20528
rect 4344 20544 4396 20596
rect 5816 20544 5868 20596
rect 6828 20544 6880 20596
rect 10876 20544 10928 20596
rect 11704 20544 11756 20596
rect 11980 20544 12032 20596
rect 12440 20544 12492 20596
rect 12716 20544 12768 20596
rect 13084 20544 13136 20596
rect 13452 20544 13504 20596
rect 13820 20544 13872 20596
rect 14556 20544 14608 20596
rect 15200 20544 15252 20596
rect 15660 20544 15712 20596
rect 16580 20544 16632 20596
rect 16948 20544 17000 20596
rect 19524 20587 19576 20596
rect 5172 20476 5224 20528
rect 5264 20476 5316 20528
rect 6644 20476 6696 20528
rect 1676 20451 1728 20460
rect 1676 20417 1685 20451
rect 1685 20417 1719 20451
rect 1719 20417 1728 20451
rect 1676 20408 1728 20417
rect 2136 20408 2188 20460
rect 2412 20451 2464 20460
rect 2412 20417 2421 20451
rect 2421 20417 2455 20451
rect 2455 20417 2464 20451
rect 2412 20408 2464 20417
rect 3516 20451 3568 20460
rect 3516 20417 3525 20451
rect 3525 20417 3559 20451
rect 3559 20417 3568 20451
rect 3516 20408 3568 20417
rect 3608 20408 3660 20460
rect 4068 20408 4120 20460
rect 5080 20451 5132 20460
rect 4528 20340 4580 20392
rect 5080 20417 5089 20451
rect 5089 20417 5123 20451
rect 5123 20417 5132 20451
rect 5080 20408 5132 20417
rect 5356 20408 5408 20460
rect 5448 20340 5500 20392
rect 7288 20476 7340 20528
rect 7472 20476 7524 20528
rect 6828 20408 6880 20460
rect 7380 20408 7432 20460
rect 7656 20408 7708 20460
rect 8208 20408 8260 20460
rect 15752 20476 15804 20528
rect 9312 20408 9364 20460
rect 10140 20451 10192 20460
rect 2872 20272 2924 20324
rect 3976 20272 4028 20324
rect 4896 20315 4948 20324
rect 4896 20281 4905 20315
rect 4905 20281 4939 20315
rect 4939 20281 4948 20315
rect 4896 20272 4948 20281
rect 5356 20272 5408 20324
rect 6644 20340 6696 20392
rect 6828 20272 6880 20324
rect 1492 20247 1544 20256
rect 1492 20213 1501 20247
rect 1501 20213 1535 20247
rect 1535 20213 1544 20247
rect 1492 20204 1544 20213
rect 2780 20247 2832 20256
rect 2780 20213 2789 20247
rect 2789 20213 2823 20247
rect 2823 20213 2832 20247
rect 2780 20204 2832 20213
rect 2964 20204 3016 20256
rect 3424 20247 3476 20256
rect 3424 20213 3433 20247
rect 3433 20213 3467 20247
rect 3467 20213 3476 20247
rect 3424 20204 3476 20213
rect 5724 20204 5776 20256
rect 7104 20340 7156 20392
rect 8392 20204 8444 20256
rect 8484 20204 8536 20256
rect 8668 20340 8720 20392
rect 9128 20340 9180 20392
rect 9680 20383 9732 20392
rect 9680 20349 9689 20383
rect 9689 20349 9723 20383
rect 9723 20349 9732 20383
rect 9680 20340 9732 20349
rect 10140 20417 10149 20451
rect 10149 20417 10183 20451
rect 10183 20417 10192 20451
rect 10140 20408 10192 20417
rect 10508 20451 10560 20460
rect 10508 20417 10517 20451
rect 10517 20417 10551 20451
rect 10551 20417 10560 20451
rect 10508 20408 10560 20417
rect 10600 20408 10652 20460
rect 12072 20451 12124 20460
rect 12072 20417 12081 20451
rect 12081 20417 12115 20451
rect 12115 20417 12124 20451
rect 12072 20408 12124 20417
rect 12164 20408 12216 20460
rect 13084 20451 13136 20460
rect 13084 20417 13093 20451
rect 13093 20417 13127 20451
rect 13127 20417 13136 20451
rect 13084 20408 13136 20417
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 13176 20408 13228 20417
rect 13636 20408 13688 20460
rect 10968 20272 11020 20324
rect 13360 20340 13412 20392
rect 14280 20408 14332 20460
rect 14648 20408 14700 20460
rect 14924 20408 14976 20460
rect 15568 20451 15620 20460
rect 15568 20417 15577 20451
rect 15577 20417 15611 20451
rect 15611 20417 15620 20451
rect 15568 20408 15620 20417
rect 15936 20451 15988 20460
rect 15936 20417 15945 20451
rect 15945 20417 15979 20451
rect 15979 20417 15988 20451
rect 15936 20408 15988 20417
rect 11888 20204 11940 20256
rect 13544 20272 13596 20324
rect 14188 20272 14240 20324
rect 15292 20272 15344 20324
rect 17132 20476 17184 20528
rect 19524 20553 19533 20587
rect 19533 20553 19567 20587
rect 19567 20553 19576 20587
rect 19524 20544 19576 20553
rect 19984 20587 20036 20596
rect 19984 20553 19993 20587
rect 19993 20553 20027 20587
rect 20027 20553 20036 20587
rect 19984 20544 20036 20553
rect 20352 20587 20404 20596
rect 20352 20553 20361 20587
rect 20361 20553 20395 20587
rect 20395 20553 20404 20587
rect 20352 20544 20404 20553
rect 21180 20544 21232 20596
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 16948 20408 17000 20460
rect 17592 20408 17644 20460
rect 17960 20408 18012 20460
rect 18236 20408 18288 20460
rect 18696 20408 18748 20460
rect 13820 20204 13872 20256
rect 16396 20204 16448 20256
rect 17040 20272 17092 20324
rect 17868 20272 17920 20324
rect 18880 20272 18932 20324
rect 19708 20451 19760 20460
rect 19708 20417 19717 20451
rect 19717 20417 19751 20451
rect 19751 20417 19760 20451
rect 19708 20408 19760 20417
rect 20996 20408 21048 20460
rect 19616 20272 19668 20324
rect 17408 20204 17460 20256
rect 17500 20204 17552 20256
rect 18420 20204 18472 20256
rect 21364 20340 21416 20392
rect 21548 20272 21600 20324
rect 21088 20247 21140 20256
rect 21088 20213 21097 20247
rect 21097 20213 21131 20247
rect 21131 20213 21140 20247
rect 21088 20204 21140 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 1952 20000 2004 20052
rect 3884 20000 3936 20052
rect 2872 19975 2924 19984
rect 2872 19941 2881 19975
rect 2881 19941 2915 19975
rect 2915 19941 2924 19975
rect 2872 19932 2924 19941
rect 3240 19975 3292 19984
rect 3240 19941 3249 19975
rect 3249 19941 3283 19975
rect 3283 19941 3292 19975
rect 3240 19932 3292 19941
rect 3332 19932 3384 19984
rect 5540 20000 5592 20052
rect 6736 20000 6788 20052
rect 10600 20000 10652 20052
rect 11244 20000 11296 20052
rect 12072 20043 12124 20052
rect 12072 20009 12081 20043
rect 12081 20009 12115 20043
rect 12115 20009 12124 20043
rect 12072 20000 12124 20009
rect 13084 20043 13136 20052
rect 8392 19932 8444 19984
rect 8576 19932 8628 19984
rect 1768 19796 1820 19848
rect 2412 19839 2464 19848
rect 1400 19728 1452 19780
rect 2412 19805 2421 19839
rect 2421 19805 2455 19839
rect 2455 19805 2464 19839
rect 2412 19796 2464 19805
rect 2596 19796 2648 19848
rect 2228 19728 2280 19780
rect 3332 19728 3384 19780
rect 3608 19728 3660 19780
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 5724 19839 5776 19848
rect 5724 19805 5733 19839
rect 5733 19805 5767 19839
rect 5767 19805 5776 19839
rect 5724 19796 5776 19805
rect 4252 19660 4304 19712
rect 4712 19728 4764 19780
rect 5540 19728 5592 19780
rect 7748 19864 7800 19916
rect 8668 19864 8720 19916
rect 12440 19932 12492 19984
rect 13084 20009 13093 20043
rect 13093 20009 13127 20043
rect 13127 20009 13136 20043
rect 13084 20000 13136 20009
rect 13360 20043 13412 20052
rect 13360 20009 13369 20043
rect 13369 20009 13403 20043
rect 13403 20009 13412 20043
rect 13360 20000 13412 20009
rect 13636 20043 13688 20052
rect 13636 20009 13645 20043
rect 13645 20009 13679 20043
rect 13679 20009 13688 20043
rect 13636 20000 13688 20009
rect 14280 20043 14332 20052
rect 14280 20009 14289 20043
rect 14289 20009 14323 20043
rect 14323 20009 14332 20043
rect 14280 20000 14332 20009
rect 14648 20043 14700 20052
rect 14648 20009 14657 20043
rect 14657 20009 14691 20043
rect 14691 20009 14700 20043
rect 14648 20000 14700 20009
rect 14924 20043 14976 20052
rect 14924 20009 14933 20043
rect 14933 20009 14967 20043
rect 14967 20009 14976 20043
rect 14924 20000 14976 20009
rect 15568 20000 15620 20052
rect 15752 20043 15804 20052
rect 15752 20009 15761 20043
rect 15761 20009 15795 20043
rect 15795 20009 15804 20043
rect 15752 20000 15804 20009
rect 16672 20000 16724 20052
rect 17224 20000 17276 20052
rect 17408 20043 17460 20052
rect 17408 20009 17417 20043
rect 17417 20009 17451 20043
rect 17451 20009 17460 20043
rect 17408 20000 17460 20009
rect 18052 20000 18104 20052
rect 18236 20043 18288 20052
rect 18236 20009 18245 20043
rect 18245 20009 18279 20043
rect 18279 20009 18288 20043
rect 18236 20000 18288 20009
rect 18328 20000 18380 20052
rect 18512 20000 18564 20052
rect 18972 20000 19024 20052
rect 19340 20000 19392 20052
rect 20536 20043 20588 20052
rect 20536 20009 20545 20043
rect 20545 20009 20579 20043
rect 20579 20009 20588 20043
rect 20536 20000 20588 20009
rect 6920 19728 6972 19780
rect 8208 19728 8260 19780
rect 10324 19796 10376 19848
rect 12256 19864 12308 19916
rect 13176 19932 13228 19984
rect 13728 19975 13780 19984
rect 13728 19941 13737 19975
rect 13737 19941 13771 19975
rect 13771 19941 13780 19975
rect 13728 19932 13780 19941
rect 15936 19932 15988 19984
rect 16856 19932 16908 19984
rect 17776 19975 17828 19984
rect 17776 19941 17785 19975
rect 17785 19941 17819 19975
rect 17819 19941 17828 19975
rect 17776 19932 17828 19941
rect 18604 19932 18656 19984
rect 19248 19932 19300 19984
rect 9588 19728 9640 19780
rect 10416 19728 10468 19780
rect 5632 19703 5684 19712
rect 5632 19669 5641 19703
rect 5641 19669 5675 19703
rect 5675 19669 5684 19703
rect 5632 19660 5684 19669
rect 6092 19660 6144 19712
rect 7104 19660 7156 19712
rect 7196 19703 7248 19712
rect 7196 19669 7205 19703
rect 7205 19669 7239 19703
rect 7239 19669 7248 19703
rect 7196 19660 7248 19669
rect 7380 19660 7432 19712
rect 8116 19660 8168 19712
rect 8300 19703 8352 19712
rect 8300 19669 8309 19703
rect 8309 19669 8343 19703
rect 8343 19669 8352 19703
rect 8300 19660 8352 19669
rect 8760 19703 8812 19712
rect 8760 19669 8769 19703
rect 8769 19669 8803 19703
rect 8803 19669 8812 19703
rect 8760 19660 8812 19669
rect 8852 19660 8904 19712
rect 11612 19839 11664 19848
rect 10876 19728 10928 19780
rect 11612 19805 11621 19839
rect 11621 19805 11655 19839
rect 11655 19805 11664 19839
rect 11612 19796 11664 19805
rect 11888 19839 11940 19848
rect 11888 19805 11897 19839
rect 11897 19805 11931 19839
rect 11931 19805 11940 19839
rect 11888 19796 11940 19805
rect 12072 19796 12124 19848
rect 12900 19839 12952 19848
rect 12900 19805 12909 19839
rect 12909 19805 12943 19839
rect 12943 19805 12952 19839
rect 12900 19796 12952 19805
rect 13268 19796 13320 19848
rect 14096 19839 14148 19848
rect 12164 19728 12216 19780
rect 12808 19728 12860 19780
rect 11796 19703 11848 19712
rect 11796 19669 11805 19703
rect 11805 19669 11839 19703
rect 11839 19669 11848 19703
rect 11796 19660 11848 19669
rect 12624 19660 12676 19712
rect 14096 19805 14105 19839
rect 14105 19805 14139 19839
rect 14139 19805 14148 19839
rect 14096 19796 14148 19805
rect 14464 19839 14516 19848
rect 14464 19805 14473 19839
rect 14473 19805 14507 19839
rect 14507 19805 14516 19839
rect 14464 19796 14516 19805
rect 14740 19839 14792 19848
rect 14740 19805 14749 19839
rect 14749 19805 14783 19839
rect 14783 19805 14792 19839
rect 14740 19796 14792 19805
rect 15016 19839 15068 19848
rect 15016 19805 15025 19839
rect 15025 19805 15059 19839
rect 15059 19805 15068 19839
rect 15016 19796 15068 19805
rect 15200 19796 15252 19848
rect 15568 19839 15620 19848
rect 15568 19805 15577 19839
rect 15577 19805 15611 19839
rect 15611 19805 15620 19839
rect 15568 19796 15620 19805
rect 15752 19796 15804 19848
rect 18328 19864 18380 19916
rect 17316 19796 17368 19848
rect 17868 19796 17920 19848
rect 16304 19703 16356 19712
rect 16304 19669 16313 19703
rect 16313 19669 16347 19703
rect 16347 19669 16356 19703
rect 16304 19660 16356 19669
rect 17592 19728 17644 19780
rect 18144 19796 18196 19848
rect 19616 19864 19668 19916
rect 18788 19796 18840 19848
rect 18696 19728 18748 19780
rect 18972 19728 19024 19780
rect 19800 19796 19852 19848
rect 20444 19864 20496 19916
rect 20352 19839 20404 19848
rect 20352 19805 20361 19839
rect 20361 19805 20395 19839
rect 20395 19805 20404 19839
rect 20352 19796 20404 19805
rect 21272 19839 21324 19848
rect 21272 19805 21281 19839
rect 21281 19805 21315 19839
rect 21315 19805 21324 19839
rect 21272 19796 21324 19805
rect 19616 19728 19668 19780
rect 19892 19771 19944 19780
rect 19892 19737 19901 19771
rect 19901 19737 19935 19771
rect 19935 19737 19944 19771
rect 19892 19728 19944 19737
rect 20076 19728 20128 19780
rect 17500 19703 17552 19712
rect 17500 19669 17509 19703
rect 17509 19669 17543 19703
rect 17543 19669 17552 19703
rect 17500 19660 17552 19669
rect 18052 19660 18104 19712
rect 21456 19703 21508 19712
rect 21456 19669 21465 19703
rect 21465 19669 21499 19703
rect 21499 19669 21508 19703
rect 21456 19660 21508 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 1584 19456 1636 19508
rect 2872 19456 2924 19508
rect 3332 19456 3384 19508
rect 112 19388 164 19440
rect 940 19388 992 19440
rect 204 19320 256 19372
rect 1308 19320 1360 19372
rect 1676 19363 1728 19372
rect 1676 19329 1685 19363
rect 1685 19329 1719 19363
rect 1719 19329 1728 19363
rect 1676 19320 1728 19329
rect 1952 19320 2004 19372
rect 3148 19388 3200 19440
rect 3792 19456 3844 19508
rect 5264 19456 5316 19508
rect 6000 19456 6052 19508
rect 7196 19456 7248 19508
rect 8668 19499 8720 19508
rect 8668 19465 8677 19499
rect 8677 19465 8711 19499
rect 8711 19465 8720 19499
rect 8668 19456 8720 19465
rect 8760 19456 8812 19508
rect 10600 19456 10652 19508
rect 12072 19456 12124 19508
rect 12440 19456 12492 19508
rect 12532 19456 12584 19508
rect 14096 19456 14148 19508
rect 15016 19456 15068 19508
rect 16948 19456 17000 19508
rect 17960 19456 18012 19508
rect 18420 19499 18472 19508
rect 2964 19320 3016 19372
rect 4344 19363 4396 19372
rect 3332 19252 3384 19304
rect 3700 19252 3752 19304
rect 3884 19295 3936 19304
rect 3884 19261 3893 19295
rect 3893 19261 3927 19295
rect 3927 19261 3936 19295
rect 3884 19252 3936 19261
rect 4344 19329 4353 19363
rect 4353 19329 4387 19363
rect 4387 19329 4396 19363
rect 4344 19320 4396 19329
rect 4436 19320 4488 19372
rect 4620 19252 4672 19304
rect 5540 19295 5592 19304
rect 5540 19261 5549 19295
rect 5549 19261 5583 19295
rect 5583 19261 5592 19295
rect 5540 19252 5592 19261
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 3148 19159 3200 19168
rect 3148 19125 3157 19159
rect 3157 19125 3191 19159
rect 3191 19125 3200 19159
rect 3148 19116 3200 19125
rect 3240 19159 3292 19168
rect 3240 19125 3249 19159
rect 3249 19125 3283 19159
rect 3283 19125 3292 19159
rect 3240 19116 3292 19125
rect 4252 19116 4304 19168
rect 5632 19184 5684 19236
rect 6276 19116 6328 19168
rect 7196 19320 7248 19372
rect 7104 19184 7156 19236
rect 7288 19295 7340 19346
rect 7564 19363 7616 19372
rect 7564 19329 7598 19363
rect 7598 19329 7616 19363
rect 10232 19388 10284 19440
rect 7564 19320 7616 19329
rect 8852 19320 8904 19372
rect 9772 19320 9824 19372
rect 11612 19320 11664 19372
rect 12256 19388 12308 19440
rect 12900 19388 12952 19440
rect 14740 19388 14792 19440
rect 14924 19431 14976 19440
rect 14924 19397 14933 19431
rect 14933 19397 14967 19431
rect 14967 19397 14976 19431
rect 14924 19388 14976 19397
rect 16396 19388 16448 19440
rect 12072 19320 12124 19372
rect 7288 19294 7297 19295
rect 7297 19294 7331 19295
rect 7331 19294 7340 19295
rect 10416 19295 10468 19304
rect 10416 19261 10425 19295
rect 10425 19261 10459 19295
rect 10459 19261 10468 19295
rect 10416 19252 10468 19261
rect 13084 19252 13136 19304
rect 14372 19320 14424 19372
rect 14556 19320 14608 19372
rect 15568 19320 15620 19372
rect 16120 19320 16172 19372
rect 16856 19320 16908 19372
rect 17316 19388 17368 19440
rect 18420 19465 18429 19499
rect 18429 19465 18463 19499
rect 18463 19465 18472 19499
rect 18420 19456 18472 19465
rect 18788 19499 18840 19508
rect 18788 19465 18797 19499
rect 18797 19465 18831 19499
rect 18831 19465 18840 19499
rect 18788 19456 18840 19465
rect 18972 19456 19024 19508
rect 19432 19456 19484 19508
rect 22284 19456 22336 19508
rect 17960 19363 18012 19372
rect 17960 19329 17969 19363
rect 17969 19329 18003 19363
rect 18003 19329 18012 19363
rect 17960 19320 18012 19329
rect 18236 19363 18288 19372
rect 18236 19329 18245 19363
rect 18245 19329 18279 19363
rect 18279 19329 18288 19363
rect 18236 19320 18288 19329
rect 18328 19320 18380 19372
rect 18696 19320 18748 19372
rect 19248 19363 19300 19372
rect 19248 19329 19257 19363
rect 19257 19329 19291 19363
rect 19291 19329 19300 19363
rect 19248 19320 19300 19329
rect 19340 19363 19392 19372
rect 19340 19329 19349 19363
rect 19349 19329 19383 19363
rect 19383 19329 19392 19363
rect 19340 19320 19392 19329
rect 19524 19320 19576 19372
rect 19984 19363 20036 19372
rect 19984 19329 19993 19363
rect 19993 19329 20027 19363
rect 20027 19329 20036 19363
rect 19984 19320 20036 19329
rect 20444 19320 20496 19372
rect 20628 19320 20680 19372
rect 21180 19320 21232 19372
rect 20812 19252 20864 19304
rect 7564 19116 7616 19168
rect 9680 19116 9732 19168
rect 11244 19159 11296 19168
rect 11244 19125 11253 19159
rect 11253 19125 11287 19159
rect 11287 19125 11296 19159
rect 11244 19116 11296 19125
rect 15292 19227 15344 19236
rect 15292 19193 15301 19227
rect 15301 19193 15335 19227
rect 15335 19193 15344 19227
rect 15292 19184 15344 19193
rect 18880 19184 18932 19236
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 12900 19116 12952 19125
rect 13176 19116 13228 19168
rect 13360 19116 13412 19168
rect 13728 19116 13780 19168
rect 14096 19116 14148 19168
rect 14464 19116 14516 19168
rect 15016 19116 15068 19168
rect 15200 19159 15252 19168
rect 15200 19125 15209 19159
rect 15209 19125 15243 19159
rect 15243 19125 15252 19159
rect 15200 19116 15252 19125
rect 15476 19159 15528 19168
rect 15476 19125 15485 19159
rect 15485 19125 15519 19159
rect 15519 19125 15528 19159
rect 15476 19116 15528 19125
rect 15660 19159 15712 19168
rect 15660 19125 15669 19159
rect 15669 19125 15703 19159
rect 15703 19125 15712 19159
rect 15660 19116 15712 19125
rect 16120 19159 16172 19168
rect 16120 19125 16129 19159
rect 16129 19125 16163 19159
rect 16163 19125 16172 19159
rect 16120 19116 16172 19125
rect 16396 19116 16448 19168
rect 16856 19159 16908 19168
rect 16856 19125 16865 19159
rect 16865 19125 16899 19159
rect 16899 19125 16908 19159
rect 16856 19116 16908 19125
rect 18328 19116 18380 19168
rect 20260 19184 20312 19236
rect 20536 19227 20588 19236
rect 20536 19193 20545 19227
rect 20545 19193 20579 19227
rect 20579 19193 20588 19227
rect 20536 19184 20588 19193
rect 19892 19116 19944 19168
rect 20168 19116 20220 19168
rect 21456 19159 21508 19168
rect 21456 19125 21465 19159
rect 21465 19125 21499 19159
rect 21499 19125 21508 19159
rect 21456 19116 21508 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 1676 18912 1728 18964
rect 2504 18912 2556 18964
rect 2688 18912 2740 18964
rect 2872 18912 2924 18964
rect 5448 18912 5500 18964
rect 5908 18912 5960 18964
rect 1768 18844 1820 18896
rect 2964 18844 3016 18896
rect 3148 18776 3200 18828
rect 3700 18776 3752 18828
rect 5724 18844 5776 18896
rect 7564 18912 7616 18964
rect 9772 18912 9824 18964
rect 10232 18955 10284 18964
rect 10232 18921 10241 18955
rect 10241 18921 10275 18955
rect 10275 18921 10284 18955
rect 10232 18912 10284 18921
rect 10876 18912 10928 18964
rect 10968 18912 11020 18964
rect 1676 18751 1728 18760
rect 1676 18717 1685 18751
rect 1685 18717 1719 18751
rect 1719 18717 1728 18751
rect 1676 18708 1728 18717
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 2596 18751 2648 18760
rect 2596 18717 2605 18751
rect 2605 18717 2639 18751
rect 2639 18717 2648 18751
rect 2596 18708 2648 18717
rect 3240 18751 3292 18760
rect 3240 18717 3249 18751
rect 3249 18717 3283 18751
rect 3283 18717 3292 18751
rect 3240 18708 3292 18717
rect 6000 18708 6052 18760
rect 2504 18640 2556 18692
rect 5908 18640 5960 18692
rect 7748 18776 7800 18828
rect 8668 18776 8720 18828
rect 6736 18751 6788 18760
rect 6736 18717 6770 18751
rect 6770 18717 6788 18751
rect 6736 18708 6788 18717
rect 6276 18640 6328 18692
rect 8300 18708 8352 18760
rect 9404 18708 9456 18760
rect 7012 18640 7064 18692
rect 9772 18683 9824 18692
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 2872 18615 2924 18624
rect 2872 18581 2881 18615
rect 2881 18581 2915 18615
rect 2915 18581 2924 18615
rect 2872 18572 2924 18581
rect 3332 18572 3384 18624
rect 4068 18572 4120 18624
rect 4712 18572 4764 18624
rect 5632 18615 5684 18624
rect 5632 18581 5641 18615
rect 5641 18581 5675 18615
rect 5675 18581 5684 18615
rect 5632 18572 5684 18581
rect 5816 18572 5868 18624
rect 7932 18615 7984 18624
rect 7932 18581 7941 18615
rect 7941 18581 7975 18615
rect 7975 18581 7984 18615
rect 8300 18615 8352 18624
rect 7932 18572 7984 18581
rect 8300 18581 8309 18615
rect 8309 18581 8343 18615
rect 8343 18581 8352 18615
rect 8300 18572 8352 18581
rect 9036 18572 9088 18624
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9772 18649 9781 18683
rect 9781 18649 9815 18683
rect 9815 18649 9824 18683
rect 9772 18640 9824 18649
rect 12072 18776 12124 18828
rect 18604 18912 18656 18964
rect 19616 18955 19668 18964
rect 19616 18921 19625 18955
rect 19625 18921 19659 18955
rect 19659 18921 19668 18955
rect 19616 18912 19668 18921
rect 20996 18912 21048 18964
rect 12348 18844 12400 18896
rect 12532 18844 12584 18896
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 10692 18708 10744 18760
rect 13360 18776 13412 18828
rect 14280 18819 14332 18828
rect 12440 18708 12492 18760
rect 12900 18708 12952 18760
rect 14280 18785 14289 18819
rect 14289 18785 14323 18819
rect 14323 18785 14332 18819
rect 14280 18776 14332 18785
rect 19432 18844 19484 18896
rect 13820 18708 13872 18760
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 19340 18776 19392 18828
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 19432 18708 19484 18717
rect 19708 18844 19760 18896
rect 20536 18844 20588 18896
rect 20444 18751 20496 18760
rect 9312 18572 9364 18581
rect 10508 18572 10560 18624
rect 10692 18572 10744 18624
rect 11612 18640 11664 18692
rect 11980 18640 12032 18692
rect 12348 18572 12400 18624
rect 12624 18572 12676 18624
rect 13452 18640 13504 18692
rect 13268 18615 13320 18624
rect 13268 18581 13277 18615
rect 13277 18581 13311 18615
rect 13311 18581 13320 18615
rect 13268 18572 13320 18581
rect 14832 18615 14884 18624
rect 14832 18581 14841 18615
rect 14841 18581 14875 18615
rect 14875 18581 14884 18615
rect 14832 18572 14884 18581
rect 19340 18572 19392 18624
rect 19524 18572 19576 18624
rect 20444 18717 20453 18751
rect 20453 18717 20487 18751
rect 20487 18717 20496 18751
rect 20444 18708 20496 18717
rect 20628 18751 20680 18760
rect 20628 18717 20637 18751
rect 20637 18717 20671 18751
rect 20671 18717 20680 18751
rect 20628 18708 20680 18717
rect 20260 18640 20312 18692
rect 20904 18683 20956 18692
rect 20904 18649 20913 18683
rect 20913 18649 20947 18683
rect 20947 18649 20956 18683
rect 20904 18640 20956 18649
rect 20352 18572 20404 18624
rect 21456 18615 21508 18624
rect 21456 18581 21465 18615
rect 21465 18581 21499 18615
rect 21499 18581 21508 18615
rect 21456 18572 21508 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 1768 18411 1820 18420
rect 1768 18377 1777 18411
rect 1777 18377 1811 18411
rect 1811 18377 1820 18411
rect 1768 18368 1820 18377
rect 5632 18368 5684 18420
rect 6000 18368 6052 18420
rect 1216 18300 1268 18352
rect 2780 18300 2832 18352
rect 2964 18300 3016 18352
rect 3332 18300 3384 18352
rect 5080 18300 5132 18352
rect 7288 18368 7340 18420
rect 7932 18368 7984 18420
rect 8208 18411 8260 18420
rect 8208 18377 8217 18411
rect 8217 18377 8251 18411
rect 8251 18377 8260 18411
rect 8208 18368 8260 18377
rect 9404 18368 9456 18420
rect 6552 18300 6604 18352
rect 12624 18411 12676 18420
rect 1768 18232 1820 18284
rect 1952 18275 2004 18284
rect 1952 18241 1961 18275
rect 1961 18241 1995 18275
rect 1995 18241 2004 18275
rect 1952 18232 2004 18241
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 2136 18028 2188 18080
rect 3240 18028 3292 18080
rect 3700 18232 3752 18284
rect 3884 18275 3936 18284
rect 3884 18241 3893 18275
rect 3893 18241 3927 18275
rect 3927 18241 3936 18275
rect 3884 18232 3936 18241
rect 3976 18232 4028 18284
rect 4988 18275 5040 18284
rect 4988 18241 4997 18275
rect 4997 18241 5031 18275
rect 5031 18241 5040 18275
rect 4988 18232 5040 18241
rect 5448 18232 5500 18284
rect 6368 18232 6420 18284
rect 3516 18164 3568 18216
rect 4712 18207 4764 18216
rect 4712 18173 4721 18207
rect 4721 18173 4755 18207
rect 4755 18173 4764 18207
rect 4712 18164 4764 18173
rect 5540 18164 5592 18216
rect 6092 18164 6144 18216
rect 7012 18232 7064 18284
rect 7196 18275 7248 18284
rect 7196 18241 7205 18275
rect 7205 18241 7239 18275
rect 7239 18241 7248 18275
rect 7196 18232 7248 18241
rect 5448 18096 5500 18148
rect 6736 18096 6788 18148
rect 4528 18071 4580 18080
rect 4528 18037 4537 18071
rect 4537 18037 4571 18071
rect 4571 18037 4580 18071
rect 4528 18028 4580 18037
rect 4620 18028 4672 18080
rect 4896 18028 4948 18080
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 7932 18232 7984 18284
rect 9496 18275 9548 18284
rect 9496 18241 9505 18275
rect 9505 18241 9539 18275
rect 9539 18241 9548 18275
rect 9496 18232 9548 18241
rect 7564 18207 7616 18216
rect 7564 18173 7573 18207
rect 7573 18173 7607 18207
rect 7607 18173 7616 18207
rect 7564 18164 7616 18173
rect 8300 18164 8352 18216
rect 8576 18207 8628 18216
rect 8576 18173 8585 18207
rect 8585 18173 8619 18207
rect 8619 18173 8628 18207
rect 8576 18164 8628 18173
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 10784 18232 10836 18284
rect 10692 18207 10744 18216
rect 9036 18139 9088 18148
rect 9036 18105 9045 18139
rect 9045 18105 9079 18139
rect 9079 18105 9088 18139
rect 9036 18096 9088 18105
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 10876 18207 10928 18216
rect 10876 18173 10885 18207
rect 10885 18173 10919 18207
rect 10919 18173 10928 18207
rect 10876 18164 10928 18173
rect 11796 18300 11848 18352
rect 12624 18377 12633 18411
rect 12633 18377 12667 18411
rect 12667 18377 12676 18411
rect 12624 18368 12676 18377
rect 13268 18368 13320 18420
rect 17960 18368 18012 18420
rect 19524 18368 19576 18420
rect 21640 18368 21692 18420
rect 11612 18232 11664 18284
rect 12900 18300 12952 18352
rect 16396 18300 16448 18352
rect 14556 18232 14608 18284
rect 20812 18300 20864 18352
rect 19708 18275 19760 18284
rect 19708 18241 19717 18275
rect 19717 18241 19751 18275
rect 19751 18241 19760 18275
rect 19708 18232 19760 18241
rect 20168 18232 20220 18284
rect 20352 18275 20404 18284
rect 20352 18241 20361 18275
rect 20361 18241 20395 18275
rect 20395 18241 20404 18275
rect 20352 18232 20404 18241
rect 20536 18232 20588 18284
rect 20720 18232 20772 18284
rect 20996 18232 21048 18284
rect 11980 18207 12032 18216
rect 11980 18173 11989 18207
rect 11989 18173 12023 18207
rect 12023 18173 12032 18207
rect 11980 18164 12032 18173
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 12716 18207 12768 18216
rect 12716 18173 12725 18207
rect 12725 18173 12759 18207
rect 12759 18173 12768 18207
rect 12716 18164 12768 18173
rect 13084 18207 13136 18216
rect 13084 18173 13093 18207
rect 13093 18173 13127 18207
rect 13127 18173 13136 18207
rect 13084 18164 13136 18173
rect 19340 18164 19392 18216
rect 20444 18164 20496 18216
rect 7748 18028 7800 18080
rect 9864 18096 9916 18148
rect 12532 18096 12584 18148
rect 9680 18028 9732 18080
rect 11060 18028 11112 18080
rect 11612 18028 11664 18080
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 20628 18096 20680 18148
rect 11704 18028 11756 18037
rect 14280 18028 14332 18080
rect 14464 18071 14516 18080
rect 14464 18037 14473 18071
rect 14473 18037 14507 18071
rect 14507 18037 14516 18071
rect 14464 18028 14516 18037
rect 15016 18028 15068 18080
rect 16028 18028 16080 18080
rect 19616 18028 19668 18080
rect 19984 18028 20036 18080
rect 20168 18071 20220 18080
rect 20168 18037 20177 18071
rect 20177 18037 20211 18071
rect 20211 18037 20220 18071
rect 20168 18028 20220 18037
rect 21364 18164 21416 18216
rect 21088 18139 21140 18148
rect 21088 18105 21097 18139
rect 21097 18105 21131 18139
rect 21131 18105 21140 18139
rect 21088 18096 21140 18105
rect 21180 18028 21232 18080
rect 21456 18071 21508 18080
rect 21456 18037 21465 18071
rect 21465 18037 21499 18071
rect 21499 18037 21508 18071
rect 21456 18028 21508 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 1676 17824 1728 17876
rect 2412 17824 2464 17876
rect 1676 17663 1728 17672
rect 1676 17629 1685 17663
rect 1685 17629 1719 17663
rect 1719 17629 1728 17663
rect 1676 17620 1728 17629
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 3240 17620 3292 17672
rect 2136 17552 2188 17604
rect 3056 17552 3108 17604
rect 3424 17824 3476 17876
rect 3516 17620 3568 17672
rect 4436 17824 4488 17876
rect 5080 17824 5132 17876
rect 5908 17824 5960 17876
rect 6644 17824 6696 17876
rect 7748 17824 7800 17876
rect 9312 17824 9364 17876
rect 4436 17688 4488 17740
rect 6368 17756 6420 17808
rect 4252 17620 4304 17672
rect 6552 17688 6604 17740
rect 8116 17688 8168 17740
rect 8300 17688 8352 17740
rect 10140 17867 10192 17876
rect 10140 17833 10149 17867
rect 10149 17833 10183 17867
rect 10183 17833 10192 17867
rect 10416 17867 10468 17876
rect 10140 17824 10192 17833
rect 10416 17833 10425 17867
rect 10425 17833 10459 17867
rect 10459 17833 10468 17867
rect 10416 17824 10468 17833
rect 11060 17867 11112 17876
rect 11060 17833 11069 17867
rect 11069 17833 11103 17867
rect 11103 17833 11112 17867
rect 11060 17824 11112 17833
rect 12164 17824 12216 17876
rect 12348 17824 12400 17876
rect 16304 17824 16356 17876
rect 19064 17824 19116 17876
rect 21272 17824 21324 17876
rect 9680 17688 9732 17740
rect 9864 17688 9916 17740
rect 5264 17620 5316 17672
rect 5448 17620 5500 17672
rect 10232 17756 10284 17808
rect 12900 17756 12952 17808
rect 19708 17756 19760 17808
rect 10048 17688 10100 17740
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 11244 17688 11296 17740
rect 11520 17731 11572 17740
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 12164 17688 12216 17740
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 18880 17688 18932 17740
rect 22100 17756 22152 17808
rect 13728 17620 13780 17672
rect 14188 17663 14240 17672
rect 14188 17629 14197 17663
rect 14197 17629 14231 17663
rect 14231 17629 14240 17663
rect 14188 17620 14240 17629
rect 14464 17663 14516 17672
rect 14464 17629 14498 17663
rect 14498 17629 14516 17663
rect 14464 17620 14516 17629
rect 17408 17620 17460 17672
rect 19708 17663 19760 17672
rect 19708 17629 19717 17663
rect 19717 17629 19751 17663
rect 19751 17629 19760 17663
rect 19708 17620 19760 17629
rect 20076 17663 20128 17672
rect 20076 17629 20085 17663
rect 20085 17629 20119 17663
rect 20119 17629 20128 17663
rect 20076 17620 20128 17629
rect 21272 17663 21324 17672
rect 2596 17484 2648 17536
rect 2780 17484 2832 17536
rect 3148 17484 3200 17536
rect 4068 17484 4120 17536
rect 4528 17484 4580 17536
rect 5540 17552 5592 17604
rect 5908 17552 5960 17604
rect 6092 17484 6144 17536
rect 6460 17552 6512 17604
rect 7012 17552 7064 17604
rect 6644 17527 6696 17536
rect 6644 17493 6653 17527
rect 6653 17493 6687 17527
rect 6687 17493 6696 17527
rect 6644 17484 6696 17493
rect 7104 17484 7156 17536
rect 7932 17527 7984 17536
rect 7932 17493 7941 17527
rect 7941 17493 7975 17527
rect 7975 17493 7984 17527
rect 7932 17484 7984 17493
rect 8208 17484 8260 17536
rect 8392 17527 8444 17536
rect 8392 17493 8401 17527
rect 8401 17493 8435 17527
rect 8435 17493 8444 17527
rect 8392 17484 8444 17493
rect 8760 17484 8812 17536
rect 9496 17484 9548 17536
rect 10140 17484 10192 17536
rect 13452 17595 13504 17604
rect 13452 17561 13461 17595
rect 13461 17561 13495 17595
rect 13495 17561 13504 17595
rect 13452 17552 13504 17561
rect 13636 17552 13688 17604
rect 19524 17552 19576 17604
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 10692 17527 10744 17536
rect 10692 17493 10701 17527
rect 10701 17493 10735 17527
rect 10735 17493 10744 17527
rect 10692 17484 10744 17493
rect 10876 17527 10928 17536
rect 10876 17493 10885 17527
rect 10885 17493 10919 17527
rect 10919 17493 10928 17527
rect 10876 17484 10928 17493
rect 11796 17527 11848 17536
rect 11796 17493 11805 17527
rect 11805 17493 11839 17527
rect 11839 17493 11848 17527
rect 11796 17484 11848 17493
rect 12440 17484 12492 17536
rect 12532 17484 12584 17536
rect 13728 17484 13780 17536
rect 14740 17484 14792 17536
rect 15200 17484 15252 17536
rect 15292 17484 15344 17536
rect 15660 17527 15712 17536
rect 15660 17493 15669 17527
rect 15669 17493 15703 17527
rect 15703 17493 15712 17527
rect 16028 17527 16080 17536
rect 15660 17484 15712 17493
rect 16028 17493 16037 17527
rect 16037 17493 16071 17527
rect 16071 17493 16080 17527
rect 16028 17484 16080 17493
rect 17868 17484 17920 17536
rect 20352 17527 20404 17536
rect 20352 17493 20361 17527
rect 20361 17493 20395 17527
rect 20395 17493 20404 17527
rect 20352 17484 20404 17493
rect 21456 17527 21508 17536
rect 21456 17493 21465 17527
rect 21465 17493 21499 17527
rect 21499 17493 21508 17527
rect 21456 17484 21508 17493
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1768 17280 1820 17332
rect 1952 17280 2004 17332
rect 2872 17280 2924 17332
rect 3332 17280 3384 17332
rect 3424 17212 3476 17264
rect 4436 17212 4488 17264
rect 4988 17280 5040 17332
rect 5908 17323 5960 17332
rect 5908 17289 5917 17323
rect 5917 17289 5951 17323
rect 5951 17289 5960 17323
rect 5908 17280 5960 17289
rect 6184 17280 6236 17332
rect 8208 17323 8260 17332
rect 8208 17289 8217 17323
rect 8217 17289 8251 17323
rect 8251 17289 8260 17323
rect 8208 17280 8260 17289
rect 8576 17280 8628 17332
rect 10140 17280 10192 17332
rect 10692 17280 10744 17332
rect 10784 17280 10836 17332
rect 12716 17280 12768 17332
rect 12992 17323 13044 17332
rect 12992 17289 13001 17323
rect 13001 17289 13035 17323
rect 13035 17289 13044 17323
rect 12992 17280 13044 17289
rect 14832 17280 14884 17332
rect 20260 17280 20312 17332
rect 20536 17280 20588 17332
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 20996 17323 21048 17332
rect 20996 17289 21005 17323
rect 21005 17289 21039 17323
rect 21039 17289 21048 17323
rect 20996 17280 21048 17289
rect 7656 17255 7708 17264
rect 7656 17221 7665 17255
rect 7665 17221 7699 17255
rect 7699 17221 7708 17255
rect 7656 17212 7708 17221
rect 8116 17212 8168 17264
rect 1768 17144 1820 17196
rect 2136 17144 2188 17196
rect 3148 17144 3200 17196
rect 3240 17187 3292 17196
rect 3240 17153 3249 17187
rect 3249 17153 3283 17187
rect 3283 17153 3292 17187
rect 3240 17144 3292 17153
rect 4068 17144 4120 17196
rect 2228 17076 2280 17128
rect 3056 17076 3108 17128
rect 5356 17187 5408 17196
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 5908 17144 5960 17196
rect 7564 17144 7616 17196
rect 7840 17144 7892 17196
rect 8668 17187 8720 17196
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 9404 17187 9456 17196
rect 8668 17144 8720 17153
rect 9404 17153 9413 17187
rect 9413 17153 9447 17187
rect 9447 17153 9456 17187
rect 9404 17144 9456 17153
rect 10232 17212 10284 17264
rect 15568 17212 15620 17264
rect 19708 17212 19760 17264
rect 11980 17144 12032 17196
rect 6000 17119 6052 17128
rect 6000 17085 6009 17119
rect 6009 17085 6043 17119
rect 6043 17085 6052 17119
rect 6000 17076 6052 17085
rect 4896 17051 4948 17060
rect 4896 17017 4905 17051
rect 4905 17017 4939 17051
rect 4939 17017 4948 17051
rect 4896 17008 4948 17017
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 1860 16940 1912 16992
rect 4804 16940 4856 16992
rect 5080 16940 5132 16992
rect 5264 17008 5316 17060
rect 7104 17076 7156 17128
rect 6736 17008 6788 17060
rect 7656 17076 7708 17128
rect 8300 17008 8352 17060
rect 9680 17076 9732 17128
rect 9772 17076 9824 17128
rect 7840 16940 7892 16992
rect 10600 16940 10652 16992
rect 13636 17144 13688 17196
rect 14188 17144 14240 17196
rect 14464 17144 14516 17196
rect 15844 17187 15896 17196
rect 11244 17051 11296 17060
rect 11244 17017 11253 17051
rect 11253 17017 11287 17051
rect 11287 17017 11296 17051
rect 11244 17008 11296 17017
rect 11704 17008 11756 17060
rect 12532 17076 12584 17128
rect 13820 17076 13872 17128
rect 15108 17119 15160 17128
rect 15108 17085 15117 17119
rect 15117 17085 15151 17119
rect 15151 17085 15160 17119
rect 15108 17076 15160 17085
rect 15200 17119 15252 17128
rect 15200 17085 15209 17119
rect 15209 17085 15243 17119
rect 15243 17085 15252 17119
rect 15200 17076 15252 17085
rect 15844 17153 15853 17187
rect 15853 17153 15887 17187
rect 15887 17153 15896 17187
rect 15844 17144 15896 17153
rect 19800 17187 19852 17196
rect 19800 17153 19809 17187
rect 19809 17153 19843 17187
rect 19843 17153 19852 17187
rect 19800 17144 19852 17153
rect 20536 17187 20588 17196
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 20812 17187 20864 17196
rect 20812 17153 20821 17187
rect 20821 17153 20855 17187
rect 20855 17153 20864 17187
rect 20812 17144 20864 17153
rect 14372 17008 14424 17060
rect 15292 17008 15344 17060
rect 16948 17076 17000 17128
rect 20444 17076 20496 17128
rect 11980 16940 12032 16992
rect 12164 16940 12216 16992
rect 12624 16940 12676 16992
rect 13360 16940 13412 16992
rect 13728 16940 13780 16992
rect 20628 17008 20680 17060
rect 20812 17008 20864 17060
rect 22836 17008 22888 17060
rect 16028 16940 16080 16992
rect 19892 16940 19944 16992
rect 20536 16940 20588 16992
rect 21456 16983 21508 16992
rect 21456 16949 21465 16983
rect 21465 16949 21499 16983
rect 21499 16949 21508 16983
rect 21456 16940 21508 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1676 16736 1728 16788
rect 2780 16779 2832 16788
rect 2780 16745 2789 16779
rect 2789 16745 2823 16779
rect 2823 16745 2832 16779
rect 2780 16736 2832 16745
rect 2504 16668 2556 16720
rect 4528 16736 4580 16788
rect 4804 16736 4856 16788
rect 6644 16779 6696 16788
rect 6644 16745 6653 16779
rect 6653 16745 6687 16779
rect 6687 16745 6696 16779
rect 6644 16736 6696 16745
rect 7196 16736 7248 16788
rect 7748 16736 7800 16788
rect 8392 16736 8444 16788
rect 9680 16736 9732 16788
rect 11060 16736 11112 16788
rect 12348 16736 12400 16788
rect 2872 16600 2924 16652
rect 1676 16575 1728 16584
rect 1676 16541 1685 16575
rect 1685 16541 1719 16575
rect 1719 16541 1728 16575
rect 1676 16532 1728 16541
rect 2228 16532 2280 16584
rect 2596 16575 2648 16584
rect 2596 16541 2605 16575
rect 2605 16541 2639 16575
rect 2639 16541 2648 16575
rect 2596 16532 2648 16541
rect 3976 16532 4028 16584
rect 1400 16464 1452 16516
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 1860 16439 1912 16448
rect 1860 16405 1869 16439
rect 1869 16405 1903 16439
rect 1903 16405 1912 16439
rect 1860 16396 1912 16405
rect 2504 16464 2556 16516
rect 2964 16464 3016 16516
rect 5632 16600 5684 16652
rect 6552 16600 6604 16652
rect 7564 16643 7616 16652
rect 4252 16532 4304 16584
rect 4436 16575 4488 16584
rect 4436 16541 4470 16575
rect 4470 16541 4488 16575
rect 4436 16532 4488 16541
rect 4712 16532 4764 16584
rect 3332 16396 3384 16448
rect 4988 16464 5040 16516
rect 6184 16575 6236 16584
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 7564 16609 7573 16643
rect 7573 16609 7607 16643
rect 7607 16609 7616 16643
rect 7564 16600 7616 16609
rect 10416 16668 10468 16720
rect 12440 16668 12492 16720
rect 8576 16600 8628 16652
rect 9036 16600 9088 16652
rect 9404 16600 9456 16652
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 11704 16643 11756 16652
rect 11704 16609 11713 16643
rect 11713 16609 11747 16643
rect 11747 16609 11756 16643
rect 11704 16600 11756 16609
rect 14464 16736 14516 16788
rect 15568 16779 15620 16788
rect 15568 16745 15577 16779
rect 15577 16745 15611 16779
rect 15611 16745 15620 16779
rect 15568 16736 15620 16745
rect 15844 16736 15896 16788
rect 16488 16736 16540 16788
rect 18788 16736 18840 16788
rect 19800 16736 19852 16788
rect 21272 16736 21324 16788
rect 18236 16711 18288 16720
rect 6184 16532 6236 16541
rect 7656 16532 7708 16584
rect 10048 16532 10100 16584
rect 13360 16532 13412 16584
rect 16028 16643 16080 16652
rect 16028 16609 16037 16643
rect 16037 16609 16071 16643
rect 16071 16609 16080 16643
rect 16028 16600 16080 16609
rect 4436 16396 4488 16448
rect 5816 16439 5868 16448
rect 5816 16405 5825 16439
rect 5825 16405 5859 16439
rect 5859 16405 5868 16439
rect 5816 16396 5868 16405
rect 6828 16396 6880 16448
rect 7012 16439 7064 16448
rect 7012 16405 7021 16439
rect 7021 16405 7055 16439
rect 7055 16405 7064 16439
rect 7012 16396 7064 16405
rect 7196 16396 7248 16448
rect 7380 16396 7432 16448
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 8576 16396 8628 16448
rect 9312 16396 9364 16448
rect 9588 16396 9640 16448
rect 9864 16439 9916 16448
rect 9864 16405 9873 16439
rect 9873 16405 9907 16439
rect 9907 16405 9916 16439
rect 11244 16464 11296 16516
rect 9864 16396 9916 16405
rect 10324 16439 10376 16448
rect 10324 16405 10333 16439
rect 10333 16405 10367 16439
rect 10367 16405 10376 16439
rect 10692 16439 10744 16448
rect 10324 16396 10376 16405
rect 10692 16405 10701 16439
rect 10701 16405 10735 16439
rect 10735 16405 10744 16439
rect 10692 16396 10744 16405
rect 10968 16396 11020 16448
rect 12348 16396 12400 16448
rect 13820 16396 13872 16448
rect 15292 16464 15344 16516
rect 16304 16600 16356 16652
rect 18236 16677 18245 16711
rect 18245 16677 18279 16711
rect 18279 16677 18288 16711
rect 18236 16668 18288 16677
rect 17316 16643 17368 16652
rect 17316 16609 17325 16643
rect 17325 16609 17359 16643
rect 17359 16609 17368 16643
rect 17316 16600 17368 16609
rect 17500 16643 17552 16652
rect 17500 16609 17509 16643
rect 17509 16609 17543 16643
rect 17543 16609 17552 16643
rect 17500 16600 17552 16609
rect 20168 16600 20220 16652
rect 15200 16396 15252 16448
rect 16396 16464 16448 16516
rect 18144 16532 18196 16584
rect 15844 16396 15896 16448
rect 17592 16439 17644 16448
rect 17592 16405 17601 16439
rect 17601 16405 17635 16439
rect 17635 16405 17644 16439
rect 20076 16464 20128 16516
rect 17592 16396 17644 16405
rect 18512 16396 18564 16448
rect 19984 16396 20036 16448
rect 20996 16532 21048 16584
rect 20720 16464 20772 16516
rect 21088 16439 21140 16448
rect 21088 16405 21097 16439
rect 21097 16405 21131 16439
rect 21131 16405 21140 16439
rect 21088 16396 21140 16405
rect 21456 16439 21508 16448
rect 21456 16405 21465 16439
rect 21465 16405 21499 16439
rect 21499 16405 21508 16439
rect 21456 16396 21508 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 1676 16192 1728 16244
rect 2320 16235 2372 16244
rect 2320 16201 2329 16235
rect 2329 16201 2363 16235
rect 2363 16201 2372 16235
rect 2320 16192 2372 16201
rect 2412 16192 2464 16244
rect 3332 16235 3384 16244
rect 3332 16201 3341 16235
rect 3341 16201 3375 16235
rect 3375 16201 3384 16235
rect 3332 16192 3384 16201
rect 3884 16192 3936 16244
rect 5908 16192 5960 16244
rect 6828 16192 6880 16244
rect 8024 16192 8076 16244
rect 9128 16192 9180 16244
rect 9312 16235 9364 16244
rect 9312 16201 9321 16235
rect 9321 16201 9355 16235
rect 9355 16201 9364 16235
rect 9312 16192 9364 16201
rect 10232 16192 10284 16244
rect 10876 16192 10928 16244
rect 11796 16192 11848 16244
rect 13820 16192 13872 16244
rect 15108 16192 15160 16244
rect 15660 16192 15712 16244
rect 15844 16235 15896 16244
rect 15844 16201 15853 16235
rect 15853 16201 15887 16235
rect 15887 16201 15896 16235
rect 15844 16192 15896 16201
rect 16304 16192 16356 16244
rect 16948 16192 17000 16244
rect 17592 16192 17644 16244
rect 18788 16235 18840 16244
rect 18788 16201 18797 16235
rect 18797 16201 18831 16235
rect 18831 16201 18840 16235
rect 18788 16192 18840 16201
rect 20444 16235 20496 16244
rect 20444 16201 20453 16235
rect 20453 16201 20487 16235
rect 20487 16201 20496 16235
rect 20444 16192 20496 16201
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 20996 16235 21048 16244
rect 20996 16201 21005 16235
rect 21005 16201 21039 16235
rect 21039 16201 21048 16235
rect 20996 16192 21048 16201
rect 112 16124 164 16176
rect 1952 16056 2004 16108
rect 1860 15988 1912 16040
rect 2044 15920 2096 15972
rect 2688 16056 2740 16108
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 2780 15852 2832 15904
rect 3976 16124 4028 16176
rect 6000 16124 6052 16176
rect 7012 16124 7064 16176
rect 9036 16167 9088 16176
rect 4712 16056 4764 16108
rect 5356 16056 5408 16108
rect 3056 16031 3108 16040
rect 3056 15997 3065 16031
rect 3065 15997 3099 16031
rect 3099 15997 3108 16031
rect 3056 15988 3108 15997
rect 3240 16031 3292 16040
rect 3240 15997 3249 16031
rect 3249 15997 3283 16031
rect 3283 15997 3292 16031
rect 3240 15988 3292 15997
rect 4068 15988 4120 16040
rect 5080 16031 5132 16040
rect 5080 15997 5089 16031
rect 5089 15997 5123 16031
rect 5123 15997 5132 16031
rect 5080 15988 5132 15997
rect 5448 15988 5500 16040
rect 5632 16031 5684 16040
rect 5632 15997 5641 16031
rect 5641 15997 5675 16031
rect 5675 15997 5684 16031
rect 5632 15988 5684 15997
rect 9036 16133 9045 16167
rect 9045 16133 9079 16167
rect 9079 16133 9088 16167
rect 9036 16124 9088 16133
rect 11428 16124 11480 16176
rect 11888 16124 11940 16176
rect 14372 16124 14424 16176
rect 18512 16124 18564 16176
rect 3148 15920 3200 15972
rect 3884 15920 3936 15972
rect 7656 16031 7708 16040
rect 7656 15997 7665 16031
rect 7665 15997 7699 16031
rect 7699 15997 7708 16031
rect 9312 16056 9364 16108
rect 9680 16099 9732 16108
rect 9680 16065 9703 16099
rect 9703 16065 9732 16099
rect 9680 16056 9732 16065
rect 10508 16056 10560 16108
rect 13360 16099 13412 16108
rect 13360 16065 13369 16099
rect 13369 16065 13403 16099
rect 13403 16065 13412 16099
rect 13360 16056 13412 16065
rect 7656 15988 7708 15997
rect 8024 15963 8076 15972
rect 8024 15929 8033 15963
rect 8033 15929 8067 15963
rect 8067 15929 8076 15963
rect 8024 15920 8076 15929
rect 3056 15852 3108 15904
rect 6828 15852 6880 15904
rect 7748 15852 7800 15904
rect 8208 15852 8260 15904
rect 13728 15988 13780 16040
rect 14280 16056 14332 16108
rect 15108 16056 15160 16108
rect 18604 16056 18656 16108
rect 20260 16099 20312 16108
rect 20260 16065 20269 16099
rect 20269 16065 20303 16099
rect 20303 16065 20312 16099
rect 20260 16056 20312 16065
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 21272 16099 21324 16108
rect 15292 16031 15344 16040
rect 15292 15997 15301 16031
rect 15301 15997 15335 16031
rect 15335 15997 15344 16031
rect 15292 15988 15344 15997
rect 16304 15988 16356 16040
rect 17132 16031 17184 16040
rect 17132 15997 17141 16031
rect 17141 15997 17175 16031
rect 17175 15997 17184 16031
rect 17132 15988 17184 15997
rect 9680 15852 9732 15904
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 11980 15895 12032 15904
rect 11980 15861 11989 15895
rect 11989 15861 12023 15895
rect 12023 15861 12032 15895
rect 11980 15852 12032 15861
rect 12072 15852 12124 15904
rect 14556 15920 14608 15972
rect 17776 15988 17828 16040
rect 19064 15988 19116 16040
rect 21272 16065 21281 16099
rect 21281 16065 21315 16099
rect 21315 16065 21324 16099
rect 21272 16056 21324 16065
rect 13820 15852 13872 15904
rect 15292 15852 15344 15904
rect 21456 15895 21508 15904
rect 21456 15861 21465 15895
rect 21465 15861 21499 15895
rect 21499 15861 21508 15895
rect 21456 15852 21508 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1768 15648 1820 15700
rect 1952 15648 2004 15700
rect 2228 15648 2280 15700
rect 2964 15648 3016 15700
rect 3240 15648 3292 15700
rect 4160 15648 4212 15700
rect 4988 15691 5040 15700
rect 4988 15657 4997 15691
rect 4997 15657 5031 15691
rect 5031 15657 5040 15691
rect 4988 15648 5040 15657
rect 5356 15648 5408 15700
rect 5724 15648 5776 15700
rect 6920 15648 6972 15700
rect 7748 15648 7800 15700
rect 8668 15648 8720 15700
rect 10784 15648 10836 15700
rect 12072 15648 12124 15700
rect 12256 15648 12308 15700
rect 13176 15648 13228 15700
rect 13820 15648 13872 15700
rect 14372 15648 14424 15700
rect 2780 15580 2832 15632
rect 204 15512 256 15564
rect 296 15376 348 15428
rect 2228 15444 2280 15496
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2596 15487 2648 15496
rect 2320 15444 2372 15453
rect 2596 15453 2605 15487
rect 2605 15453 2639 15487
rect 2639 15453 2648 15487
rect 2596 15444 2648 15453
rect 2872 15512 2924 15564
rect 4068 15512 4120 15564
rect 4620 15512 4672 15564
rect 5080 15512 5132 15564
rect 6000 15555 6052 15564
rect 6000 15521 6009 15555
rect 6009 15521 6043 15555
rect 6043 15521 6052 15555
rect 6000 15512 6052 15521
rect 7104 15555 7156 15564
rect 7104 15521 7113 15555
rect 7113 15521 7147 15555
rect 7147 15521 7156 15555
rect 7104 15512 7156 15521
rect 10508 15555 10560 15564
rect 10508 15521 10517 15555
rect 10517 15521 10551 15555
rect 10551 15521 10560 15555
rect 10508 15512 10560 15521
rect 12716 15580 12768 15632
rect 12808 15580 12860 15632
rect 13728 15580 13780 15632
rect 17316 15648 17368 15700
rect 12624 15555 12676 15564
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 13176 15512 13228 15564
rect 14372 15512 14424 15564
rect 18604 15648 18656 15700
rect 19432 15648 19484 15700
rect 20536 15648 20588 15700
rect 21272 15648 21324 15700
rect 18512 15580 18564 15632
rect 2780 15444 2832 15496
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 3056 15444 3108 15496
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 2412 15376 2464 15428
rect 4988 15444 5040 15496
rect 5356 15419 5408 15428
rect 5356 15385 5365 15419
rect 5365 15385 5399 15419
rect 5399 15385 5408 15419
rect 5356 15376 5408 15385
rect 7932 15444 7984 15496
rect 8208 15444 8260 15496
rect 9680 15444 9732 15496
rect 10232 15444 10284 15496
rect 11704 15444 11756 15496
rect 11980 15444 12032 15496
rect 12532 15444 12584 15496
rect 14280 15444 14332 15496
rect 15108 15444 15160 15496
rect 3056 15308 3108 15360
rect 3332 15308 3384 15360
rect 4160 15351 4212 15360
rect 4160 15317 4169 15351
rect 4169 15317 4203 15351
rect 4203 15317 4212 15351
rect 4160 15308 4212 15317
rect 4896 15308 4948 15360
rect 6000 15308 6052 15360
rect 6552 15351 6604 15360
rect 6552 15317 6561 15351
rect 6561 15317 6595 15351
rect 6595 15317 6604 15351
rect 6552 15308 6604 15317
rect 6920 15351 6972 15360
rect 6920 15317 6929 15351
rect 6929 15317 6963 15351
rect 6963 15317 6972 15351
rect 6920 15308 6972 15317
rect 7012 15351 7064 15360
rect 7012 15317 7021 15351
rect 7021 15317 7055 15351
rect 7055 15317 7064 15351
rect 8668 15376 8720 15428
rect 9220 15419 9272 15428
rect 7012 15308 7064 15317
rect 8116 15308 8168 15360
rect 9220 15385 9254 15419
rect 9254 15385 9272 15419
rect 9220 15376 9272 15385
rect 10876 15376 10928 15428
rect 11428 15376 11480 15428
rect 12072 15376 12124 15428
rect 13452 15376 13504 15428
rect 9404 15308 9456 15360
rect 12992 15308 13044 15360
rect 13636 15351 13688 15360
rect 13636 15317 13645 15351
rect 13645 15317 13679 15351
rect 13679 15317 13688 15351
rect 13636 15308 13688 15317
rect 14188 15308 14240 15360
rect 14556 15351 14608 15360
rect 14556 15317 14565 15351
rect 14565 15317 14599 15351
rect 14599 15317 14608 15351
rect 14556 15308 14608 15317
rect 15016 15308 15068 15360
rect 16948 15444 17000 15496
rect 19248 15512 19300 15564
rect 19432 15444 19484 15496
rect 19524 15444 19576 15496
rect 20076 15487 20128 15496
rect 20076 15453 20085 15487
rect 20085 15453 20119 15487
rect 20119 15453 20128 15487
rect 20076 15444 20128 15453
rect 15752 15376 15804 15428
rect 17776 15376 17828 15428
rect 17132 15308 17184 15360
rect 18788 15351 18840 15360
rect 18788 15317 18797 15351
rect 18797 15317 18831 15351
rect 18831 15317 18840 15351
rect 18788 15308 18840 15317
rect 21180 15351 21232 15360
rect 21180 15317 21189 15351
rect 21189 15317 21223 15351
rect 21223 15317 21232 15351
rect 21180 15308 21232 15317
rect 21456 15351 21508 15360
rect 21456 15317 21465 15351
rect 21465 15317 21499 15351
rect 21499 15317 21508 15351
rect 21456 15308 21508 15317
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 1676 15011 1728 15020
rect 1676 14977 1685 15011
rect 1685 14977 1719 15011
rect 1719 14977 1728 15011
rect 1676 14968 1728 14977
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 2412 15147 2464 15156
rect 2412 15113 2421 15147
rect 2421 15113 2455 15147
rect 2455 15113 2464 15147
rect 2412 15104 2464 15113
rect 6552 15104 6604 15156
rect 7012 15104 7064 15156
rect 7380 15147 7432 15156
rect 7380 15113 7389 15147
rect 7389 15113 7423 15147
rect 7423 15113 7432 15147
rect 7380 15104 7432 15113
rect 7748 15104 7800 15156
rect 8300 15104 8352 15156
rect 8484 15147 8536 15156
rect 8484 15113 8493 15147
rect 8493 15113 8527 15147
rect 8527 15113 8536 15147
rect 8484 15104 8536 15113
rect 8576 15147 8628 15156
rect 8576 15113 8585 15147
rect 8585 15113 8619 15147
rect 8619 15113 8628 15147
rect 8576 15104 8628 15113
rect 9588 15104 9640 15156
rect 9864 15104 9916 15156
rect 4068 15036 4120 15088
rect 5540 15036 5592 15088
rect 4252 14968 4304 15020
rect 4528 14968 4580 15020
rect 4804 14968 4856 15020
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 5908 14968 5960 15020
rect 9128 15036 9180 15088
rect 8208 14968 8260 15020
rect 5264 14943 5316 14952
rect 5264 14909 5273 14943
rect 5273 14909 5307 14943
rect 5307 14909 5316 14943
rect 5264 14900 5316 14909
rect 5632 14900 5684 14952
rect 7196 14900 7248 14952
rect 7564 14943 7616 14952
rect 7564 14909 7573 14943
rect 7573 14909 7607 14943
rect 7607 14909 7616 14943
rect 7564 14900 7616 14909
rect 9220 14943 9272 14952
rect 9220 14909 9229 14943
rect 9229 14909 9263 14943
rect 9263 14909 9272 14943
rect 9220 14900 9272 14909
rect 1860 14875 1912 14884
rect 1860 14841 1869 14875
rect 1869 14841 1903 14875
rect 1903 14841 1912 14875
rect 1860 14832 1912 14841
rect 2872 14832 2924 14884
rect 4528 14875 4580 14884
rect 4528 14841 4537 14875
rect 4537 14841 4571 14875
rect 4571 14841 4580 14875
rect 4528 14832 4580 14841
rect 6460 14875 6512 14884
rect 6460 14841 6469 14875
rect 6469 14841 6503 14875
rect 6503 14841 6512 14875
rect 6460 14832 6512 14841
rect 6552 14832 6604 14884
rect 6828 14832 6880 14884
rect 7012 14832 7064 14884
rect 9128 14832 9180 14884
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 4344 14764 4396 14816
rect 5356 14764 5408 14816
rect 6000 14764 6052 14816
rect 7840 14807 7892 14816
rect 7840 14773 7849 14807
rect 7849 14773 7883 14807
rect 7883 14773 7892 14807
rect 7840 14764 7892 14773
rect 9680 14900 9732 14952
rect 10416 15036 10468 15088
rect 12256 15036 12308 15088
rect 13820 15104 13872 15156
rect 14464 15147 14516 15156
rect 14464 15113 14473 15147
rect 14473 15113 14507 15147
rect 14507 15113 14516 15147
rect 14464 15104 14516 15113
rect 16948 15147 17000 15156
rect 16948 15113 16957 15147
rect 16957 15113 16991 15147
rect 16991 15113 17000 15147
rect 16948 15104 17000 15113
rect 11704 14968 11756 15020
rect 10324 14943 10376 14952
rect 10324 14909 10333 14943
rect 10333 14909 10367 14943
rect 10367 14909 10376 14943
rect 10324 14900 10376 14909
rect 10416 14943 10468 14952
rect 10416 14909 10425 14943
rect 10425 14909 10459 14943
rect 10459 14909 10468 14943
rect 10416 14900 10468 14909
rect 10784 14900 10836 14952
rect 9404 14764 9456 14816
rect 9496 14764 9548 14816
rect 10968 14807 11020 14816
rect 10968 14773 10977 14807
rect 10977 14773 11011 14807
rect 11011 14773 11020 14807
rect 10968 14764 11020 14773
rect 12716 14943 12768 14952
rect 12716 14909 12725 14943
rect 12725 14909 12759 14943
rect 12759 14909 12768 14943
rect 12716 14900 12768 14909
rect 13636 15036 13688 15088
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 14832 15036 14884 15088
rect 17316 15036 17368 15088
rect 19524 15104 19576 15156
rect 20260 15104 20312 15156
rect 19984 15036 20036 15088
rect 22652 15104 22704 15156
rect 22192 15036 22244 15088
rect 14372 14968 14424 15020
rect 15016 15011 15068 15020
rect 15016 14977 15025 15011
rect 15025 14977 15059 15011
rect 15059 14977 15068 15011
rect 15016 14968 15068 14977
rect 16028 15011 16080 15020
rect 16028 14977 16037 15011
rect 16037 14977 16071 15011
rect 16071 14977 16080 15011
rect 16028 14968 16080 14977
rect 18052 14968 18104 15020
rect 19708 15011 19760 15020
rect 19708 14977 19717 15011
rect 19717 14977 19751 15011
rect 19751 14977 19760 15011
rect 19708 14968 19760 14977
rect 20720 14968 20772 15020
rect 20996 14968 21048 15020
rect 13728 14900 13780 14952
rect 14004 14943 14056 14952
rect 14004 14909 14013 14943
rect 14013 14909 14047 14943
rect 14047 14909 14056 14943
rect 14004 14900 14056 14909
rect 15752 14943 15804 14952
rect 15752 14909 15761 14943
rect 15761 14909 15795 14943
rect 15795 14909 15804 14943
rect 15752 14900 15804 14909
rect 15936 14943 15988 14952
rect 15936 14909 15945 14943
rect 15945 14909 15979 14943
rect 15979 14909 15988 14943
rect 15936 14900 15988 14909
rect 18604 14900 18656 14952
rect 21364 14900 21416 14952
rect 21088 14875 21140 14884
rect 21088 14841 21097 14875
rect 21097 14841 21131 14875
rect 21131 14841 21140 14875
rect 21088 14832 21140 14841
rect 12624 14764 12676 14816
rect 12900 14764 12952 14816
rect 13360 14807 13412 14816
rect 13360 14773 13369 14807
rect 13369 14773 13403 14807
rect 13403 14773 13412 14807
rect 13360 14764 13412 14773
rect 15200 14807 15252 14816
rect 15200 14773 15209 14807
rect 15209 14773 15243 14807
rect 15243 14773 15252 14807
rect 15200 14764 15252 14773
rect 16856 14764 16908 14816
rect 17960 14764 18012 14816
rect 22284 14832 22336 14884
rect 21456 14807 21508 14816
rect 21456 14773 21465 14807
rect 21465 14773 21499 14807
rect 21499 14773 21508 14807
rect 21456 14764 21508 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 1676 14560 1728 14612
rect 2228 14560 2280 14612
rect 2964 14560 3016 14612
rect 4804 14603 4856 14612
rect 4804 14569 4813 14603
rect 4813 14569 4847 14603
rect 4847 14569 4856 14603
rect 4804 14560 4856 14569
rect 5264 14560 5316 14612
rect 6828 14560 6880 14612
rect 6920 14560 6972 14612
rect 8576 14560 8628 14612
rect 10508 14560 10560 14612
rect 2044 14492 2096 14544
rect 2780 14492 2832 14544
rect 10692 14492 10744 14544
rect 3240 14467 3292 14476
rect 2044 14399 2096 14408
rect 2044 14365 2053 14399
rect 2053 14365 2087 14399
rect 2087 14365 2096 14399
rect 2044 14356 2096 14365
rect 3240 14433 3249 14467
rect 3249 14433 3283 14467
rect 3283 14433 3292 14467
rect 3240 14424 3292 14433
rect 8484 14467 8536 14476
rect 2412 14356 2464 14408
rect 3884 14288 3936 14340
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 4344 14263 4396 14272
rect 4344 14229 4353 14263
rect 4353 14229 4387 14263
rect 4387 14229 4396 14263
rect 4344 14220 4396 14229
rect 4436 14263 4488 14272
rect 4436 14229 4445 14263
rect 4445 14229 4479 14263
rect 4479 14229 4488 14263
rect 5632 14356 5684 14408
rect 6460 14356 6512 14408
rect 7288 14356 7340 14408
rect 7564 14399 7616 14408
rect 7564 14365 7593 14399
rect 7593 14365 7616 14399
rect 8484 14433 8493 14467
rect 8493 14433 8527 14467
rect 8527 14433 8536 14467
rect 8484 14424 8536 14433
rect 8944 14424 8996 14476
rect 7564 14356 7616 14365
rect 7932 14356 7984 14408
rect 8300 14356 8352 14408
rect 10324 14424 10376 14476
rect 10784 14424 10836 14476
rect 13820 14424 13872 14476
rect 15752 14560 15804 14612
rect 16856 14492 16908 14544
rect 17500 14560 17552 14612
rect 19524 14560 19576 14612
rect 20720 14603 20772 14612
rect 20720 14569 20729 14603
rect 20729 14569 20763 14603
rect 20763 14569 20772 14603
rect 20720 14560 20772 14569
rect 20996 14603 21048 14612
rect 20996 14569 21005 14603
rect 21005 14569 21039 14603
rect 21039 14569 21048 14603
rect 20996 14560 21048 14569
rect 17132 14467 17184 14476
rect 9496 14399 9548 14408
rect 9496 14365 9505 14399
rect 9505 14365 9539 14399
rect 9539 14365 9548 14399
rect 9496 14356 9548 14365
rect 10692 14356 10744 14408
rect 11888 14399 11940 14408
rect 11888 14365 11906 14399
rect 11906 14365 11940 14399
rect 11888 14356 11940 14365
rect 4988 14288 5040 14340
rect 10876 14288 10928 14340
rect 11704 14288 11756 14340
rect 13636 14356 13688 14408
rect 14188 14356 14240 14408
rect 17132 14433 17141 14467
rect 17141 14433 17175 14467
rect 17175 14433 17184 14467
rect 17132 14424 17184 14433
rect 19064 14492 19116 14544
rect 17776 14424 17828 14476
rect 20996 14356 21048 14408
rect 4436 14220 4488 14229
rect 5448 14220 5500 14272
rect 7104 14220 7156 14272
rect 7840 14220 7892 14272
rect 9312 14220 9364 14272
rect 9864 14220 9916 14272
rect 10324 14263 10376 14272
rect 10324 14229 10333 14263
rect 10333 14229 10367 14263
rect 10367 14229 10376 14263
rect 10324 14220 10376 14229
rect 12716 14288 12768 14340
rect 12808 14220 12860 14272
rect 14832 14288 14884 14340
rect 15108 14288 15160 14340
rect 15844 14331 15896 14340
rect 15568 14220 15620 14272
rect 15844 14297 15878 14331
rect 15878 14297 15896 14331
rect 15844 14288 15896 14297
rect 17132 14288 17184 14340
rect 17408 14263 17460 14272
rect 17408 14229 17417 14263
rect 17417 14229 17451 14263
rect 17451 14229 17460 14263
rect 18512 14288 18564 14340
rect 20076 14288 20128 14340
rect 22928 14288 22980 14340
rect 17408 14220 17460 14229
rect 18328 14220 18380 14272
rect 18880 14263 18932 14272
rect 18880 14229 18889 14263
rect 18889 14229 18923 14263
rect 18923 14229 18932 14263
rect 18880 14220 18932 14229
rect 19616 14263 19668 14272
rect 19616 14229 19625 14263
rect 19625 14229 19659 14263
rect 19659 14229 19668 14263
rect 19616 14220 19668 14229
rect 19984 14263 20036 14272
rect 19984 14229 19993 14263
rect 19993 14229 20027 14263
rect 20027 14229 20036 14263
rect 19984 14220 20036 14229
rect 21456 14263 21508 14272
rect 21456 14229 21465 14263
rect 21465 14229 21499 14263
rect 21499 14229 21508 14263
rect 21456 14220 21508 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 2412 14016 2464 14068
rect 3424 14016 3476 14068
rect 3240 13948 3292 14000
rect 4804 13948 4856 14000
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 3884 13880 3936 13932
rect 4068 13880 4120 13932
rect 4252 13923 4304 13932
rect 4252 13889 4261 13923
rect 4261 13889 4295 13923
rect 4295 13889 4304 13923
rect 4252 13880 4304 13889
rect 4988 14016 5040 14068
rect 5632 14059 5684 14068
rect 5632 14025 5641 14059
rect 5641 14025 5675 14059
rect 5675 14025 5684 14059
rect 5632 14016 5684 14025
rect 5908 13948 5960 14000
rect 7840 14016 7892 14068
rect 9404 14059 9456 14068
rect 6828 13948 6880 14000
rect 9404 14025 9413 14059
rect 9413 14025 9447 14059
rect 9447 14025 9456 14059
rect 9404 14016 9456 14025
rect 9496 14016 9548 14068
rect 9864 14059 9916 14068
rect 7932 13880 7984 13932
rect 8116 13880 8168 13932
rect 9036 13880 9088 13932
rect 2504 13744 2556 13796
rect 3332 13812 3384 13864
rect 4160 13855 4212 13864
rect 4160 13821 4169 13855
rect 4169 13821 4203 13855
rect 4203 13821 4212 13855
rect 4160 13812 4212 13821
rect 5264 13812 5316 13864
rect 4252 13744 4304 13796
rect 5356 13744 5408 13796
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 8392 13812 8444 13864
rect 9864 14025 9873 14059
rect 9873 14025 9907 14059
rect 9907 14025 9916 14059
rect 9864 14016 9916 14025
rect 10508 14016 10560 14068
rect 11060 14059 11112 14068
rect 11060 14025 11069 14059
rect 11069 14025 11103 14059
rect 11103 14025 11112 14059
rect 11060 14016 11112 14025
rect 11796 14016 11848 14068
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 12256 14016 12308 14068
rect 12716 14016 12768 14068
rect 12900 14016 12952 14068
rect 13452 14059 13504 14068
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 13728 14016 13780 14068
rect 9772 13948 9824 14000
rect 11520 13991 11572 14000
rect 10232 13923 10284 13932
rect 10232 13889 10241 13923
rect 10241 13889 10275 13923
rect 10275 13889 10284 13923
rect 10232 13880 10284 13889
rect 11520 13957 11529 13991
rect 11529 13957 11563 13991
rect 11563 13957 11572 13991
rect 11520 13948 11572 13957
rect 11980 13880 12032 13932
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 2320 13676 2372 13728
rect 3976 13676 4028 13728
rect 4528 13676 4580 13728
rect 4988 13676 5040 13728
rect 5816 13676 5868 13728
rect 6092 13744 6144 13796
rect 6184 13744 6236 13796
rect 6644 13744 6696 13796
rect 8944 13787 8996 13796
rect 8944 13753 8953 13787
rect 8953 13753 8987 13787
rect 8987 13753 8996 13787
rect 8944 13744 8996 13753
rect 10416 13855 10468 13864
rect 10416 13821 10425 13855
rect 10425 13821 10459 13855
rect 10459 13821 10468 13855
rect 10876 13855 10928 13864
rect 10416 13812 10468 13821
rect 10876 13821 10885 13855
rect 10885 13821 10919 13855
rect 10919 13821 10928 13855
rect 10876 13812 10928 13821
rect 11336 13812 11388 13864
rect 11796 13812 11848 13864
rect 12256 13855 12308 13864
rect 12256 13821 12265 13855
rect 12265 13821 12299 13855
rect 12299 13821 12308 13855
rect 12256 13812 12308 13821
rect 13452 13880 13504 13932
rect 13820 13923 13872 13932
rect 13820 13889 13829 13923
rect 13829 13889 13863 13923
rect 13863 13889 13872 13923
rect 13820 13880 13872 13889
rect 14280 13880 14332 13932
rect 14372 13923 14424 13932
rect 14372 13889 14381 13923
rect 14381 13889 14415 13923
rect 14415 13889 14424 13923
rect 15936 14016 15988 14068
rect 17408 14016 17460 14068
rect 20996 14059 21048 14068
rect 20996 14025 21005 14059
rect 21005 14025 21039 14059
rect 21039 14025 21048 14059
rect 20996 14016 21048 14025
rect 15752 13948 15804 14000
rect 14372 13880 14424 13889
rect 11612 13744 11664 13796
rect 14004 13812 14056 13864
rect 14188 13812 14240 13864
rect 15016 13812 15068 13864
rect 15752 13812 15804 13864
rect 15936 13880 15988 13932
rect 17592 13880 17644 13932
rect 18788 13948 18840 14000
rect 17960 13923 18012 13932
rect 17960 13889 17994 13923
rect 17994 13889 18012 13923
rect 17960 13880 18012 13889
rect 19064 13880 19116 13932
rect 19524 13923 19576 13932
rect 19524 13889 19533 13923
rect 19533 13889 19567 13923
rect 19567 13889 19576 13923
rect 19524 13880 19576 13889
rect 16396 13812 16448 13864
rect 20168 13855 20220 13864
rect 16212 13744 16264 13796
rect 17408 13744 17460 13796
rect 18972 13744 19024 13796
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 20352 13855 20404 13864
rect 20352 13821 20361 13855
rect 20361 13821 20395 13855
rect 20395 13821 20404 13855
rect 20720 13880 20772 13932
rect 20996 13880 21048 13932
rect 20352 13812 20404 13821
rect 21272 13744 21324 13796
rect 7840 13676 7892 13728
rect 8668 13676 8720 13728
rect 9128 13676 9180 13728
rect 9312 13676 9364 13728
rect 9956 13676 10008 13728
rect 13820 13676 13872 13728
rect 14372 13676 14424 13728
rect 15752 13676 15804 13728
rect 17500 13676 17552 13728
rect 18880 13676 18932 13728
rect 19892 13719 19944 13728
rect 19892 13685 19901 13719
rect 19901 13685 19935 13719
rect 19935 13685 19944 13719
rect 19892 13676 19944 13685
rect 21456 13719 21508 13728
rect 21456 13685 21465 13719
rect 21465 13685 21499 13719
rect 21499 13685 21508 13719
rect 21456 13676 21508 13685
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 4436 13472 4488 13524
rect 4528 13472 4580 13524
rect 4344 13404 4396 13456
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 2044 13311 2096 13320
rect 2044 13277 2053 13311
rect 2053 13277 2087 13311
rect 2087 13277 2096 13311
rect 2044 13268 2096 13277
rect 4528 13336 4580 13388
rect 4804 13379 4856 13388
rect 4804 13345 4813 13379
rect 4813 13345 4847 13379
rect 4847 13345 4856 13379
rect 4804 13336 4856 13345
rect 5448 13336 5500 13388
rect 6092 13472 6144 13524
rect 8576 13472 8628 13524
rect 12072 13472 12124 13524
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 13084 13472 13136 13524
rect 13544 13472 13596 13524
rect 13820 13472 13872 13524
rect 15936 13472 15988 13524
rect 16028 13472 16080 13524
rect 18972 13515 19024 13524
rect 18972 13481 18981 13515
rect 18981 13481 19015 13515
rect 19015 13481 19024 13515
rect 18972 13472 19024 13481
rect 19064 13472 19116 13524
rect 19708 13472 19760 13524
rect 7012 13404 7064 13456
rect 3976 13268 4028 13320
rect 4068 13268 4120 13320
rect 5632 13268 5684 13320
rect 848 13200 900 13252
rect 4344 13200 4396 13252
rect 4436 13200 4488 13252
rect 5540 13200 5592 13252
rect 6000 13243 6052 13252
rect 6000 13209 6009 13243
rect 6009 13209 6043 13243
rect 6043 13209 6052 13243
rect 6000 13200 6052 13209
rect 6552 13268 6604 13320
rect 7104 13336 7156 13388
rect 9220 13404 9272 13456
rect 10600 13404 10652 13456
rect 9496 13268 9548 13320
rect 9772 13268 9824 13320
rect 6644 13200 6696 13252
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 1860 13175 1912 13184
rect 1860 13141 1869 13175
rect 1869 13141 1903 13175
rect 1903 13141 1912 13175
rect 1860 13132 1912 13141
rect 2228 13175 2280 13184
rect 2228 13141 2237 13175
rect 2237 13141 2271 13175
rect 2271 13141 2280 13175
rect 2228 13132 2280 13141
rect 2780 13132 2832 13184
rect 3884 13132 3936 13184
rect 5264 13132 5316 13184
rect 5448 13175 5500 13184
rect 5448 13141 5457 13175
rect 5457 13141 5491 13175
rect 5491 13141 5500 13175
rect 6184 13175 6236 13184
rect 5448 13132 5500 13141
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 6184 13132 6236 13141
rect 6552 13175 6604 13184
rect 6552 13141 6561 13175
rect 6561 13141 6595 13175
rect 6595 13141 6604 13175
rect 6552 13132 6604 13141
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 8116 13132 8168 13184
rect 9312 13132 9364 13184
rect 9588 13200 9640 13252
rect 10048 13243 10100 13252
rect 10048 13209 10066 13243
rect 10066 13209 10100 13243
rect 12256 13404 12308 13456
rect 12532 13447 12584 13456
rect 12532 13413 12541 13447
rect 12541 13413 12575 13447
rect 12575 13413 12584 13447
rect 12532 13404 12584 13413
rect 14372 13404 14424 13456
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 11796 13268 11848 13320
rect 12164 13336 12216 13388
rect 12808 13379 12860 13388
rect 12808 13345 12817 13379
rect 12817 13345 12851 13379
rect 12851 13345 12860 13379
rect 12808 13336 12860 13345
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 12992 13336 13044 13345
rect 15844 13336 15896 13388
rect 16948 13336 17000 13388
rect 17592 13379 17644 13388
rect 10048 13200 10100 13209
rect 10692 13200 10744 13252
rect 10600 13132 10652 13184
rect 11152 13132 11204 13184
rect 11336 13132 11388 13184
rect 11612 13200 11664 13252
rect 13360 13268 13412 13320
rect 13636 13311 13688 13320
rect 13636 13277 13645 13311
rect 13645 13277 13679 13311
rect 13679 13277 13688 13311
rect 13636 13268 13688 13277
rect 13820 13268 13872 13320
rect 15108 13268 15160 13320
rect 15384 13268 15436 13320
rect 17592 13345 17601 13379
rect 17601 13345 17635 13379
rect 17635 13345 17644 13379
rect 17592 13336 17644 13345
rect 18880 13336 18932 13388
rect 20536 13336 20588 13388
rect 17500 13268 17552 13320
rect 19708 13268 19760 13320
rect 19892 13268 19944 13320
rect 21272 13311 21324 13320
rect 21272 13277 21281 13311
rect 21281 13277 21315 13311
rect 21315 13277 21324 13311
rect 21272 13268 21324 13277
rect 12164 13132 12216 13184
rect 14464 13200 14516 13252
rect 15200 13200 15252 13252
rect 17684 13200 17736 13252
rect 18236 13200 18288 13252
rect 20628 13200 20680 13252
rect 16304 13132 16356 13184
rect 17224 13175 17276 13184
rect 17224 13141 17233 13175
rect 17233 13141 17267 13175
rect 17267 13141 17276 13175
rect 17224 13132 17276 13141
rect 18328 13132 18380 13184
rect 18788 13132 18840 13184
rect 21088 13175 21140 13184
rect 21088 13141 21097 13175
rect 21097 13141 21131 13175
rect 21131 13141 21140 13175
rect 21088 13132 21140 13141
rect 21456 13175 21508 13184
rect 21456 13141 21465 13175
rect 21465 13141 21499 13175
rect 21499 13141 21508 13175
rect 21456 13132 21508 13141
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 1676 12928 1728 12980
rect 3240 12971 3292 12980
rect 3240 12937 3249 12971
rect 3249 12937 3283 12971
rect 3283 12937 3292 12971
rect 3240 12928 3292 12937
rect 3332 12928 3384 12980
rect 6368 12928 6420 12980
rect 7380 12928 7432 12980
rect 8300 12971 8352 12980
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 8668 12928 8720 12980
rect 9128 12971 9180 12980
rect 9128 12937 9137 12971
rect 9137 12937 9171 12971
rect 9171 12937 9180 12971
rect 9128 12928 9180 12937
rect 9496 12971 9548 12980
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 9680 12928 9732 12980
rect 9864 12971 9916 12980
rect 9864 12937 9873 12971
rect 9873 12937 9907 12971
rect 9907 12937 9916 12971
rect 9864 12928 9916 12937
rect 10968 12928 11020 12980
rect 11428 12928 11480 12980
rect 2228 12860 2280 12912
rect 3332 12792 3384 12844
rect 2872 12767 2924 12776
rect 2872 12733 2881 12767
rect 2881 12733 2915 12767
rect 2915 12733 2924 12767
rect 2872 12724 2924 12733
rect 4252 12860 4304 12912
rect 5632 12860 5684 12912
rect 6184 12860 6236 12912
rect 4620 12792 4672 12844
rect 5356 12792 5408 12844
rect 5540 12792 5592 12844
rect 5724 12792 5776 12844
rect 5908 12792 5960 12844
rect 6644 12835 6696 12844
rect 6644 12801 6678 12835
rect 6678 12801 6696 12835
rect 6644 12792 6696 12801
rect 7196 12860 7248 12912
rect 7656 12860 7708 12912
rect 8024 12860 8076 12912
rect 4344 12767 4396 12776
rect 4344 12733 4353 12767
rect 4353 12733 4387 12767
rect 4387 12733 4396 12767
rect 4344 12724 4396 12733
rect 5632 12724 5684 12776
rect 6000 12724 6052 12776
rect 8576 12860 8628 12912
rect 11060 12860 11112 12912
rect 12164 12928 12216 12980
rect 13360 12971 13412 12980
rect 13360 12937 13369 12971
rect 13369 12937 13403 12971
rect 13403 12937 13412 12971
rect 13360 12928 13412 12937
rect 15200 12971 15252 12980
rect 15200 12937 15209 12971
rect 15209 12937 15243 12971
rect 15243 12937 15252 12971
rect 15200 12928 15252 12937
rect 18236 12971 18288 12980
rect 18236 12937 18245 12971
rect 18245 12937 18279 12971
rect 18279 12937 18288 12971
rect 18236 12928 18288 12937
rect 19524 12928 19576 12980
rect 20168 12971 20220 12980
rect 20168 12937 20177 12971
rect 20177 12937 20211 12971
rect 20211 12937 20220 12971
rect 20168 12928 20220 12937
rect 20444 12928 20496 12980
rect 20812 12928 20864 12980
rect 20996 12971 21048 12980
rect 20996 12937 21005 12971
rect 21005 12937 21039 12971
rect 21039 12937 21048 12971
rect 20996 12928 21048 12937
rect 9864 12792 9916 12844
rect 12992 12860 13044 12912
rect 14280 12860 14332 12912
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 13176 12792 13228 12844
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 8484 12767 8536 12776
rect 8484 12733 8493 12767
rect 8493 12733 8527 12767
rect 8527 12733 8536 12767
rect 9220 12767 9272 12776
rect 8484 12724 8536 12733
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 10324 12767 10376 12776
rect 10324 12733 10333 12767
rect 10333 12733 10367 12767
rect 10367 12733 10376 12767
rect 10324 12724 10376 12733
rect 10784 12724 10836 12776
rect 12532 12724 12584 12776
rect 12808 12724 12860 12776
rect 15476 12860 15528 12912
rect 15660 12835 15712 12844
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 16212 12792 16264 12844
rect 18972 12860 19024 12912
rect 18236 12792 18288 12844
rect 18328 12835 18380 12844
rect 18328 12801 18337 12835
rect 18337 12801 18371 12835
rect 18371 12801 18380 12835
rect 18328 12792 18380 12801
rect 18880 12792 18932 12844
rect 20812 12835 20864 12844
rect 4252 12656 4304 12708
rect 4712 12656 4764 12708
rect 4896 12656 4948 12708
rect 8576 12656 8628 12708
rect 2504 12588 2556 12640
rect 3792 12588 3844 12640
rect 3976 12588 4028 12640
rect 4988 12588 5040 12640
rect 5356 12588 5408 12640
rect 6276 12588 6328 12640
rect 6368 12588 6420 12640
rect 9128 12588 9180 12640
rect 10876 12588 10928 12640
rect 11060 12588 11112 12640
rect 13084 12588 13136 12640
rect 15108 12656 15160 12708
rect 16580 12656 16632 12708
rect 16764 12631 16816 12640
rect 16764 12597 16773 12631
rect 16773 12597 16807 12631
rect 16807 12597 16816 12631
rect 16764 12588 16816 12597
rect 17040 12631 17092 12640
rect 17040 12597 17049 12631
rect 17049 12597 17083 12631
rect 17083 12597 17092 12631
rect 17040 12588 17092 12597
rect 17408 12631 17460 12640
rect 17408 12597 17417 12631
rect 17417 12597 17451 12631
rect 17451 12597 17460 12631
rect 17408 12588 17460 12597
rect 18052 12724 18104 12776
rect 20812 12801 20821 12835
rect 20821 12801 20855 12835
rect 20855 12801 20864 12835
rect 20812 12792 20864 12801
rect 20996 12792 21048 12844
rect 21272 12835 21324 12844
rect 21272 12801 21281 12835
rect 21281 12801 21315 12835
rect 21315 12801 21324 12835
rect 21272 12792 21324 12801
rect 19524 12656 19576 12708
rect 20536 12656 20588 12708
rect 21548 12656 21600 12708
rect 20444 12588 20496 12640
rect 21456 12631 21508 12640
rect 21456 12597 21465 12631
rect 21465 12597 21499 12631
rect 21499 12597 21508 12631
rect 21456 12588 21508 12597
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 1492 12427 1544 12436
rect 1492 12393 1501 12427
rect 1501 12393 1535 12427
rect 1535 12393 1544 12427
rect 1492 12384 1544 12393
rect 3976 12427 4028 12436
rect 3976 12393 3985 12427
rect 3985 12393 4019 12427
rect 4019 12393 4028 12427
rect 3976 12384 4028 12393
rect 4252 12384 4304 12436
rect 6368 12384 6420 12436
rect 7380 12384 7432 12436
rect 7932 12384 7984 12436
rect 8300 12384 8352 12436
rect 8760 12384 8812 12436
rect 9496 12427 9548 12436
rect 9496 12393 9505 12427
rect 9505 12393 9539 12427
rect 9539 12393 9548 12427
rect 9496 12384 9548 12393
rect 10600 12427 10652 12436
rect 10600 12393 10609 12427
rect 10609 12393 10643 12427
rect 10643 12393 10652 12427
rect 10600 12384 10652 12393
rect 10968 12384 11020 12436
rect 11244 12384 11296 12436
rect 11980 12384 12032 12436
rect 12256 12384 12308 12436
rect 3240 12316 3292 12368
rect 4160 12316 4212 12368
rect 6644 12316 6696 12368
rect 3332 12248 3384 12300
rect 3700 12248 3752 12300
rect 3884 12248 3936 12300
rect 4528 12291 4580 12300
rect 4528 12257 4537 12291
rect 4537 12257 4571 12291
rect 4571 12257 4580 12291
rect 4528 12248 4580 12257
rect 7288 12316 7340 12368
rect 8208 12316 8260 12368
rect 9220 12316 9272 12368
rect 9772 12316 9824 12368
rect 9864 12316 9916 12368
rect 12532 12316 12584 12368
rect 12900 12316 12952 12368
rect 12992 12316 13044 12368
rect 13360 12316 13412 12368
rect 7104 12291 7156 12300
rect 7104 12257 7113 12291
rect 7113 12257 7147 12291
rect 7147 12257 7156 12291
rect 7104 12248 7156 12257
rect 7748 12248 7800 12300
rect 10784 12248 10836 12300
rect 11060 12291 11112 12300
rect 11060 12257 11069 12291
rect 11069 12257 11103 12291
rect 11103 12257 11112 12291
rect 11060 12248 11112 12257
rect 12440 12248 12492 12300
rect 13176 12248 13228 12300
rect 1952 12180 2004 12232
rect 2136 12180 2188 12232
rect 2504 12223 2556 12232
rect 2504 12189 2538 12223
rect 2538 12189 2556 12223
rect 1492 12112 1544 12164
rect 2504 12180 2556 12189
rect 2872 12180 2924 12232
rect 4068 12180 4120 12232
rect 4712 12180 4764 12232
rect 4896 12180 4948 12232
rect 7656 12180 7708 12232
rect 8852 12180 8904 12232
rect 9220 12180 9272 12232
rect 1860 12087 1912 12096
rect 1860 12053 1869 12087
rect 1869 12053 1903 12087
rect 1903 12053 1912 12087
rect 1860 12044 1912 12053
rect 4160 12044 4212 12096
rect 4896 12044 4948 12096
rect 5356 12112 5408 12164
rect 6920 12112 6972 12164
rect 8300 12112 8352 12164
rect 12348 12180 12400 12232
rect 11336 12155 11388 12164
rect 11336 12121 11370 12155
rect 11370 12121 11388 12155
rect 11336 12112 11388 12121
rect 11796 12112 11848 12164
rect 13544 12384 13596 12436
rect 14280 12384 14332 12436
rect 15660 12384 15712 12436
rect 16396 12427 16448 12436
rect 16396 12393 16405 12427
rect 16405 12393 16439 12427
rect 16439 12393 16448 12427
rect 16396 12384 16448 12393
rect 18052 12427 18104 12436
rect 18052 12393 18061 12427
rect 18061 12393 18095 12427
rect 18095 12393 18104 12427
rect 18052 12384 18104 12393
rect 20628 12384 20680 12436
rect 20812 12384 20864 12436
rect 22284 12384 22336 12436
rect 16948 12291 17000 12300
rect 16948 12257 16957 12291
rect 16957 12257 16991 12291
rect 16991 12257 17000 12291
rect 16948 12248 17000 12257
rect 17960 12316 18012 12368
rect 20260 12316 20312 12368
rect 22560 12316 22612 12368
rect 17592 12248 17644 12300
rect 20352 12248 20404 12300
rect 22100 12248 22152 12300
rect 22376 12248 22428 12300
rect 13820 12180 13872 12232
rect 14832 12180 14884 12232
rect 15384 12180 15436 12232
rect 16212 12180 16264 12232
rect 18880 12223 18932 12232
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 20536 12223 20588 12232
rect 5632 12044 5684 12096
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 7012 12044 7064 12096
rect 8024 12044 8076 12096
rect 8208 12087 8260 12096
rect 8208 12053 8217 12087
rect 8217 12053 8251 12087
rect 8251 12053 8260 12087
rect 8208 12044 8260 12053
rect 8576 12044 8628 12096
rect 8668 12044 8720 12096
rect 9864 12087 9916 12096
rect 9864 12053 9873 12087
rect 9873 12053 9907 12087
rect 9907 12053 9916 12087
rect 9864 12044 9916 12053
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 10232 12087 10284 12096
rect 10232 12053 10241 12087
rect 10241 12053 10275 12087
rect 10275 12053 10284 12087
rect 10232 12044 10284 12053
rect 10324 12087 10376 12096
rect 10324 12053 10333 12087
rect 10333 12053 10367 12087
rect 10367 12053 10376 12087
rect 10324 12044 10376 12053
rect 10784 12044 10836 12096
rect 13452 12112 13504 12164
rect 14648 12112 14700 12164
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 12900 12044 12952 12096
rect 13084 12044 13136 12096
rect 13820 12087 13872 12096
rect 13820 12053 13829 12087
rect 13829 12053 13863 12087
rect 13863 12053 13872 12087
rect 13820 12044 13872 12053
rect 16120 12112 16172 12164
rect 16764 12155 16816 12164
rect 16764 12121 16773 12155
rect 16773 12121 16807 12155
rect 16807 12121 16816 12155
rect 16764 12112 16816 12121
rect 17040 12112 17092 12164
rect 15292 12044 15344 12096
rect 15384 12044 15436 12096
rect 15936 12087 15988 12096
rect 15936 12053 15945 12087
rect 15945 12053 15979 12087
rect 15979 12053 15988 12087
rect 15936 12044 15988 12053
rect 16028 12087 16080 12096
rect 16028 12053 16037 12087
rect 16037 12053 16071 12087
rect 16071 12053 16080 12087
rect 16028 12044 16080 12053
rect 17224 12044 17276 12096
rect 20168 12112 20220 12164
rect 20536 12189 20545 12223
rect 20545 12189 20579 12223
rect 20579 12189 20588 12223
rect 20536 12180 20588 12189
rect 21640 12180 21692 12232
rect 20444 12112 20496 12164
rect 21088 12155 21140 12164
rect 18420 12087 18472 12096
rect 18420 12053 18429 12087
rect 18429 12053 18463 12087
rect 18463 12053 18472 12087
rect 18420 12044 18472 12053
rect 19340 12044 19392 12096
rect 19892 12087 19944 12096
rect 19892 12053 19901 12087
rect 19901 12053 19935 12087
rect 19935 12053 19944 12087
rect 20260 12087 20312 12096
rect 19892 12044 19944 12053
rect 20260 12053 20269 12087
rect 20269 12053 20303 12087
rect 20303 12053 20312 12087
rect 20260 12044 20312 12053
rect 21088 12121 21097 12155
rect 21097 12121 21131 12155
rect 21131 12121 21140 12155
rect 21088 12112 21140 12121
rect 21456 12087 21508 12096
rect 21456 12053 21465 12087
rect 21465 12053 21499 12087
rect 21499 12053 21508 12087
rect 21456 12044 21508 12053
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 2320 11840 2372 11892
rect 2412 11840 2464 11892
rect 2688 11840 2740 11892
rect 3424 11840 3476 11892
rect 4344 11840 4396 11892
rect 5356 11883 5408 11892
rect 5356 11849 5365 11883
rect 5365 11849 5399 11883
rect 5399 11849 5408 11883
rect 5356 11840 5408 11849
rect 2780 11772 2832 11824
rect 2872 11772 2924 11824
rect 4804 11772 4856 11824
rect 5540 11772 5592 11824
rect 6184 11772 6236 11824
rect 7196 11840 7248 11892
rect 7748 11883 7800 11892
rect 2412 11704 2464 11756
rect 3424 11704 3476 11756
rect 4528 11747 4580 11756
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 3884 11679 3936 11688
rect 1860 11568 1912 11620
rect 1400 11500 1452 11552
rect 2504 11568 2556 11620
rect 3884 11645 3893 11679
rect 3893 11645 3927 11679
rect 3927 11645 3936 11679
rect 3884 11636 3936 11645
rect 4068 11611 4120 11620
rect 4068 11577 4077 11611
rect 4077 11577 4111 11611
rect 4111 11577 4120 11611
rect 4068 11568 4120 11577
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4988 11747 5040 11756
rect 4528 11704 4580 11713
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 7656 11815 7708 11824
rect 7656 11781 7665 11815
rect 7665 11781 7699 11815
rect 7699 11781 7708 11815
rect 7656 11772 7708 11781
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 8944 11772 8996 11824
rect 8024 11704 8076 11756
rect 9312 11772 9364 11824
rect 9772 11704 9824 11756
rect 11060 11772 11112 11824
rect 10508 11704 10560 11756
rect 11244 11840 11296 11892
rect 12532 11840 12584 11892
rect 12624 11840 12676 11892
rect 12992 11840 13044 11892
rect 15108 11883 15160 11892
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 16028 11840 16080 11892
rect 17132 11840 17184 11892
rect 17408 11840 17460 11892
rect 18236 11883 18288 11892
rect 18236 11849 18245 11883
rect 18245 11849 18279 11883
rect 18279 11849 18288 11883
rect 18236 11840 18288 11849
rect 20352 11883 20404 11892
rect 20352 11849 20361 11883
rect 20361 11849 20395 11883
rect 20395 11849 20404 11883
rect 20352 11840 20404 11849
rect 20444 11883 20496 11892
rect 20444 11849 20453 11883
rect 20453 11849 20487 11883
rect 20487 11849 20496 11883
rect 20444 11840 20496 11849
rect 22836 11840 22888 11892
rect 11428 11772 11480 11824
rect 12900 11772 12952 11824
rect 13176 11772 13228 11824
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 6736 11568 6788 11620
rect 3792 11500 3844 11552
rect 4712 11500 4764 11552
rect 6000 11500 6052 11552
rect 7012 11636 7064 11688
rect 7840 11500 7892 11552
rect 12348 11704 12400 11756
rect 12624 11704 12676 11756
rect 13360 11704 13412 11756
rect 13636 11704 13688 11756
rect 8484 11568 8536 11620
rect 8852 11500 8904 11552
rect 9864 11543 9916 11552
rect 9864 11509 9873 11543
rect 9873 11509 9907 11543
rect 9907 11509 9916 11543
rect 9864 11500 9916 11509
rect 11428 11568 11480 11620
rect 12164 11568 12216 11620
rect 12256 11568 12308 11620
rect 13176 11636 13228 11688
rect 14464 11772 14516 11824
rect 18328 11772 18380 11824
rect 15476 11704 15528 11756
rect 16396 11704 16448 11756
rect 16580 11704 16632 11756
rect 17500 11704 17552 11756
rect 17684 11704 17736 11756
rect 18052 11704 18104 11756
rect 18788 11772 18840 11824
rect 19340 11772 19392 11824
rect 21272 11772 21324 11824
rect 14280 11636 14332 11688
rect 14648 11679 14700 11688
rect 14648 11645 14657 11679
rect 14657 11645 14691 11679
rect 14691 11645 14700 11679
rect 14648 11636 14700 11645
rect 14924 11636 14976 11688
rect 15200 11636 15252 11688
rect 16212 11636 16264 11688
rect 16764 11636 16816 11688
rect 17592 11679 17644 11688
rect 14372 11568 14424 11620
rect 16120 11568 16172 11620
rect 17592 11645 17601 11679
rect 17601 11645 17635 11679
rect 17635 11645 17644 11679
rect 17592 11636 17644 11645
rect 17776 11679 17828 11688
rect 17776 11645 17785 11679
rect 17785 11645 17819 11679
rect 17819 11645 17828 11679
rect 17776 11636 17828 11645
rect 17684 11568 17736 11620
rect 11060 11500 11112 11552
rect 11612 11500 11664 11552
rect 12900 11500 12952 11552
rect 13268 11500 13320 11552
rect 15200 11543 15252 11552
rect 15200 11509 15209 11543
rect 15209 11509 15243 11543
rect 15243 11509 15252 11543
rect 16396 11543 16448 11552
rect 15200 11500 15252 11509
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16396 11500 16448 11509
rect 16856 11500 16908 11552
rect 17316 11500 17368 11552
rect 17408 11500 17460 11552
rect 18144 11500 18196 11552
rect 19064 11704 19116 11756
rect 20260 11704 20312 11756
rect 20812 11636 20864 11688
rect 21548 11679 21600 11688
rect 21548 11645 21557 11679
rect 21557 11645 21591 11679
rect 21591 11645 21600 11679
rect 21548 11636 21600 11645
rect 18972 11500 19024 11552
rect 19156 11500 19208 11552
rect 22744 11568 22796 11620
rect 22836 11568 22888 11620
rect 21364 11500 21416 11552
rect 22100 11500 22152 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1952 11296 2004 11348
rect 4436 11296 4488 11348
rect 5264 11296 5316 11348
rect 1676 11271 1728 11280
rect 1676 11237 1685 11271
rect 1685 11237 1719 11271
rect 1719 11237 1728 11271
rect 1676 11228 1728 11237
rect 3608 11271 3660 11280
rect 3608 11237 3617 11271
rect 3617 11237 3651 11271
rect 3651 11237 3660 11271
rect 3608 11228 3660 11237
rect 3332 11160 3384 11212
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 2504 11135 2556 11144
rect 2504 11101 2538 11135
rect 2538 11101 2556 11135
rect 1860 11067 1912 11076
rect 1860 11033 1869 11067
rect 1869 11033 1903 11067
rect 1903 11033 1912 11067
rect 1860 11024 1912 11033
rect 2044 11067 2096 11076
rect 2044 11033 2053 11067
rect 2053 11033 2087 11067
rect 2087 11033 2096 11067
rect 2044 11024 2096 11033
rect 2504 11092 2556 11101
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 4528 11203 4580 11212
rect 4528 11169 4537 11203
rect 4537 11169 4571 11203
rect 4571 11169 4580 11203
rect 5816 11296 5868 11348
rect 5632 11228 5684 11280
rect 7472 11296 7524 11348
rect 8760 11339 8812 11348
rect 8760 11305 8769 11339
rect 8769 11305 8803 11339
rect 8803 11305 8812 11339
rect 8760 11296 8812 11305
rect 7012 11228 7064 11280
rect 4528 11160 4580 11169
rect 6092 11203 6144 11212
rect 6092 11169 6101 11203
rect 6101 11169 6135 11203
rect 6135 11169 6144 11203
rect 6368 11203 6420 11212
rect 6092 11160 6144 11169
rect 6368 11169 6377 11203
rect 6377 11169 6411 11203
rect 6411 11169 6420 11203
rect 6368 11160 6420 11169
rect 6920 11092 6972 11144
rect 7104 11160 7156 11212
rect 9036 11160 9088 11212
rect 9128 11203 9180 11212
rect 9128 11169 9137 11203
rect 9137 11169 9171 11203
rect 9171 11169 9180 11203
rect 10692 11296 10744 11348
rect 11428 11296 11480 11348
rect 11704 11296 11756 11348
rect 12348 11339 12400 11348
rect 10876 11271 10928 11280
rect 10876 11237 10885 11271
rect 10885 11237 10919 11271
rect 10919 11237 10928 11271
rect 10876 11228 10928 11237
rect 12348 11305 12357 11339
rect 12357 11305 12391 11339
rect 12391 11305 12400 11339
rect 12348 11296 12400 11305
rect 13176 11339 13228 11348
rect 13176 11305 13185 11339
rect 13185 11305 13219 11339
rect 13219 11305 13228 11339
rect 13176 11296 13228 11305
rect 13360 11339 13412 11348
rect 13360 11305 13369 11339
rect 13369 11305 13403 11339
rect 13403 11305 13412 11339
rect 13360 11296 13412 11305
rect 13820 11339 13872 11348
rect 13820 11305 13829 11339
rect 13829 11305 13863 11339
rect 13863 11305 13872 11339
rect 13820 11296 13872 11305
rect 14464 11296 14516 11348
rect 14648 11296 14700 11348
rect 15476 11296 15528 11348
rect 15936 11296 15988 11348
rect 17132 11296 17184 11348
rect 17316 11296 17368 11348
rect 11796 11203 11848 11212
rect 9128 11160 9180 11169
rect 11796 11169 11805 11203
rect 11805 11169 11839 11203
rect 11839 11169 11848 11203
rect 11796 11160 11848 11169
rect 2964 11024 3016 11076
rect 3424 11024 3476 11076
rect 4528 11024 4580 11076
rect 4804 11067 4856 11076
rect 4804 11033 4838 11067
rect 4838 11033 4856 11067
rect 4804 11024 4856 11033
rect 5632 11024 5684 11076
rect 6368 11024 6420 11076
rect 6552 11024 6604 11076
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 8576 11092 8628 11144
rect 8944 11135 8996 11144
rect 8944 11101 8953 11135
rect 8953 11101 8987 11135
rect 8987 11101 8996 11135
rect 8944 11092 8996 11101
rect 3148 10956 3200 11008
rect 6184 10956 6236 11008
rect 7012 10956 7064 11008
rect 7564 11024 7616 11076
rect 8484 11024 8536 11076
rect 11704 11092 11756 11144
rect 12072 11092 12124 11144
rect 12348 11160 12400 11212
rect 17868 11296 17920 11348
rect 18052 11296 18104 11348
rect 12716 11092 12768 11144
rect 14464 11160 14516 11212
rect 15016 11160 15068 11212
rect 15200 11203 15252 11212
rect 15200 11169 15209 11203
rect 15209 11169 15243 11203
rect 15243 11169 15252 11203
rect 15200 11160 15252 11169
rect 15292 11203 15344 11212
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 16120 11203 16172 11212
rect 15292 11160 15344 11169
rect 16120 11169 16129 11203
rect 16129 11169 16163 11203
rect 16163 11169 16172 11203
rect 16120 11160 16172 11169
rect 13636 11067 13688 11076
rect 7656 10956 7708 11008
rect 8208 10956 8260 11008
rect 10508 10999 10560 11008
rect 10508 10965 10517 10999
rect 10517 10965 10551 10999
rect 10551 10965 10560 10999
rect 10508 10956 10560 10965
rect 10600 10999 10652 11008
rect 10600 10965 10609 10999
rect 10609 10965 10643 10999
rect 10643 10965 10652 10999
rect 11152 10999 11204 11008
rect 10600 10956 10652 10965
rect 11152 10965 11161 10999
rect 11161 10965 11195 10999
rect 11195 10965 11204 10999
rect 11152 10956 11204 10965
rect 11704 10956 11756 11008
rect 11980 10956 12032 11008
rect 13636 11033 13645 11067
rect 13645 11033 13679 11067
rect 13679 11033 13688 11067
rect 13636 11024 13688 11033
rect 13176 10956 13228 11008
rect 16028 11092 16080 11144
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 16856 11135 16908 11144
rect 16856 11101 16865 11135
rect 16865 11101 16899 11135
rect 16899 11101 16908 11135
rect 16856 11092 16908 11101
rect 15016 11024 15068 11076
rect 16948 11024 17000 11076
rect 17132 11160 17184 11212
rect 17684 11203 17736 11212
rect 17684 11169 17693 11203
rect 17693 11169 17727 11203
rect 17727 11169 17736 11203
rect 17684 11160 17736 11169
rect 18788 11296 18840 11348
rect 19064 11271 19116 11280
rect 19064 11237 19073 11271
rect 19073 11237 19107 11271
rect 19107 11237 19116 11271
rect 19064 11228 19116 11237
rect 19248 11228 19300 11280
rect 17316 11092 17368 11144
rect 17592 11024 17644 11076
rect 18696 11024 18748 11076
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 16028 10999 16080 11008
rect 16028 10965 16037 10999
rect 16037 10965 16071 10999
rect 16071 10965 16080 10999
rect 16028 10956 16080 10965
rect 16212 10956 16264 11008
rect 17316 10956 17368 11008
rect 18236 10956 18288 11008
rect 18512 10956 18564 11008
rect 21272 11203 21324 11212
rect 21272 11169 21281 11203
rect 21281 11169 21315 11203
rect 21315 11169 21324 11203
rect 21272 11160 21324 11169
rect 20352 11135 20404 11144
rect 20352 11101 20370 11135
rect 20370 11101 20404 11135
rect 20352 11092 20404 11101
rect 20720 11092 20772 11144
rect 19800 10956 19852 11008
rect 20352 10956 20404 11008
rect 20812 10956 20864 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 2504 10752 2556 10804
rect 2780 10752 2832 10804
rect 4804 10752 4856 10804
rect 5172 10752 5224 10804
rect 6552 10752 6604 10804
rect 6828 10752 6880 10804
rect 7564 10752 7616 10804
rect 7748 10752 7800 10804
rect 7932 10752 7984 10804
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 8392 10752 8444 10804
rect 8668 10752 8720 10804
rect 9772 10795 9824 10804
rect 9772 10761 9781 10795
rect 9781 10761 9815 10795
rect 9815 10761 9824 10795
rect 9772 10752 9824 10761
rect 10600 10752 10652 10804
rect 11888 10752 11940 10804
rect 12072 10752 12124 10804
rect 12348 10752 12400 10804
rect 13084 10752 13136 10804
rect 13544 10752 13596 10804
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 1768 10684 1820 10736
rect 1860 10616 1912 10668
rect 3608 10684 3660 10736
rect 2964 10591 3016 10600
rect 2964 10557 2973 10591
rect 2973 10557 3007 10591
rect 3007 10557 3016 10591
rect 2964 10548 3016 10557
rect 4344 10616 4396 10668
rect 5356 10616 5408 10668
rect 6736 10616 6788 10668
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 4252 10591 4304 10600
rect 4252 10557 4261 10591
rect 4261 10557 4295 10591
rect 4295 10557 4304 10591
rect 4252 10548 4304 10557
rect 5908 10548 5960 10600
rect 7380 10727 7432 10736
rect 7380 10693 7389 10727
rect 7389 10693 7423 10727
rect 7423 10693 7432 10727
rect 7380 10684 7432 10693
rect 7012 10616 7064 10668
rect 7288 10616 7340 10668
rect 7840 10616 7892 10668
rect 8024 10616 8076 10668
rect 8944 10684 8996 10736
rect 9036 10684 9088 10736
rect 9312 10684 9364 10736
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 2228 10412 2280 10464
rect 3424 10412 3476 10464
rect 6184 10480 6236 10532
rect 6460 10480 6512 10532
rect 7656 10480 7708 10532
rect 6000 10412 6052 10464
rect 6368 10412 6420 10464
rect 6828 10412 6880 10464
rect 7104 10412 7156 10464
rect 8024 10523 8076 10532
rect 8024 10489 8033 10523
rect 8033 10489 8067 10523
rect 8067 10489 8076 10523
rect 8024 10480 8076 10489
rect 7932 10412 7984 10464
rect 9588 10616 9640 10668
rect 8300 10548 8352 10600
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 9772 10480 9824 10532
rect 10324 10548 10376 10600
rect 11704 10684 11756 10736
rect 11980 10684 12032 10736
rect 12164 10684 12216 10736
rect 12716 10684 12768 10736
rect 15936 10752 15988 10804
rect 16120 10795 16172 10804
rect 16120 10761 16129 10795
rect 16129 10761 16163 10795
rect 16163 10761 16172 10795
rect 16120 10752 16172 10761
rect 16948 10752 17000 10804
rect 17592 10752 17644 10804
rect 18052 10795 18104 10804
rect 18052 10761 18061 10795
rect 18061 10761 18095 10795
rect 18095 10761 18104 10795
rect 18052 10752 18104 10761
rect 18420 10752 18472 10804
rect 19892 10752 19944 10804
rect 20260 10795 20312 10804
rect 20260 10761 20269 10795
rect 20269 10761 20303 10795
rect 20303 10761 20312 10795
rect 20260 10752 20312 10761
rect 15200 10684 15252 10736
rect 16212 10684 16264 10736
rect 11152 10616 11204 10668
rect 12256 10616 12308 10668
rect 12440 10616 12492 10668
rect 14280 10616 14332 10668
rect 15752 10616 15804 10668
rect 16948 10616 17000 10668
rect 17868 10684 17920 10736
rect 17960 10684 18012 10736
rect 11244 10548 11296 10600
rect 12072 10548 12124 10600
rect 14648 10548 14700 10600
rect 15936 10548 15988 10600
rect 16856 10548 16908 10600
rect 17316 10591 17368 10600
rect 17316 10557 17325 10591
rect 17325 10557 17359 10591
rect 17359 10557 17368 10591
rect 17316 10548 17368 10557
rect 18604 10616 18656 10668
rect 18972 10659 19024 10668
rect 18328 10548 18380 10600
rect 18972 10625 18981 10659
rect 18981 10625 19015 10659
rect 19015 10625 19024 10659
rect 18972 10616 19024 10625
rect 18788 10548 18840 10600
rect 20720 10684 20772 10736
rect 21180 10684 21232 10736
rect 19800 10659 19852 10668
rect 19800 10625 19809 10659
rect 19809 10625 19843 10659
rect 19843 10625 19852 10659
rect 19800 10616 19852 10625
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 21456 10659 21508 10668
rect 21456 10625 21465 10659
rect 21465 10625 21499 10659
rect 21499 10625 21508 10659
rect 21456 10616 21508 10625
rect 19248 10548 19300 10600
rect 10232 10412 10284 10464
rect 10324 10412 10376 10464
rect 10416 10412 10468 10464
rect 10692 10412 10744 10464
rect 11704 10412 11756 10464
rect 12256 10455 12308 10464
rect 12256 10421 12265 10455
rect 12265 10421 12299 10455
rect 12299 10421 12308 10455
rect 12256 10412 12308 10421
rect 14464 10480 14516 10532
rect 13728 10455 13780 10464
rect 13728 10421 13737 10455
rect 13737 10421 13771 10455
rect 13771 10421 13780 10455
rect 13728 10412 13780 10421
rect 16120 10412 16172 10464
rect 16396 10455 16448 10464
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 17776 10480 17828 10532
rect 20168 10548 20220 10600
rect 20260 10548 20312 10600
rect 20628 10412 20680 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 2964 10208 3016 10260
rect 1492 10072 1544 10124
rect 2044 10072 2096 10124
rect 4988 10208 5040 10260
rect 5540 10208 5592 10260
rect 7196 10208 7248 10260
rect 3608 10115 3660 10124
rect 3608 10081 3617 10115
rect 3617 10081 3651 10115
rect 3651 10081 3660 10115
rect 3608 10072 3660 10081
rect 1952 9936 2004 9988
rect 2964 9979 3016 9988
rect 2964 9945 2982 9979
rect 2982 9945 3016 9979
rect 2964 9936 3016 9945
rect 1860 9911 1912 9920
rect 1860 9877 1869 9911
rect 1869 9877 1903 9911
rect 1903 9877 1912 9911
rect 1860 9868 1912 9877
rect 2044 9868 2096 9920
rect 5172 10072 5224 10124
rect 5448 10072 5500 10124
rect 7104 10183 7156 10192
rect 7104 10149 7113 10183
rect 7113 10149 7147 10183
rect 7147 10149 7156 10183
rect 7104 10140 7156 10149
rect 6368 10072 6420 10124
rect 6552 10072 6604 10124
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 4068 10047 4120 10056
rect 3792 10004 3844 10013
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4436 10004 4488 10056
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 5448 9936 5500 9988
rect 10876 10208 10928 10260
rect 9404 10140 9456 10192
rect 9680 10140 9732 10192
rect 8392 10072 8444 10124
rect 10508 10072 10560 10124
rect 10600 10072 10652 10124
rect 12164 10140 12216 10192
rect 14372 10208 14424 10260
rect 16028 10208 16080 10260
rect 16212 10251 16264 10260
rect 16212 10217 16221 10251
rect 16221 10217 16255 10251
rect 16255 10217 16264 10251
rect 16212 10208 16264 10217
rect 12808 10072 12860 10124
rect 13728 10072 13780 10124
rect 14188 10115 14240 10124
rect 14188 10081 14197 10115
rect 14197 10081 14231 10115
rect 14231 10081 14240 10115
rect 14188 10072 14240 10081
rect 15016 10115 15068 10124
rect 15016 10081 15025 10115
rect 15025 10081 15059 10115
rect 15059 10081 15068 10115
rect 15016 10072 15068 10081
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 8024 10004 8076 10056
rect 8668 10004 8720 10056
rect 9036 10004 9088 10056
rect 4436 9868 4488 9920
rect 5540 9868 5592 9920
rect 5816 9868 5868 9920
rect 6276 9868 6328 9920
rect 7840 9936 7892 9988
rect 8852 9936 8904 9988
rect 7380 9868 7432 9920
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 11888 10004 11940 10056
rect 12900 10004 12952 10056
rect 14556 10004 14608 10056
rect 11520 9979 11572 9988
rect 11520 9945 11529 9979
rect 11529 9945 11563 9979
rect 11563 9945 11572 9979
rect 11520 9936 11572 9945
rect 9220 9868 9272 9920
rect 9496 9868 9548 9920
rect 9864 9868 9916 9920
rect 10140 9911 10192 9920
rect 10140 9877 10149 9911
rect 10149 9877 10183 9911
rect 10183 9877 10192 9911
rect 10140 9868 10192 9877
rect 10692 9911 10744 9920
rect 10692 9877 10701 9911
rect 10701 9877 10735 9911
rect 10735 9877 10744 9911
rect 10692 9868 10744 9877
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 11152 9911 11204 9920
rect 11152 9877 11161 9911
rect 11161 9877 11195 9911
rect 11195 9877 11204 9911
rect 12164 9911 12216 9920
rect 11152 9868 11204 9877
rect 12164 9877 12173 9911
rect 12173 9877 12207 9911
rect 12207 9877 12216 9911
rect 12164 9868 12216 9877
rect 14188 9936 14240 9988
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 16212 10004 16264 10056
rect 17684 10208 17736 10260
rect 18696 10251 18748 10260
rect 18696 10217 18705 10251
rect 18705 10217 18739 10251
rect 18739 10217 18748 10251
rect 18696 10208 18748 10217
rect 19616 10208 19668 10260
rect 19892 10208 19944 10260
rect 20260 10251 20312 10260
rect 20260 10217 20269 10251
rect 20269 10217 20303 10251
rect 20303 10217 20312 10251
rect 20260 10208 20312 10217
rect 17316 10115 17368 10124
rect 17316 10081 17325 10115
rect 17325 10081 17359 10115
rect 17359 10081 17368 10115
rect 17316 10072 17368 10081
rect 19340 10140 19392 10192
rect 20444 10140 20496 10192
rect 21272 10140 21324 10192
rect 19616 10115 19668 10124
rect 19616 10081 19625 10115
rect 19625 10081 19659 10115
rect 19659 10081 19668 10115
rect 19616 10072 19668 10081
rect 19708 10004 19760 10056
rect 20812 10072 20864 10124
rect 20996 10115 21048 10124
rect 20996 10081 21005 10115
rect 21005 10081 21039 10115
rect 21039 10081 21048 10115
rect 20996 10072 21048 10081
rect 20628 10004 20680 10056
rect 17684 9936 17736 9988
rect 17776 9936 17828 9988
rect 18972 9979 19024 9988
rect 18972 9945 18981 9979
rect 18981 9945 19015 9979
rect 19015 9945 19024 9979
rect 18972 9936 19024 9945
rect 20352 9936 20404 9988
rect 20444 9979 20496 9988
rect 20444 9945 20453 9979
rect 20453 9945 20487 9979
rect 20487 9945 20496 9979
rect 20444 9936 20496 9945
rect 12624 9868 12676 9920
rect 13912 9868 13964 9920
rect 14740 9868 14792 9920
rect 15016 9868 15068 9920
rect 15476 9868 15528 9920
rect 16304 9868 16356 9920
rect 17132 9868 17184 9920
rect 17868 9868 17920 9920
rect 19156 9868 19208 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 1768 9664 1820 9716
rect 2136 9664 2188 9716
rect 3332 9664 3384 9716
rect 4344 9664 4396 9716
rect 5356 9664 5408 9716
rect 6184 9664 6236 9716
rect 3792 9639 3844 9648
rect 3792 9605 3810 9639
rect 3810 9605 3844 9639
rect 3792 9596 3844 9605
rect 5540 9596 5592 9648
rect 7104 9664 7156 9716
rect 7748 9664 7800 9716
rect 8392 9664 8444 9716
rect 9772 9664 9824 9716
rect 10784 9664 10836 9716
rect 11060 9664 11112 9716
rect 11704 9664 11756 9716
rect 11888 9664 11940 9716
rect 12256 9664 12308 9716
rect 12808 9664 12860 9716
rect 13084 9664 13136 9716
rect 19156 9664 19208 9716
rect 19800 9664 19852 9716
rect 20168 9664 20220 9716
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 4528 9528 4580 9580
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 2136 9460 2188 9512
rect 4252 9460 4304 9512
rect 4344 9460 4396 9512
rect 4896 9460 4948 9512
rect 2412 9435 2464 9444
rect 2412 9401 2421 9435
rect 2421 9401 2455 9435
rect 2455 9401 2464 9435
rect 2412 9392 2464 9401
rect 1676 9324 1728 9376
rect 2964 9392 3016 9444
rect 2872 9324 2924 9376
rect 3056 9324 3108 9376
rect 4804 9392 4856 9444
rect 5172 9503 5224 9512
rect 5172 9469 5181 9503
rect 5181 9469 5215 9503
rect 5215 9469 5224 9503
rect 5172 9460 5224 9469
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 7840 9596 7892 9648
rect 6828 9571 6880 9580
rect 5816 9528 5868 9537
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 6920 9528 6972 9580
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 7932 9528 7984 9580
rect 8392 9571 8444 9580
rect 5908 9503 5960 9512
rect 5908 9469 5917 9503
rect 5917 9469 5951 9503
rect 5951 9469 5960 9503
rect 5908 9460 5960 9469
rect 6276 9460 6328 9512
rect 7380 9460 7432 9512
rect 8392 9537 8415 9571
rect 8415 9537 8444 9571
rect 8392 9528 8444 9537
rect 9312 9596 9364 9648
rect 9588 9528 9640 9580
rect 9772 9528 9824 9580
rect 11704 9528 11756 9580
rect 12440 9596 12492 9648
rect 13728 9639 13780 9648
rect 12532 9528 12584 9580
rect 4344 9367 4396 9376
rect 4344 9333 4353 9367
rect 4353 9333 4387 9367
rect 4387 9333 4396 9367
rect 4344 9324 4396 9333
rect 7564 9324 7616 9376
rect 7932 9324 7984 9376
rect 9680 9324 9732 9376
rect 10508 9460 10560 9512
rect 11796 9503 11848 9512
rect 11796 9469 11805 9503
rect 11805 9469 11839 9503
rect 11839 9469 11848 9503
rect 11796 9460 11848 9469
rect 12716 9528 12768 9580
rect 13176 9528 13228 9580
rect 13728 9605 13762 9639
rect 13762 9605 13780 9639
rect 13728 9596 13780 9605
rect 14464 9596 14516 9648
rect 17592 9639 17644 9648
rect 17592 9605 17604 9639
rect 17604 9605 17644 9639
rect 17592 9596 17644 9605
rect 17684 9596 17736 9648
rect 17868 9596 17920 9648
rect 20444 9596 20496 9648
rect 20996 9596 21048 9648
rect 21272 9596 21324 9648
rect 14188 9528 14240 9580
rect 14556 9528 14608 9580
rect 17040 9528 17092 9580
rect 17132 9528 17184 9580
rect 17316 9571 17368 9580
rect 17316 9537 17325 9571
rect 17325 9537 17359 9571
rect 17359 9537 17368 9571
rect 17316 9528 17368 9537
rect 13084 9460 13136 9512
rect 12164 9392 12216 9444
rect 13452 9503 13504 9512
rect 13452 9469 13461 9503
rect 13461 9469 13495 9503
rect 13495 9469 13504 9503
rect 13452 9460 13504 9469
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 15476 9460 15528 9512
rect 15936 9503 15988 9512
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 15936 9460 15988 9469
rect 13360 9392 13412 9444
rect 14924 9392 14976 9444
rect 16672 9460 16724 9512
rect 17132 9392 17184 9444
rect 19340 9528 19392 9580
rect 19432 9571 19484 9580
rect 19432 9537 19441 9571
rect 19441 9537 19475 9571
rect 19475 9537 19484 9571
rect 19432 9528 19484 9537
rect 19708 9528 19760 9580
rect 19800 9528 19852 9580
rect 19616 9392 19668 9444
rect 20260 9460 20312 9512
rect 20444 9460 20496 9512
rect 20812 9503 20864 9512
rect 20812 9469 20821 9503
rect 20821 9469 20855 9503
rect 20855 9469 20864 9503
rect 20812 9460 20864 9469
rect 20628 9392 20680 9444
rect 21088 9392 21140 9444
rect 10416 9324 10468 9376
rect 12716 9324 12768 9376
rect 14740 9324 14792 9376
rect 15292 9324 15344 9376
rect 16672 9367 16724 9376
rect 16672 9333 16681 9367
rect 16681 9333 16715 9367
rect 16715 9333 16724 9367
rect 16672 9324 16724 9333
rect 16764 9324 16816 9376
rect 17224 9324 17276 9376
rect 18788 9324 18840 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 2136 9163 2188 9172
rect 2136 9129 2145 9163
rect 2145 9129 2179 9163
rect 2179 9129 2188 9163
rect 2136 9120 2188 9129
rect 3424 9120 3476 9172
rect 3884 9120 3936 9172
rect 4160 9120 4212 9172
rect 2504 9052 2556 9104
rect 2688 9052 2740 9104
rect 3976 9052 4028 9104
rect 1676 8984 1728 9036
rect 2412 8984 2464 9036
rect 4068 8984 4120 9036
rect 5172 9052 5224 9104
rect 2688 8916 2740 8968
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 2964 8848 3016 8900
rect 5908 9120 5960 9172
rect 6644 9120 6696 9172
rect 7380 9163 7432 9172
rect 7380 9129 7389 9163
rect 7389 9129 7423 9163
rect 7423 9129 7432 9163
rect 7380 9120 7432 9129
rect 7748 9120 7800 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9128 9120 9180 9129
rect 9588 9120 9640 9172
rect 11060 9120 11112 9172
rect 13084 9163 13136 9172
rect 13084 9129 13093 9163
rect 13093 9129 13127 9163
rect 13127 9129 13136 9163
rect 13084 9120 13136 9129
rect 13176 9163 13228 9172
rect 13176 9129 13185 9163
rect 13185 9129 13219 9163
rect 13219 9129 13228 9163
rect 13176 9120 13228 9129
rect 13820 9120 13872 9172
rect 14556 9163 14608 9172
rect 14556 9129 14565 9163
rect 14565 9129 14599 9163
rect 14599 9129 14608 9163
rect 14556 9120 14608 9129
rect 15936 9120 15988 9172
rect 10600 9052 10652 9104
rect 11704 9052 11756 9104
rect 5356 8984 5408 9036
rect 6276 9027 6328 9036
rect 6276 8993 6285 9027
rect 6285 8993 6319 9027
rect 6319 8993 6328 9027
rect 6276 8984 6328 8993
rect 6644 8984 6696 9036
rect 6736 8984 6788 9036
rect 10508 8984 10560 9036
rect 14464 9052 14516 9104
rect 12624 9027 12676 9036
rect 12624 8993 12633 9027
rect 12633 8993 12667 9027
rect 12667 8993 12676 9027
rect 12624 8984 12676 8993
rect 5172 8916 5224 8968
rect 5264 8959 5316 8968
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 6092 8959 6144 8968
rect 5264 8916 5316 8925
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 6552 8916 6604 8968
rect 7472 8916 7524 8968
rect 7748 8916 7800 8968
rect 8668 8916 8720 8968
rect 9588 8916 9640 8968
rect 11152 8916 11204 8968
rect 11704 8959 11756 8968
rect 11704 8925 11713 8959
rect 11713 8925 11747 8959
rect 11747 8925 11756 8959
rect 11704 8916 11756 8925
rect 12532 8916 12584 8968
rect 13360 8984 13412 9036
rect 14280 8984 14332 9036
rect 17040 9120 17092 9172
rect 18880 9120 18932 9172
rect 20720 9163 20772 9172
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 17500 9052 17552 9104
rect 18052 9052 18104 9104
rect 12900 8916 12952 8968
rect 13728 8916 13780 8968
rect 15476 8916 15528 8968
rect 16304 8959 16356 8968
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 17040 8916 17092 8968
rect 20628 8984 20680 9036
rect 18880 8959 18932 8968
rect 2504 8780 2556 8832
rect 3332 8780 3384 8832
rect 4804 8780 4856 8832
rect 5540 8780 5592 8832
rect 7932 8848 7984 8900
rect 9680 8848 9732 8900
rect 9864 8891 9916 8900
rect 9864 8857 9873 8891
rect 9873 8857 9907 8891
rect 9907 8857 9916 8891
rect 9864 8848 9916 8857
rect 6828 8780 6880 8832
rect 8024 8780 8076 8832
rect 9496 8780 9548 8832
rect 12256 8848 12308 8900
rect 13176 8780 13228 8832
rect 13452 8780 13504 8832
rect 14096 8780 14148 8832
rect 14556 8780 14608 8832
rect 15108 8891 15160 8900
rect 15108 8857 15142 8891
rect 15142 8857 15160 8891
rect 18880 8925 18889 8959
rect 18889 8925 18923 8959
rect 18923 8925 18932 8959
rect 18880 8916 18932 8925
rect 19064 8916 19116 8968
rect 19340 8916 19392 8968
rect 19524 8959 19576 8968
rect 19524 8925 19558 8959
rect 19558 8925 19576 8959
rect 19524 8916 19576 8925
rect 15108 8848 15160 8857
rect 19432 8848 19484 8900
rect 17684 8823 17736 8832
rect 17684 8789 17693 8823
rect 17693 8789 17727 8823
rect 17727 8789 17736 8823
rect 17684 8780 17736 8789
rect 18144 8823 18196 8832
rect 18144 8789 18153 8823
rect 18153 8789 18187 8823
rect 18187 8789 18196 8823
rect 18144 8780 18196 8789
rect 19340 8780 19392 8832
rect 20536 8780 20588 8832
rect 21088 8823 21140 8832
rect 21088 8789 21097 8823
rect 21097 8789 21131 8823
rect 21131 8789 21140 8823
rect 21088 8780 21140 8789
rect 21180 8823 21232 8832
rect 21180 8789 21189 8823
rect 21189 8789 21223 8823
rect 21223 8789 21232 8823
rect 21180 8780 21232 8789
rect 22008 8780 22060 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2136 8576 2188 8628
rect 4896 8576 4948 8628
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 5264 8576 5316 8628
rect 6276 8576 6328 8628
rect 6644 8576 6696 8628
rect 7288 8576 7340 8628
rect 8116 8576 8168 8628
rect 8852 8576 8904 8628
rect 4620 8508 4672 8560
rect 6000 8508 6052 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 2872 8440 2924 8492
rect 3240 8440 3292 8492
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 2412 8415 2464 8424
rect 2412 8381 2421 8415
rect 2421 8381 2455 8415
rect 2455 8381 2464 8415
rect 2412 8372 2464 8381
rect 2596 8372 2648 8424
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2964 8415 3016 8424
rect 2780 8372 2832 8381
rect 2964 8381 2973 8415
rect 2973 8381 3007 8415
rect 3007 8381 3016 8415
rect 2964 8372 3016 8381
rect 3884 8372 3936 8424
rect 1860 8279 1912 8288
rect 1860 8245 1869 8279
rect 1869 8245 1903 8279
rect 1903 8245 1912 8279
rect 1860 8236 1912 8245
rect 2872 8236 2924 8288
rect 4068 8236 4120 8288
rect 5448 8372 5500 8424
rect 6736 8440 6788 8492
rect 6552 8372 6604 8424
rect 8944 8508 8996 8560
rect 9404 8576 9456 8628
rect 9680 8576 9732 8628
rect 10048 8576 10100 8628
rect 11796 8576 11848 8628
rect 12716 8619 12768 8628
rect 12716 8585 12725 8619
rect 12725 8585 12759 8619
rect 12759 8585 12768 8619
rect 12716 8576 12768 8585
rect 13176 8576 13228 8628
rect 13728 8576 13780 8628
rect 14004 8576 14056 8628
rect 14924 8619 14976 8628
rect 14924 8585 14933 8619
rect 14933 8585 14967 8619
rect 14967 8585 14976 8619
rect 14924 8576 14976 8585
rect 15292 8576 15344 8628
rect 17132 8576 17184 8628
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 18144 8576 18196 8628
rect 19432 8619 19484 8628
rect 19432 8585 19441 8619
rect 19441 8585 19475 8619
rect 19475 8585 19484 8619
rect 19432 8576 19484 8585
rect 19708 8576 19760 8628
rect 20352 8576 20404 8628
rect 20720 8576 20772 8628
rect 7748 8415 7800 8424
rect 7748 8381 7757 8415
rect 7757 8381 7791 8415
rect 7791 8381 7800 8415
rect 7748 8372 7800 8381
rect 9496 8440 9548 8492
rect 10600 8508 10652 8560
rect 10876 8508 10928 8560
rect 12256 8508 12308 8560
rect 11336 8440 11388 8492
rect 12164 8483 12216 8492
rect 12164 8449 12173 8483
rect 12173 8449 12207 8483
rect 12207 8449 12216 8483
rect 12164 8440 12216 8449
rect 12992 8440 13044 8492
rect 4804 8304 4856 8356
rect 5172 8236 5224 8288
rect 8116 8304 8168 8356
rect 8668 8372 8720 8424
rect 11704 8372 11756 8424
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 7472 8236 7524 8288
rect 7564 8236 7616 8288
rect 9588 8304 9640 8356
rect 11152 8304 11204 8356
rect 12440 8372 12492 8424
rect 13176 8372 13228 8424
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 15476 8508 15528 8560
rect 17960 8508 18012 8560
rect 18972 8551 19024 8560
rect 18972 8517 18990 8551
rect 18990 8517 19024 8551
rect 18972 8508 19024 8517
rect 19156 8508 19208 8560
rect 21272 8508 21324 8560
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 13544 8372 13596 8381
rect 15016 8415 15068 8424
rect 13084 8347 13136 8356
rect 13084 8313 13093 8347
rect 13093 8313 13127 8347
rect 13127 8313 13136 8347
rect 13084 8304 13136 8313
rect 13820 8347 13872 8356
rect 13820 8313 13829 8347
rect 13829 8313 13863 8347
rect 13863 8313 13872 8347
rect 15016 8381 15025 8415
rect 15025 8381 15059 8415
rect 15059 8381 15068 8415
rect 15016 8372 15068 8381
rect 15936 8415 15988 8424
rect 15936 8381 15945 8415
rect 15945 8381 15979 8415
rect 15979 8381 15988 8415
rect 15936 8372 15988 8381
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 17500 8440 17552 8492
rect 19616 8440 19668 8492
rect 19892 8483 19944 8492
rect 19892 8449 19901 8483
rect 19901 8449 19935 8483
rect 19935 8449 19944 8483
rect 19892 8440 19944 8449
rect 16304 8372 16356 8424
rect 17040 8372 17092 8424
rect 17684 8372 17736 8424
rect 19340 8372 19392 8424
rect 20444 8372 20496 8424
rect 20720 8372 20772 8424
rect 21364 8372 21416 8424
rect 13820 8304 13872 8313
rect 15108 8304 15160 8356
rect 15200 8304 15252 8356
rect 17132 8304 17184 8356
rect 17592 8304 17644 8356
rect 9036 8236 9088 8288
rect 9956 8236 10008 8288
rect 11796 8279 11848 8288
rect 11796 8245 11805 8279
rect 11805 8245 11839 8279
rect 11839 8245 11848 8279
rect 11796 8236 11848 8245
rect 12992 8236 13044 8288
rect 14556 8236 14608 8288
rect 17224 8236 17276 8288
rect 17500 8236 17552 8288
rect 17684 8236 17736 8288
rect 21364 8279 21416 8288
rect 21364 8245 21373 8279
rect 21373 8245 21407 8279
rect 21407 8245 21416 8279
rect 21364 8236 21416 8245
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 2044 8032 2096 8084
rect 2964 8032 3016 8084
rect 4896 8032 4948 8084
rect 5816 8032 5868 8084
rect 6092 8075 6144 8084
rect 20 7964 72 8016
rect 940 7964 992 8016
rect 1124 7964 1176 8016
rect 1676 7896 1728 7948
rect 1860 7896 1912 7948
rect 3148 7964 3200 8016
rect 5356 7964 5408 8016
rect 6092 8041 6101 8075
rect 6101 8041 6135 8075
rect 6135 8041 6144 8075
rect 6092 8032 6144 8041
rect 7380 8032 7432 8084
rect 2964 7896 3016 7948
rect 3608 7896 3660 7948
rect 4160 7896 4212 7948
rect 7288 7964 7340 8016
rect 7472 7964 7524 8016
rect 1492 7828 1544 7880
rect 2872 7828 2924 7880
rect 3976 7828 4028 7880
rect 4068 7828 4120 7880
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 5356 7828 5408 7880
rect 5724 7828 5776 7880
rect 6828 7896 6880 7948
rect 8024 7896 8076 7948
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 7564 7828 7616 7880
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 10416 8032 10468 8084
rect 10784 8032 10836 8084
rect 11152 8032 11204 8084
rect 11704 8032 11756 8084
rect 9036 7964 9088 8016
rect 9772 7964 9824 8016
rect 10140 7964 10192 8016
rect 10876 7964 10928 8016
rect 8668 7896 8720 7948
rect 9404 7896 9456 7948
rect 9680 7896 9732 7948
rect 10048 7896 10100 7948
rect 10600 7896 10652 7948
rect 12992 8032 13044 8084
rect 2504 7760 2556 7812
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 2044 7735 2096 7744
rect 2044 7701 2053 7735
rect 2053 7701 2087 7735
rect 2087 7701 2096 7735
rect 2044 7692 2096 7701
rect 3700 7692 3752 7744
rect 3884 7692 3936 7744
rect 4712 7760 4764 7812
rect 8116 7760 8168 7812
rect 5080 7692 5132 7744
rect 5632 7735 5684 7744
rect 5632 7701 5641 7735
rect 5641 7701 5675 7735
rect 5675 7701 5684 7735
rect 5632 7692 5684 7701
rect 5816 7692 5868 7744
rect 7012 7692 7064 7744
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 7840 7692 7892 7744
rect 8024 7692 8076 7744
rect 8852 7760 8904 7812
rect 9128 7828 9180 7880
rect 10692 7828 10744 7880
rect 11796 7828 11848 7880
rect 14004 8032 14056 8084
rect 15200 8032 15252 8084
rect 16212 8032 16264 8084
rect 17408 8032 17460 8084
rect 18880 8032 18932 8084
rect 20168 8075 20220 8084
rect 20168 8041 20177 8075
rect 20177 8041 20211 8075
rect 20211 8041 20220 8075
rect 20168 8032 20220 8041
rect 21088 8032 21140 8084
rect 21456 8075 21508 8084
rect 21456 8041 21465 8075
rect 21465 8041 21499 8075
rect 21499 8041 21508 8075
rect 21456 8032 21508 8041
rect 15108 7964 15160 8016
rect 17592 8007 17644 8016
rect 14740 7939 14792 7948
rect 9220 7760 9272 7812
rect 8668 7692 8720 7744
rect 10232 7692 10284 7744
rect 12348 7760 12400 7812
rect 14740 7905 14749 7939
rect 14749 7905 14783 7939
rect 14783 7905 14792 7939
rect 14740 7896 14792 7905
rect 17132 7896 17184 7948
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 15016 7828 15068 7880
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 17316 7828 17368 7880
rect 17592 7973 17601 8007
rect 17601 7973 17635 8007
rect 17635 7973 17644 8007
rect 17592 7964 17644 7973
rect 18972 7964 19024 8016
rect 20260 8007 20312 8016
rect 17500 7896 17552 7948
rect 20260 7973 20269 8007
rect 20269 7973 20303 8007
rect 20303 7973 20312 8007
rect 20260 7964 20312 7973
rect 20444 7964 20496 8016
rect 20168 7896 20220 7948
rect 20720 7939 20772 7948
rect 20720 7905 20729 7939
rect 20729 7905 20763 7939
rect 20763 7905 20772 7939
rect 20720 7896 20772 7905
rect 21456 7896 21508 7948
rect 21732 7896 21784 7948
rect 22468 7896 22520 7948
rect 22836 7896 22888 7948
rect 17776 7828 17828 7880
rect 20444 7871 20496 7880
rect 15844 7803 15896 7812
rect 15844 7769 15853 7803
rect 15853 7769 15887 7803
rect 15887 7769 15896 7803
rect 15844 7760 15896 7769
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 18512 7760 18564 7812
rect 18696 7760 18748 7812
rect 22836 7760 22888 7812
rect 10968 7735 11020 7744
rect 10968 7701 10977 7735
rect 10977 7701 11011 7735
rect 11011 7701 11020 7735
rect 10968 7692 11020 7701
rect 11060 7692 11112 7744
rect 11796 7692 11848 7744
rect 12256 7692 12308 7744
rect 13084 7692 13136 7744
rect 14464 7692 14516 7744
rect 14556 7692 14608 7744
rect 15016 7735 15068 7744
rect 15016 7701 15025 7735
rect 15025 7701 15059 7735
rect 15059 7701 15068 7735
rect 15016 7692 15068 7701
rect 15384 7735 15436 7744
rect 15384 7701 15393 7735
rect 15393 7701 15427 7735
rect 15427 7701 15436 7735
rect 15384 7692 15436 7701
rect 18788 7692 18840 7744
rect 19340 7692 19392 7744
rect 19708 7735 19760 7744
rect 19708 7701 19717 7735
rect 19717 7701 19751 7735
rect 19751 7701 19760 7735
rect 19708 7692 19760 7701
rect 21272 7692 21324 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 1768 7488 1820 7540
rect 2504 7488 2556 7540
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 4252 7531 4304 7540
rect 2780 7488 2832 7497
rect 4252 7497 4261 7531
rect 4261 7497 4295 7531
rect 4295 7497 4304 7531
rect 4252 7488 4304 7497
rect 4712 7531 4764 7540
rect 4712 7497 4721 7531
rect 4721 7497 4755 7531
rect 4755 7497 4764 7531
rect 4712 7488 4764 7497
rect 6736 7488 6788 7540
rect 7564 7531 7616 7540
rect 940 7420 992 7472
rect 1860 7284 1912 7336
rect 2412 7284 2464 7336
rect 1676 7259 1728 7268
rect 1676 7225 1685 7259
rect 1685 7225 1719 7259
rect 1719 7225 1728 7259
rect 1676 7216 1728 7225
rect 2872 7420 2924 7472
rect 7564 7497 7573 7531
rect 7573 7497 7607 7531
rect 7607 7497 7616 7531
rect 7564 7488 7616 7497
rect 8024 7488 8076 7540
rect 9036 7488 9088 7540
rect 10232 7488 10284 7540
rect 2964 7352 3016 7404
rect 3608 7352 3660 7404
rect 4068 7352 4120 7404
rect 4252 7352 4304 7404
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 4712 7352 4764 7404
rect 4896 7352 4948 7404
rect 5448 7352 5500 7404
rect 1768 7191 1820 7200
rect 1768 7157 1777 7191
rect 1777 7157 1811 7191
rect 1811 7157 1820 7191
rect 1768 7148 1820 7157
rect 2780 7148 2832 7200
rect 4436 7216 4488 7268
rect 7380 7352 7432 7404
rect 8116 7420 8168 7472
rect 8392 7420 8444 7472
rect 8668 7420 8720 7472
rect 8852 7420 8904 7472
rect 10048 7420 10100 7472
rect 10600 7420 10652 7472
rect 6552 7284 6604 7336
rect 7840 7327 7892 7336
rect 4344 7148 4396 7200
rect 4712 7148 4764 7200
rect 5172 7148 5224 7200
rect 5540 7148 5592 7200
rect 5816 7148 5868 7200
rect 7380 7216 7432 7268
rect 6920 7148 6972 7200
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 7840 7293 7849 7327
rect 7849 7293 7883 7327
rect 7883 7293 7892 7327
rect 7840 7284 7892 7293
rect 10140 7352 10192 7404
rect 8024 7216 8076 7268
rect 9404 7284 9456 7336
rect 10784 7420 10836 7472
rect 11152 7420 11204 7472
rect 11060 7352 11112 7404
rect 11796 7488 11848 7540
rect 12164 7531 12216 7540
rect 12164 7497 12173 7531
rect 12173 7497 12207 7531
rect 12207 7497 12216 7531
rect 12164 7488 12216 7497
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 11428 7420 11480 7472
rect 12256 7420 12308 7472
rect 11980 7352 12032 7404
rect 12808 7352 12860 7404
rect 11796 7284 11848 7336
rect 9128 7216 9180 7268
rect 9864 7216 9916 7268
rect 11152 7216 11204 7268
rect 12348 7216 12400 7268
rect 12900 7284 12952 7336
rect 14004 7488 14056 7540
rect 15016 7488 15068 7540
rect 17684 7488 17736 7540
rect 19340 7531 19392 7540
rect 19340 7497 19349 7531
rect 19349 7497 19383 7531
rect 19383 7497 19392 7531
rect 19340 7488 19392 7497
rect 19708 7488 19760 7540
rect 20352 7531 20404 7540
rect 20352 7497 20361 7531
rect 20361 7497 20395 7531
rect 20395 7497 20404 7531
rect 20352 7488 20404 7497
rect 20812 7488 20864 7540
rect 14740 7420 14792 7472
rect 16396 7420 16448 7472
rect 19524 7420 19576 7472
rect 20628 7420 20680 7472
rect 20996 7420 21048 7472
rect 14280 7352 14332 7404
rect 15016 7352 15068 7404
rect 15384 7395 15436 7404
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 17224 7352 17276 7404
rect 17408 7395 17460 7404
rect 17408 7361 17442 7395
rect 17442 7361 17460 7395
rect 17408 7352 17460 7361
rect 18972 7395 19024 7404
rect 18972 7361 18981 7395
rect 18981 7361 19015 7395
rect 19015 7361 19024 7395
rect 18972 7352 19024 7361
rect 20352 7352 20404 7404
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 13452 7284 13504 7336
rect 9404 7191 9456 7200
rect 9404 7157 9413 7191
rect 9413 7157 9447 7191
rect 9447 7157 9456 7191
rect 9404 7148 9456 7157
rect 10140 7148 10192 7200
rect 11428 7148 11480 7200
rect 11704 7191 11756 7200
rect 11704 7157 11713 7191
rect 11713 7157 11747 7191
rect 11747 7157 11756 7191
rect 11704 7148 11756 7157
rect 13084 7148 13136 7200
rect 13360 7191 13412 7200
rect 13360 7157 13369 7191
rect 13369 7157 13403 7191
rect 13403 7157 13412 7191
rect 13360 7148 13412 7157
rect 13728 7148 13780 7200
rect 14280 7148 14332 7200
rect 15292 7284 15344 7336
rect 16028 7284 16080 7336
rect 16672 7284 16724 7336
rect 17040 7284 17092 7336
rect 18880 7327 18932 7336
rect 16304 7216 16356 7268
rect 18512 7259 18564 7268
rect 18512 7225 18521 7259
rect 18521 7225 18555 7259
rect 18555 7225 18564 7259
rect 18880 7293 18889 7327
rect 18889 7293 18923 7327
rect 18923 7293 18932 7327
rect 18880 7284 18932 7293
rect 19892 7327 19944 7336
rect 19892 7293 19901 7327
rect 19901 7293 19935 7327
rect 19935 7293 19944 7327
rect 19892 7284 19944 7293
rect 18512 7216 18564 7225
rect 20260 7216 20312 7268
rect 15752 7191 15804 7200
rect 15752 7157 15761 7191
rect 15761 7157 15795 7191
rect 15795 7157 15804 7191
rect 15752 7148 15804 7157
rect 16488 7148 16540 7200
rect 17132 7148 17184 7200
rect 21088 7148 21140 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 2044 6944 2096 6996
rect 3056 6944 3108 6996
rect 6828 6944 6880 6996
rect 6920 6944 6972 6996
rect 7656 6944 7708 6996
rect 9588 6944 9640 6996
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 2780 6876 2832 6928
rect 3240 6919 3292 6928
rect 3240 6885 3249 6919
rect 3249 6885 3283 6919
rect 3283 6885 3292 6919
rect 3240 6876 3292 6885
rect 3976 6876 4028 6928
rect 3700 6808 3752 6860
rect 5264 6808 5316 6860
rect 6552 6876 6604 6928
rect 7196 6876 7248 6928
rect 9864 6944 9916 6996
rect 5816 6808 5868 6860
rect 112 6740 164 6792
rect 940 6740 992 6792
rect 1216 6740 1268 6792
rect 1860 6672 1912 6724
rect 2780 6740 2832 6792
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 4344 6740 4396 6792
rect 2044 6715 2096 6724
rect 2044 6681 2053 6715
rect 2053 6681 2087 6715
rect 2087 6681 2096 6715
rect 2044 6672 2096 6681
rect 3516 6672 3568 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 2780 6604 2832 6613
rect 3240 6604 3292 6656
rect 3332 6604 3384 6656
rect 5724 6740 5776 6792
rect 7196 6740 7248 6792
rect 7472 6740 7524 6792
rect 9036 6808 9088 6860
rect 11152 6944 11204 6996
rect 11796 6987 11848 6996
rect 11796 6953 11805 6987
rect 11805 6953 11839 6987
rect 11839 6953 11848 6987
rect 11796 6944 11848 6953
rect 12256 6944 12308 6996
rect 12532 6876 12584 6928
rect 11152 6808 11204 6860
rect 11888 6808 11940 6860
rect 12348 6851 12400 6860
rect 12348 6817 12357 6851
rect 12357 6817 12391 6851
rect 12391 6817 12400 6851
rect 12348 6808 12400 6817
rect 14740 6876 14792 6928
rect 15384 6944 15436 6996
rect 16396 6944 16448 6996
rect 17132 6944 17184 6996
rect 17500 6944 17552 6996
rect 9220 6740 9272 6792
rect 9312 6740 9364 6792
rect 9680 6740 9732 6792
rect 5264 6672 5316 6724
rect 4160 6604 4212 6656
rect 4344 6647 4396 6656
rect 4344 6613 4353 6647
rect 4353 6613 4387 6647
rect 4387 6613 4396 6647
rect 4344 6604 4396 6613
rect 4712 6604 4764 6656
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 6000 6647 6052 6656
rect 6000 6613 6009 6647
rect 6009 6613 6043 6647
rect 6043 6613 6052 6647
rect 6644 6672 6696 6724
rect 8024 6672 8076 6724
rect 10416 6672 10468 6724
rect 10784 6740 10836 6792
rect 12164 6783 12216 6792
rect 12164 6749 12173 6783
rect 12173 6749 12207 6783
rect 12207 6749 12216 6783
rect 12164 6740 12216 6749
rect 13636 6808 13688 6860
rect 14188 6851 14240 6860
rect 14188 6817 14197 6851
rect 14197 6817 14231 6851
rect 14231 6817 14240 6851
rect 14188 6808 14240 6817
rect 16028 6876 16080 6928
rect 12900 6740 12952 6792
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 15200 6851 15252 6860
rect 15200 6817 15209 6851
rect 15209 6817 15243 6851
rect 15243 6817 15252 6851
rect 15200 6808 15252 6817
rect 15384 6808 15436 6860
rect 15568 6808 15620 6860
rect 18144 6808 18196 6860
rect 18512 6876 18564 6928
rect 18880 6944 18932 6996
rect 21272 6944 21324 6996
rect 20996 6851 21048 6860
rect 20996 6817 21005 6851
rect 21005 6817 21039 6851
rect 21039 6817 21048 6851
rect 20996 6808 21048 6817
rect 16212 6740 16264 6792
rect 16672 6740 16724 6792
rect 17224 6740 17276 6792
rect 17500 6740 17552 6792
rect 6000 6604 6052 6613
rect 6736 6647 6788 6656
rect 6736 6613 6745 6647
rect 6745 6613 6779 6647
rect 6779 6613 6788 6647
rect 6736 6604 6788 6613
rect 7380 6604 7432 6656
rect 8208 6604 8260 6656
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 8944 6604 8996 6656
rect 9312 6604 9364 6656
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 10232 6604 10284 6656
rect 11244 6604 11296 6656
rect 11704 6604 11756 6656
rect 11796 6604 11848 6656
rect 14556 6672 14608 6724
rect 15568 6672 15620 6724
rect 17684 6672 17736 6724
rect 18788 6740 18840 6792
rect 13820 6647 13872 6656
rect 13820 6613 13829 6647
rect 13829 6613 13863 6647
rect 13863 6613 13872 6647
rect 13820 6604 13872 6613
rect 14832 6647 14884 6656
rect 14832 6613 14841 6647
rect 14841 6613 14875 6647
rect 14875 6613 14884 6647
rect 14832 6604 14884 6613
rect 15936 6647 15988 6656
rect 15936 6613 15945 6647
rect 15945 6613 15979 6647
rect 15979 6613 15988 6647
rect 15936 6604 15988 6613
rect 16948 6604 17000 6656
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 17868 6647 17920 6656
rect 17868 6613 17877 6647
rect 17877 6613 17911 6647
rect 17911 6613 17920 6647
rect 19064 6740 19116 6792
rect 19156 6672 19208 6724
rect 20260 6740 20312 6792
rect 22100 6740 22152 6792
rect 19432 6672 19484 6724
rect 19800 6672 19852 6724
rect 22468 6672 22520 6724
rect 17868 6604 17920 6613
rect 20260 6604 20312 6656
rect 20444 6604 20496 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 2596 6332 2648 6384
rect 2964 6332 3016 6384
rect 3240 6400 3292 6452
rect 3700 6332 3752 6384
rect 4068 6332 4120 6384
rect 4988 6332 5040 6384
rect 6460 6400 6512 6452
rect 6552 6400 6604 6452
rect 6276 6332 6328 6384
rect 2872 6264 2924 6316
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 3240 6196 3292 6248
rect 4160 6264 4212 6316
rect 6092 6264 6144 6316
rect 6184 6307 6236 6316
rect 6184 6273 6193 6307
rect 6193 6273 6227 6307
rect 6227 6273 6236 6307
rect 7012 6332 7064 6384
rect 7380 6400 7432 6452
rect 7656 6443 7708 6452
rect 7656 6409 7665 6443
rect 7665 6409 7699 6443
rect 7699 6409 7708 6443
rect 7656 6400 7708 6409
rect 7748 6400 7800 6452
rect 8392 6443 8444 6452
rect 7564 6375 7616 6384
rect 7564 6341 7573 6375
rect 7573 6341 7607 6375
rect 7607 6341 7616 6375
rect 7564 6332 7616 6341
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 8668 6400 8720 6452
rect 10968 6443 11020 6452
rect 10968 6409 10977 6443
rect 10977 6409 11011 6443
rect 11011 6409 11020 6443
rect 10968 6400 11020 6409
rect 11060 6443 11112 6452
rect 11060 6409 11069 6443
rect 11069 6409 11103 6443
rect 11103 6409 11112 6443
rect 11060 6400 11112 6409
rect 6184 6264 6236 6273
rect 4712 6196 4764 6248
rect 5632 6196 5684 6248
rect 5264 6128 5316 6180
rect 6828 6196 6880 6248
rect 7564 6196 7616 6248
rect 7840 6196 7892 6248
rect 8668 6264 8720 6316
rect 8944 6264 8996 6316
rect 9496 6264 9548 6316
rect 12624 6400 12676 6452
rect 13268 6443 13320 6452
rect 13268 6409 13277 6443
rect 13277 6409 13311 6443
rect 13311 6409 13320 6443
rect 13268 6400 13320 6409
rect 13360 6400 13412 6452
rect 13820 6332 13872 6384
rect 14188 6332 14240 6384
rect 12716 6264 12768 6316
rect 13360 6264 13412 6316
rect 13912 6264 13964 6316
rect 15752 6400 15804 6452
rect 16948 6443 17000 6452
rect 16948 6409 16957 6443
rect 16957 6409 16991 6443
rect 16991 6409 17000 6443
rect 16948 6400 17000 6409
rect 18512 6400 18564 6452
rect 18972 6443 19024 6452
rect 18972 6409 18981 6443
rect 18981 6409 19015 6443
rect 19015 6409 19024 6443
rect 18972 6400 19024 6409
rect 19524 6400 19576 6452
rect 20260 6443 20312 6452
rect 14832 6332 14884 6384
rect 16120 6332 16172 6384
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 11152 6239 11204 6248
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 2320 6060 2372 6112
rect 3148 6060 3200 6112
rect 4988 6060 5040 6112
rect 5080 6060 5132 6112
rect 6552 6060 6604 6112
rect 7472 6060 7524 6112
rect 8760 6128 8812 6180
rect 9312 6128 9364 6180
rect 10140 6128 10192 6180
rect 11152 6205 11161 6239
rect 11161 6205 11195 6239
rect 11195 6205 11204 6239
rect 11152 6196 11204 6205
rect 12440 6196 12492 6248
rect 7840 6060 7892 6112
rect 8300 6060 8352 6112
rect 10600 6060 10652 6112
rect 10784 6060 10836 6112
rect 12624 6060 12676 6112
rect 12900 6060 12952 6112
rect 13360 6103 13412 6112
rect 13360 6069 13369 6103
rect 13369 6069 13403 6103
rect 13403 6069 13412 6103
rect 13360 6060 13412 6069
rect 16396 6264 16448 6316
rect 17224 6264 17276 6316
rect 17684 6264 17736 6316
rect 18052 6264 18104 6316
rect 16488 6239 16540 6248
rect 15200 6171 15252 6180
rect 15200 6137 15209 6171
rect 15209 6137 15243 6171
rect 15243 6137 15252 6171
rect 16488 6205 16497 6239
rect 16497 6205 16531 6239
rect 16531 6205 16540 6239
rect 16488 6196 16540 6205
rect 17316 6196 17368 6248
rect 17500 6196 17552 6248
rect 18144 6239 18196 6248
rect 18144 6205 18153 6239
rect 18153 6205 18187 6239
rect 18187 6205 18196 6239
rect 18144 6196 18196 6205
rect 19064 6332 19116 6384
rect 20260 6409 20269 6443
rect 20269 6409 20303 6443
rect 20303 6409 20312 6443
rect 20260 6400 20312 6409
rect 21180 6400 21232 6452
rect 18788 6307 18840 6316
rect 18788 6273 18797 6307
rect 18797 6273 18831 6307
rect 18831 6273 18840 6307
rect 18788 6264 18840 6273
rect 20812 6332 20864 6384
rect 19340 6264 19392 6316
rect 19432 6239 19484 6248
rect 15200 6128 15252 6137
rect 16212 6128 16264 6180
rect 19432 6205 19441 6239
rect 19441 6205 19475 6239
rect 19475 6205 19484 6239
rect 19432 6196 19484 6205
rect 20444 6264 20496 6316
rect 20536 6196 20588 6248
rect 20720 6239 20772 6248
rect 20720 6205 20729 6239
rect 20729 6205 20763 6239
rect 20763 6205 20772 6239
rect 20720 6196 20772 6205
rect 19064 6128 19116 6180
rect 19892 6128 19944 6180
rect 20168 6128 20220 6180
rect 16028 6103 16080 6112
rect 16028 6069 16037 6103
rect 16037 6069 16071 6103
rect 16071 6069 16080 6103
rect 16028 6060 16080 6069
rect 16120 6060 16172 6112
rect 17316 6060 17368 6112
rect 17684 6060 17736 6112
rect 18328 6103 18380 6112
rect 18328 6069 18337 6103
rect 18337 6069 18371 6103
rect 18371 6069 18380 6103
rect 18328 6060 18380 6069
rect 18604 6060 18656 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 1492 5856 1544 5908
rect 940 5788 992 5840
rect 1400 5720 1452 5772
rect 1676 5720 1728 5772
rect 2596 5720 2648 5772
rect 3148 5788 3200 5840
rect 3332 5788 3384 5840
rect 3516 5856 3568 5908
rect 5816 5899 5868 5908
rect 5816 5865 5825 5899
rect 5825 5865 5859 5899
rect 5859 5865 5868 5899
rect 5816 5856 5868 5865
rect 5908 5856 5960 5908
rect 6460 5856 6512 5908
rect 10048 5856 10100 5908
rect 6000 5788 6052 5840
rect 4436 5763 4488 5772
rect 3148 5652 3200 5704
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 5632 5720 5684 5772
rect 7840 5788 7892 5840
rect 10416 5856 10468 5908
rect 10968 5856 11020 5908
rect 11060 5856 11112 5908
rect 11336 5856 11388 5908
rect 12440 5856 12492 5908
rect 12624 5856 12676 5908
rect 4712 5695 4764 5704
rect 2228 5584 2280 5636
rect 3056 5584 3108 5636
rect 2136 5516 2188 5568
rect 2780 5559 2832 5568
rect 2780 5525 2789 5559
rect 2789 5525 2823 5559
rect 2823 5525 2832 5559
rect 4252 5584 4304 5636
rect 4712 5661 4746 5695
rect 4746 5661 4764 5695
rect 4712 5652 4764 5661
rect 5724 5652 5776 5704
rect 4988 5584 5040 5636
rect 2780 5516 2832 5525
rect 3792 5516 3844 5568
rect 6460 5652 6512 5704
rect 7196 5652 7248 5704
rect 6920 5584 6972 5636
rect 8116 5584 8168 5636
rect 6276 5559 6328 5568
rect 6276 5525 6285 5559
rect 6285 5525 6319 5559
rect 6319 5525 6328 5559
rect 6276 5516 6328 5525
rect 6368 5516 6420 5568
rect 7012 5516 7064 5568
rect 7840 5516 7892 5568
rect 8208 5516 8260 5568
rect 8944 5763 8996 5772
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 8484 5652 8536 5661
rect 8944 5729 8953 5763
rect 8953 5729 8987 5763
rect 8987 5729 8996 5763
rect 8944 5720 8996 5729
rect 10784 5720 10836 5772
rect 9036 5652 9088 5704
rect 10140 5652 10192 5704
rect 11796 5788 11848 5840
rect 11152 5720 11204 5772
rect 14280 5788 14332 5840
rect 15568 5831 15620 5840
rect 15568 5797 15577 5831
rect 15577 5797 15611 5831
rect 15611 5797 15620 5831
rect 15568 5788 15620 5797
rect 13728 5720 13780 5772
rect 9588 5584 9640 5636
rect 9864 5584 9916 5636
rect 12256 5652 12308 5704
rect 13820 5652 13872 5704
rect 14372 5652 14424 5704
rect 15200 5695 15252 5704
rect 15200 5661 15218 5695
rect 15218 5661 15252 5695
rect 15200 5652 15252 5661
rect 10784 5584 10836 5636
rect 16580 5856 16632 5908
rect 17684 5856 17736 5908
rect 18144 5788 18196 5840
rect 18328 5788 18380 5840
rect 18972 5856 19024 5908
rect 21088 5856 21140 5908
rect 19064 5788 19116 5840
rect 20812 5788 20864 5840
rect 15752 5652 15804 5704
rect 16120 5720 16172 5772
rect 16488 5720 16540 5772
rect 17132 5720 17184 5772
rect 17776 5720 17828 5772
rect 17960 5720 18012 5772
rect 17684 5652 17736 5704
rect 18052 5652 18104 5704
rect 18328 5652 18380 5704
rect 18880 5652 18932 5704
rect 20812 5652 20864 5704
rect 20996 5652 21048 5704
rect 16304 5584 16356 5636
rect 17500 5584 17552 5636
rect 11060 5559 11112 5568
rect 11060 5525 11069 5559
rect 11069 5525 11103 5559
rect 11103 5525 11112 5559
rect 11520 5559 11572 5568
rect 11060 5516 11112 5525
rect 11520 5525 11529 5559
rect 11529 5525 11563 5559
rect 11563 5525 11572 5559
rect 11520 5516 11572 5525
rect 11796 5516 11848 5568
rect 12624 5559 12676 5568
rect 12624 5525 12633 5559
rect 12633 5525 12667 5559
rect 12667 5525 12676 5559
rect 12624 5516 12676 5525
rect 13636 5516 13688 5568
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 15568 5516 15620 5568
rect 16580 5559 16632 5568
rect 16580 5525 16589 5559
rect 16589 5525 16623 5559
rect 16623 5525 16632 5559
rect 16948 5559 17000 5568
rect 16580 5516 16632 5525
rect 16948 5525 16957 5559
rect 16957 5525 16991 5559
rect 16991 5525 17000 5559
rect 16948 5516 17000 5525
rect 17316 5516 17368 5568
rect 18972 5627 19024 5636
rect 18972 5593 18981 5627
rect 18981 5593 19015 5627
rect 19015 5593 19024 5627
rect 18972 5584 19024 5593
rect 19708 5584 19760 5636
rect 22928 5584 22980 5636
rect 18052 5559 18104 5568
rect 18052 5525 18061 5559
rect 18061 5525 18095 5559
rect 18095 5525 18104 5559
rect 18052 5516 18104 5525
rect 18236 5516 18288 5568
rect 18512 5559 18564 5568
rect 18512 5525 18521 5559
rect 18521 5525 18555 5559
rect 18555 5525 18564 5559
rect 18512 5516 18564 5525
rect 20720 5559 20772 5568
rect 20720 5525 20729 5559
rect 20729 5525 20763 5559
rect 20763 5525 20772 5559
rect 21088 5559 21140 5568
rect 20720 5516 20772 5525
rect 21088 5525 21097 5559
rect 21097 5525 21131 5559
rect 21131 5525 21140 5559
rect 21088 5516 21140 5525
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 3056 5312 3108 5364
rect 5264 5312 5316 5364
rect 5724 5312 5776 5364
rect 5816 5312 5868 5364
rect 1584 5244 1636 5296
rect 3424 5244 3476 5296
rect 3884 5244 3936 5296
rect 4252 5244 4304 5296
rect 4988 5244 5040 5296
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 2596 5176 2648 5228
rect 5080 5176 5132 5228
rect 7012 5312 7064 5364
rect 7564 5355 7616 5364
rect 7564 5321 7573 5355
rect 7573 5321 7607 5355
rect 7607 5321 7616 5355
rect 7564 5312 7616 5321
rect 8208 5355 8260 5364
rect 8208 5321 8217 5355
rect 8217 5321 8251 5355
rect 8251 5321 8260 5355
rect 8208 5312 8260 5321
rect 8300 5355 8352 5364
rect 8300 5321 8309 5355
rect 8309 5321 8343 5355
rect 8343 5321 8352 5355
rect 8300 5312 8352 5321
rect 9772 5312 9824 5364
rect 10140 5355 10192 5364
rect 10140 5321 10149 5355
rect 10149 5321 10183 5355
rect 10183 5321 10192 5355
rect 10140 5312 10192 5321
rect 10508 5312 10560 5364
rect 11060 5312 11112 5364
rect 11336 5355 11388 5364
rect 11336 5321 11345 5355
rect 11345 5321 11379 5355
rect 11379 5321 11388 5355
rect 11336 5312 11388 5321
rect 12164 5312 12216 5364
rect 12348 5312 12400 5364
rect 12624 5312 12676 5364
rect 12716 5312 12768 5364
rect 2228 5151 2280 5160
rect 2228 5117 2237 5151
rect 2237 5117 2271 5151
rect 2271 5117 2280 5151
rect 2228 5108 2280 5117
rect 1032 4972 1084 5024
rect 3884 5108 3936 5160
rect 4712 5040 4764 5092
rect 6092 5176 6144 5228
rect 6276 5176 6328 5228
rect 7288 5244 7340 5296
rect 5632 5108 5684 5160
rect 6460 5108 6512 5160
rect 7564 5176 7616 5228
rect 7748 5176 7800 5228
rect 8024 5244 8076 5296
rect 8484 5176 8536 5228
rect 8668 5176 8720 5228
rect 9036 5219 9088 5228
rect 9036 5185 9070 5219
rect 9070 5185 9088 5219
rect 9036 5176 9088 5185
rect 9312 5176 9364 5228
rect 9496 5176 9548 5228
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 11796 5176 11848 5228
rect 12900 5176 12952 5228
rect 13820 5176 13872 5228
rect 14372 5219 14424 5228
rect 14372 5185 14381 5219
rect 14381 5185 14415 5219
rect 14415 5185 14424 5219
rect 14372 5176 14424 5185
rect 14924 5312 14976 5364
rect 15016 5355 15068 5364
rect 15016 5321 15025 5355
rect 15025 5321 15059 5355
rect 15059 5321 15068 5355
rect 15200 5355 15252 5364
rect 15016 5312 15068 5321
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 15660 5312 15712 5364
rect 17592 5312 17644 5364
rect 15844 5244 15896 5296
rect 16396 5244 16448 5296
rect 16580 5244 16632 5296
rect 17132 5244 17184 5296
rect 10784 5151 10836 5160
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 7288 5040 7340 5092
rect 8760 5040 8812 5092
rect 10692 5040 10744 5092
rect 11612 5108 11664 5160
rect 11060 5040 11112 5092
rect 12256 5040 12308 5092
rect 3240 4972 3292 5024
rect 4160 4972 4212 5024
rect 4620 4972 4672 5024
rect 5632 4972 5684 5024
rect 6184 4972 6236 5024
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 7656 5015 7708 5024
rect 7656 4981 7665 5015
rect 7665 4981 7699 5015
rect 7699 4981 7708 5015
rect 7656 4972 7708 4981
rect 7840 4972 7892 5024
rect 10140 4972 10192 5024
rect 11428 4972 11480 5024
rect 11612 4972 11664 5024
rect 12716 4972 12768 5024
rect 14464 5108 14516 5160
rect 15844 5108 15896 5160
rect 16764 5108 16816 5160
rect 16948 5108 17000 5160
rect 17960 5244 18012 5296
rect 20720 5312 20772 5364
rect 17868 5219 17920 5228
rect 17868 5185 17877 5219
rect 17877 5185 17911 5219
rect 17911 5185 17920 5219
rect 17868 5176 17920 5185
rect 18420 5176 18472 5228
rect 21548 5219 21600 5228
rect 21548 5185 21557 5219
rect 21557 5185 21591 5219
rect 21591 5185 21600 5219
rect 21548 5176 21600 5185
rect 18328 5151 18380 5160
rect 13268 5040 13320 5092
rect 14372 5040 14424 5092
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 12992 4972 13044 4981
rect 15016 4972 15068 5024
rect 16396 4972 16448 5024
rect 16580 4972 16632 5024
rect 16856 4972 16908 5024
rect 18328 5117 18337 5151
rect 18337 5117 18371 5151
rect 18371 5117 18380 5151
rect 18328 5108 18380 5117
rect 20444 5151 20496 5160
rect 20444 5117 20453 5151
rect 20453 5117 20487 5151
rect 20487 5117 20496 5151
rect 20444 5108 20496 5117
rect 22100 5108 22152 5160
rect 20352 5040 20404 5092
rect 19524 4972 19576 5024
rect 19708 5015 19760 5024
rect 19708 4981 19717 5015
rect 19717 4981 19751 5015
rect 19751 4981 19760 5015
rect 19708 4972 19760 4981
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 2596 4768 2648 4820
rect 3332 4768 3384 4820
rect 4436 4768 4488 4820
rect 4896 4768 4948 4820
rect 5264 4768 5316 4820
rect 2044 4700 2096 4752
rect 1124 4564 1176 4616
rect 1952 4564 2004 4616
rect 3884 4632 3936 4684
rect 3056 4539 3108 4548
rect 3056 4505 3074 4539
rect 3074 4505 3108 4539
rect 3608 4607 3660 4616
rect 3608 4573 3617 4607
rect 3617 4573 3651 4607
rect 3651 4573 3660 4607
rect 3608 4564 3660 4573
rect 3792 4564 3844 4616
rect 4436 4607 4488 4616
rect 4436 4573 4445 4607
rect 4445 4573 4479 4607
rect 4479 4573 4488 4607
rect 4436 4564 4488 4573
rect 5080 4632 5132 4684
rect 5724 4700 5776 4752
rect 6276 4700 6328 4752
rect 6828 4768 6880 4820
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 5908 4675 5960 4684
rect 5908 4641 5917 4675
rect 5917 4641 5951 4675
rect 5951 4641 5960 4675
rect 5908 4632 5960 4641
rect 6184 4632 6236 4684
rect 6460 4632 6512 4684
rect 8300 4768 8352 4820
rect 9220 4768 9272 4820
rect 11704 4811 11756 4820
rect 11704 4777 11713 4811
rect 11713 4777 11747 4811
rect 11747 4777 11756 4811
rect 11704 4768 11756 4777
rect 12900 4811 12952 4820
rect 12900 4777 12909 4811
rect 12909 4777 12943 4811
rect 12943 4777 12952 4811
rect 12900 4768 12952 4777
rect 13084 4768 13136 4820
rect 15292 4768 15344 4820
rect 16764 4811 16816 4820
rect 16764 4777 16773 4811
rect 16773 4777 16807 4811
rect 16807 4777 16816 4811
rect 16764 4768 16816 4777
rect 17868 4768 17920 4820
rect 21640 4768 21692 4820
rect 8576 4700 8628 4752
rect 9312 4700 9364 4752
rect 8116 4675 8168 4684
rect 8116 4641 8125 4675
rect 8125 4641 8159 4675
rect 8159 4641 8168 4675
rect 8116 4632 8168 4641
rect 9128 4632 9180 4684
rect 10784 4700 10836 4752
rect 10968 4700 11020 4752
rect 12624 4700 12676 4752
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 10416 4675 10468 4684
rect 10416 4641 10425 4675
rect 10425 4641 10459 4675
rect 10459 4641 10468 4675
rect 10416 4632 10468 4641
rect 11244 4632 11296 4684
rect 13820 4700 13872 4752
rect 14740 4700 14792 4752
rect 13728 4632 13780 4684
rect 14372 4632 14424 4684
rect 18420 4700 18472 4752
rect 5448 4564 5500 4616
rect 6092 4564 6144 4616
rect 3056 4496 3108 4505
rect 4160 4496 4212 4548
rect 4620 4496 4672 4548
rect 2044 4428 2096 4480
rect 3608 4428 3660 4480
rect 3976 4471 4028 4480
rect 3976 4437 3985 4471
rect 3985 4437 4019 4471
rect 4019 4437 4028 4471
rect 3976 4428 4028 4437
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 4804 4471 4856 4480
rect 4804 4437 4813 4471
rect 4813 4437 4847 4471
rect 4847 4437 4856 4471
rect 4804 4428 4856 4437
rect 4896 4471 4948 4480
rect 4896 4437 4905 4471
rect 4905 4437 4939 4471
rect 4939 4437 4948 4471
rect 5816 4496 5868 4548
rect 7748 4564 7800 4616
rect 8576 4564 8628 4616
rect 4896 4428 4948 4437
rect 5448 4428 5500 4480
rect 7288 4496 7340 4548
rect 9772 4564 9824 4616
rect 10600 4607 10652 4616
rect 10600 4573 10609 4607
rect 10609 4573 10643 4607
rect 10643 4573 10652 4607
rect 10600 4564 10652 4573
rect 11428 4564 11480 4616
rect 12256 4564 12308 4616
rect 7012 4428 7064 4480
rect 8024 4471 8076 4480
rect 8024 4437 8033 4471
rect 8033 4437 8067 4471
rect 8067 4437 8076 4471
rect 9956 4496 10008 4548
rect 10232 4496 10284 4548
rect 8024 4428 8076 4437
rect 9220 4428 9272 4480
rect 10784 4471 10836 4480
rect 10784 4437 10793 4471
rect 10793 4437 10827 4471
rect 10827 4437 10836 4471
rect 10784 4428 10836 4437
rect 11336 4539 11388 4548
rect 11336 4505 11345 4539
rect 11345 4505 11379 4539
rect 11379 4505 11388 4539
rect 11336 4496 11388 4505
rect 12348 4496 12400 4548
rect 12532 4539 12584 4548
rect 12532 4505 12541 4539
rect 12541 4505 12575 4539
rect 12575 4505 12584 4539
rect 12532 4496 12584 4505
rect 13176 4496 13228 4548
rect 14464 4496 14516 4548
rect 14924 4496 14976 4548
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 19708 4632 19760 4684
rect 17960 4564 18012 4616
rect 18328 4564 18380 4616
rect 18696 4564 18748 4616
rect 19524 4607 19576 4616
rect 19524 4573 19533 4607
rect 19533 4573 19567 4607
rect 19567 4573 19576 4607
rect 19524 4564 19576 4573
rect 22560 4632 22612 4684
rect 15660 4539 15712 4548
rect 15660 4505 15694 4539
rect 15694 4505 15712 4539
rect 15660 4496 15712 4505
rect 18512 4496 18564 4548
rect 11888 4428 11940 4480
rect 12256 4428 12308 4480
rect 12624 4428 12676 4480
rect 13084 4428 13136 4480
rect 13360 4471 13412 4480
rect 13360 4437 13369 4471
rect 13369 4437 13403 4471
rect 13403 4437 13412 4471
rect 13360 4428 13412 4437
rect 14372 4471 14424 4480
rect 14372 4437 14381 4471
rect 14381 4437 14415 4471
rect 14415 4437 14424 4471
rect 14372 4428 14424 4437
rect 16948 4428 17000 4480
rect 18696 4471 18748 4480
rect 18696 4437 18705 4471
rect 18705 4437 18739 4471
rect 18739 4437 18748 4471
rect 18696 4428 18748 4437
rect 18788 4471 18840 4480
rect 18788 4437 18797 4471
rect 18797 4437 18831 4471
rect 18831 4437 18840 4471
rect 21364 4564 21416 4616
rect 18788 4428 18840 4437
rect 20720 4428 20772 4480
rect 21272 4428 21324 4480
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 1860 4267 1912 4276
rect 1860 4233 1869 4267
rect 1869 4233 1903 4267
rect 1903 4233 1912 4267
rect 1860 4224 1912 4233
rect 2780 4224 2832 4276
rect 3056 4224 3108 4276
rect 3884 4224 3936 4276
rect 4712 4224 4764 4276
rect 5540 4224 5592 4276
rect 3148 4156 3200 4208
rect 5908 4224 5960 4276
rect 8300 4224 8352 4276
rect 9496 4267 9548 4276
rect 9496 4233 9505 4267
rect 9505 4233 9539 4267
rect 9539 4233 9548 4267
rect 9496 4224 9548 4233
rect 11704 4224 11756 4276
rect 11796 4224 11848 4276
rect 12164 4224 12216 4276
rect 12624 4224 12676 4276
rect 12992 4224 13044 4276
rect 13728 4224 13780 4276
rect 16304 4224 16356 4276
rect 16856 4267 16908 4276
rect 16856 4233 16865 4267
rect 16865 4233 16899 4267
rect 16899 4233 16908 4267
rect 16856 4224 16908 4233
rect 16948 4224 17000 4276
rect 6276 4156 6328 4208
rect 6460 4156 6512 4208
rect 7104 4156 7156 4208
rect 1676 4063 1728 4072
rect 1676 4029 1685 4063
rect 1685 4029 1719 4063
rect 1719 4029 1728 4063
rect 1676 4020 1728 4029
rect 4896 4088 4948 4140
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 5540 4088 5592 4140
rect 2964 4020 3016 4072
rect 4620 4063 4672 4072
rect 4620 4029 4629 4063
rect 4629 4029 4663 4063
rect 4663 4029 4672 4063
rect 4620 4020 4672 4029
rect 4712 4063 4764 4072
rect 4712 4029 4721 4063
rect 4721 4029 4755 4063
rect 4755 4029 4764 4063
rect 4712 4020 4764 4029
rect 2872 3952 2924 4004
rect 3332 3952 3384 4004
rect 5448 4020 5500 4072
rect 6000 4020 6052 4072
rect 6184 4020 6236 4072
rect 6368 4063 6420 4072
rect 6368 4029 6377 4063
rect 6377 4029 6411 4063
rect 6411 4029 6420 4063
rect 6368 4020 6420 4029
rect 8116 4088 8168 4140
rect 8484 4131 8536 4140
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 9312 4088 9364 4140
rect 4804 3884 4856 3936
rect 5724 3884 5776 3936
rect 8116 3884 8168 3936
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 8760 3952 8812 4004
rect 9588 4020 9640 4072
rect 10784 4088 10836 4140
rect 9956 4063 10008 4072
rect 9956 4029 9965 4063
rect 9965 4029 9999 4063
rect 9999 4029 10008 4063
rect 9956 4020 10008 4029
rect 10968 4020 11020 4072
rect 12624 4131 12676 4140
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 13544 4156 13596 4208
rect 16120 4156 16172 4208
rect 12808 4088 12860 4140
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 13820 4088 13872 4140
rect 9680 3884 9732 3936
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 12532 3952 12584 4004
rect 13452 3952 13504 4004
rect 14924 4063 14976 4072
rect 13728 3952 13780 4004
rect 14924 4029 14933 4063
rect 14933 4029 14967 4063
rect 14967 4029 14976 4063
rect 14924 4020 14976 4029
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 15568 4020 15620 4072
rect 15936 4063 15988 4072
rect 15936 4029 15945 4063
rect 15945 4029 15979 4063
rect 15979 4029 15988 4063
rect 16396 4088 16448 4140
rect 16948 4088 17000 4140
rect 17224 4088 17276 4140
rect 15936 4020 15988 4029
rect 15660 3952 15712 4004
rect 16948 3952 17000 4004
rect 17592 4224 17644 4276
rect 18144 4224 18196 4276
rect 20444 4224 20496 4276
rect 17960 4020 18012 4072
rect 18972 4088 19024 4140
rect 19800 4131 19852 4140
rect 19800 4097 19809 4131
rect 19809 4097 19843 4131
rect 19843 4097 19852 4131
rect 19800 4088 19852 4097
rect 19984 4088 20036 4140
rect 20996 4156 21048 4208
rect 21088 4199 21140 4208
rect 21088 4165 21097 4199
rect 21097 4165 21131 4199
rect 21131 4165 21140 4199
rect 21456 4199 21508 4208
rect 21088 4156 21140 4165
rect 21456 4165 21465 4199
rect 21465 4165 21499 4199
rect 21499 4165 21508 4199
rect 21456 4156 21508 4165
rect 22008 4156 22060 4208
rect 22560 4156 22612 4208
rect 17776 3952 17828 4004
rect 18052 3952 18104 4004
rect 18236 3995 18288 4004
rect 18236 3961 18245 3995
rect 18245 3961 18279 3995
rect 18279 3961 18288 3995
rect 18236 3952 18288 3961
rect 12348 3927 12400 3936
rect 12348 3893 12357 3927
rect 12357 3893 12391 3927
rect 12391 3893 12400 3927
rect 12348 3884 12400 3893
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 12900 3884 12952 3936
rect 14556 3884 14608 3936
rect 14740 3884 14792 3936
rect 17224 3884 17276 3936
rect 19708 3952 19760 4004
rect 20168 3952 20220 4004
rect 20720 4088 20772 4140
rect 20536 4020 20588 4072
rect 22008 4020 22060 4072
rect 19432 3927 19484 3936
rect 19432 3893 19441 3927
rect 19441 3893 19475 3927
rect 19475 3893 19484 3927
rect 19432 3884 19484 3893
rect 20444 3884 20496 3936
rect 22192 3952 22244 4004
rect 21364 3927 21416 3936
rect 21364 3893 21373 3927
rect 21373 3893 21407 3927
rect 21407 3893 21416 3927
rect 21364 3884 21416 3893
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 2044 3680 2096 3732
rect 5540 3680 5592 3732
rect 5908 3680 5960 3732
rect 8300 3680 8352 3732
rect 8668 3680 8720 3732
rect 10140 3723 10192 3732
rect 10140 3689 10149 3723
rect 10149 3689 10183 3723
rect 10183 3689 10192 3723
rect 10140 3680 10192 3689
rect 1676 3655 1728 3664
rect 1676 3621 1685 3655
rect 1685 3621 1719 3655
rect 1719 3621 1728 3655
rect 1676 3612 1728 3621
rect 2320 3612 2372 3664
rect 1860 3544 1912 3596
rect 4712 3612 4764 3664
rect 2596 3587 2648 3596
rect 2596 3553 2605 3587
rect 2605 3553 2639 3587
rect 2639 3553 2648 3587
rect 2596 3544 2648 3553
rect 3056 3544 3108 3596
rect 3516 3544 3568 3596
rect 8116 3612 8168 3664
rect 1492 3519 1544 3528
rect 1492 3485 1501 3519
rect 1501 3485 1535 3519
rect 1535 3485 1544 3519
rect 1492 3476 1544 3485
rect 2504 3476 2556 3528
rect 4620 3476 4672 3528
rect 7012 3544 7064 3596
rect 9312 3612 9364 3664
rect 10048 3612 10100 3664
rect 10692 3680 10744 3732
rect 11244 3680 11296 3732
rect 11888 3723 11940 3732
rect 11888 3689 11897 3723
rect 11897 3689 11931 3723
rect 11931 3689 11940 3723
rect 11888 3680 11940 3689
rect 12348 3680 12400 3732
rect 13176 3680 13228 3732
rect 13268 3680 13320 3732
rect 14464 3680 14516 3732
rect 14924 3680 14976 3732
rect 13912 3612 13964 3664
rect 16856 3723 16908 3732
rect 16856 3689 16865 3723
rect 16865 3689 16899 3723
rect 16899 3689 16908 3723
rect 16856 3680 16908 3689
rect 18696 3680 18748 3732
rect 18788 3680 18840 3732
rect 19892 3680 19944 3732
rect 20168 3680 20220 3732
rect 20536 3680 20588 3732
rect 20720 3680 20772 3732
rect 22652 3680 22704 3732
rect 5080 3519 5132 3528
rect 5080 3485 5114 3519
rect 5114 3485 5132 3519
rect 3884 3408 3936 3460
rect 5080 3476 5132 3485
rect 5448 3476 5500 3528
rect 6552 3476 6604 3528
rect 6828 3476 6880 3528
rect 8392 3544 8444 3596
rect 8668 3544 8720 3596
rect 12532 3587 12584 3596
rect 8760 3476 8812 3528
rect 6000 3408 6052 3460
rect 6184 3408 6236 3460
rect 7012 3408 7064 3460
rect 3240 3383 3292 3392
rect 3240 3349 3249 3383
rect 3249 3349 3283 3383
rect 3283 3349 3292 3383
rect 3240 3340 3292 3349
rect 3332 3383 3384 3392
rect 3332 3349 3341 3383
rect 3341 3349 3375 3383
rect 3375 3349 3384 3383
rect 4344 3383 4396 3392
rect 3332 3340 3384 3349
rect 4344 3349 4353 3383
rect 4353 3349 4387 3383
rect 4387 3349 4396 3383
rect 4344 3340 4396 3349
rect 5448 3340 5500 3392
rect 5540 3340 5592 3392
rect 7288 3340 7340 3392
rect 7840 3340 7892 3392
rect 8300 3340 8352 3392
rect 9128 3476 9180 3528
rect 9312 3476 9364 3528
rect 9956 3476 10008 3528
rect 12532 3553 12541 3587
rect 12541 3553 12575 3587
rect 12575 3553 12584 3587
rect 12532 3544 12584 3553
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 15936 3612 15988 3664
rect 17132 3612 17184 3664
rect 12440 3476 12492 3528
rect 9496 3408 9548 3460
rect 9680 3408 9732 3460
rect 11244 3408 11296 3460
rect 12808 3451 12860 3460
rect 12808 3417 12842 3451
rect 12842 3417 12860 3451
rect 17224 3544 17276 3596
rect 18604 3612 18656 3664
rect 18880 3612 18932 3664
rect 20996 3612 21048 3664
rect 19248 3544 19300 3596
rect 15660 3476 15712 3528
rect 15844 3476 15896 3528
rect 16028 3476 16080 3528
rect 17040 3476 17092 3528
rect 17316 3476 17368 3528
rect 20904 3544 20956 3596
rect 9956 3340 10008 3392
rect 10968 3340 11020 3392
rect 12808 3408 12860 3417
rect 13360 3340 13412 3392
rect 13728 3340 13780 3392
rect 14280 3340 14332 3392
rect 14464 3383 14516 3392
rect 14464 3349 14473 3383
rect 14473 3349 14507 3383
rect 14507 3349 14516 3383
rect 14464 3340 14516 3349
rect 14924 3340 14976 3392
rect 16856 3408 16908 3460
rect 15936 3340 15988 3392
rect 16396 3383 16448 3392
rect 16396 3349 16405 3383
rect 16405 3349 16439 3383
rect 16439 3349 16448 3383
rect 16396 3340 16448 3349
rect 19156 3408 19208 3460
rect 19616 3476 19668 3528
rect 19892 3476 19944 3528
rect 20076 3476 20128 3528
rect 20628 3519 20680 3528
rect 20628 3485 20637 3519
rect 20637 3485 20671 3519
rect 20671 3485 20680 3519
rect 20628 3476 20680 3485
rect 20720 3519 20772 3528
rect 20720 3485 20729 3519
rect 20729 3485 20763 3519
rect 20763 3485 20772 3519
rect 20720 3476 20772 3485
rect 21088 3476 21140 3528
rect 20904 3408 20956 3460
rect 20168 3340 20220 3392
rect 21364 3340 21416 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 2412 3179 2464 3188
rect 2412 3145 2421 3179
rect 2421 3145 2455 3179
rect 2455 3145 2464 3179
rect 2412 3136 2464 3145
rect 2688 3179 2740 3188
rect 2688 3145 2697 3179
rect 2697 3145 2731 3179
rect 2731 3145 2740 3179
rect 2688 3136 2740 3145
rect 3148 3136 3200 3188
rect 3332 3136 3384 3188
rect 5724 3179 5776 3188
rect 5724 3145 5733 3179
rect 5733 3145 5767 3179
rect 5767 3145 5776 3179
rect 5724 3136 5776 3145
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 6828 3136 6880 3188
rect 7012 3136 7064 3188
rect 3424 3111 3476 3120
rect 3424 3077 3433 3111
rect 3433 3077 3467 3111
rect 3467 3077 3476 3111
rect 3424 3068 3476 3077
rect 2136 3000 2188 3052
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 2688 2932 2740 2984
rect 848 2864 900 2916
rect 3516 3000 3568 3052
rect 7196 3068 7248 3120
rect 7380 3068 7432 3120
rect 7932 3068 7984 3120
rect 8116 3068 8168 3120
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 4160 3043 4212 3052
rect 3884 3000 3936 3009
rect 4160 3009 4194 3043
rect 4194 3009 4212 3043
rect 4160 3000 4212 3009
rect 8208 3043 8260 3052
rect 4896 2932 4948 2984
rect 5908 2975 5960 2984
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 7748 2975 7800 2984
rect 7748 2941 7757 2975
rect 7757 2941 7791 2975
rect 7791 2941 7800 2975
rect 7748 2932 7800 2941
rect 3148 2796 3200 2848
rect 5816 2864 5868 2916
rect 5356 2796 5408 2848
rect 6000 2796 6052 2848
rect 8208 3009 8217 3043
rect 8217 3009 8251 3043
rect 8251 3009 8260 3043
rect 8208 3000 8260 3009
rect 8760 3136 8812 3188
rect 9772 3136 9824 3188
rect 10140 3179 10192 3188
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 9220 3068 9272 3120
rect 10876 3136 10928 3188
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 12072 3136 12124 3188
rect 12808 3136 12860 3188
rect 13452 3136 13504 3188
rect 10692 3000 10744 3052
rect 11152 3068 11204 3120
rect 12164 3068 12216 3120
rect 13728 3136 13780 3188
rect 13820 3136 13872 3188
rect 14372 3136 14424 3188
rect 13176 3000 13228 3052
rect 14648 3000 14700 3052
rect 9312 2932 9364 2984
rect 11980 2932 12032 2984
rect 13820 2975 13872 2984
rect 13820 2941 13829 2975
rect 13829 2941 13863 2975
rect 13863 2941 13872 2975
rect 13820 2932 13872 2941
rect 14372 2975 14424 2984
rect 14372 2941 14381 2975
rect 14381 2941 14415 2975
rect 14415 2941 14424 2975
rect 14372 2932 14424 2941
rect 15016 3136 15068 3188
rect 15292 3136 15344 3188
rect 14924 3043 14976 3052
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 15200 3068 15252 3120
rect 15292 3043 15344 3052
rect 15292 3009 15301 3043
rect 15301 3009 15335 3043
rect 15335 3009 15344 3043
rect 15292 3000 15344 3009
rect 16396 3136 16448 3188
rect 15936 3068 15988 3120
rect 16212 3043 16264 3052
rect 16212 3009 16221 3043
rect 16221 3009 16255 3043
rect 16255 3009 16264 3043
rect 16212 3000 16264 3009
rect 16488 3000 16540 3052
rect 17040 3000 17092 3052
rect 18144 3136 18196 3188
rect 17592 3000 17644 3052
rect 18052 3000 18104 3052
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 19248 3136 19300 3188
rect 21088 3136 21140 3188
rect 19156 3000 19208 3052
rect 19616 3043 19668 3052
rect 19616 3009 19625 3043
rect 19625 3009 19659 3043
rect 19659 3009 19668 3043
rect 19616 3000 19668 3009
rect 20260 3043 20312 3052
rect 20260 3009 20269 3043
rect 20269 3009 20303 3043
rect 20303 3009 20312 3043
rect 20260 3000 20312 3009
rect 20352 3043 20404 3052
rect 20352 3009 20361 3043
rect 20361 3009 20395 3043
rect 20395 3009 20404 3043
rect 20352 3000 20404 3009
rect 21640 3000 21692 3052
rect 22744 3000 22796 3052
rect 8576 2796 8628 2848
rect 9588 2907 9640 2916
rect 9588 2873 9597 2907
rect 9597 2873 9631 2907
rect 9631 2873 9640 2907
rect 9588 2864 9640 2873
rect 11244 2864 11296 2916
rect 11152 2796 11204 2848
rect 11704 2796 11756 2848
rect 12164 2796 12216 2848
rect 13084 2796 13136 2848
rect 13452 2796 13504 2848
rect 17408 2932 17460 2984
rect 15568 2864 15620 2916
rect 16488 2864 16540 2916
rect 17316 2864 17368 2916
rect 18972 2932 19024 2984
rect 20812 2932 20864 2984
rect 18052 2864 18104 2916
rect 20628 2864 20680 2916
rect 14740 2839 14792 2848
rect 14740 2805 14749 2839
rect 14749 2805 14783 2839
rect 14783 2805 14792 2839
rect 14740 2796 14792 2805
rect 15200 2839 15252 2848
rect 15200 2805 15209 2839
rect 15209 2805 15243 2839
rect 15243 2805 15252 2839
rect 15200 2796 15252 2805
rect 15476 2796 15528 2848
rect 15936 2839 15988 2848
rect 15936 2805 15945 2839
rect 15945 2805 15979 2839
rect 15979 2805 15988 2839
rect 15936 2796 15988 2805
rect 16396 2839 16448 2848
rect 16396 2805 16405 2839
rect 16405 2805 16439 2839
rect 16439 2805 16448 2839
rect 16396 2796 16448 2805
rect 17132 2839 17184 2848
rect 17132 2805 17141 2839
rect 17141 2805 17175 2839
rect 17175 2805 17184 2839
rect 17132 2796 17184 2805
rect 18236 2796 18288 2848
rect 18788 2796 18840 2848
rect 19156 2796 19208 2848
rect 19524 2796 19576 2848
rect 20260 2796 20312 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 3148 2592 3200 2644
rect 4712 2524 4764 2576
rect 4988 2592 5040 2644
rect 6552 2592 6604 2644
rect 8024 2592 8076 2644
rect 8208 2592 8260 2644
rect 11888 2592 11940 2644
rect 12624 2592 12676 2644
rect 5264 2524 5316 2576
rect 1952 2499 2004 2508
rect 1952 2465 1961 2499
rect 1961 2465 1995 2499
rect 1995 2465 2004 2499
rect 1952 2456 2004 2465
rect 3148 2499 3200 2508
rect 3148 2465 3157 2499
rect 3157 2465 3191 2499
rect 3191 2465 3200 2499
rect 3148 2456 3200 2465
rect 3700 2456 3752 2508
rect 8484 2524 8536 2576
rect 9404 2524 9456 2576
rect 11152 2524 11204 2576
rect 12256 2524 12308 2576
rect 13912 2592 13964 2644
rect 14004 2592 14056 2644
rect 15844 2592 15896 2644
rect 16764 2592 16816 2644
rect 13636 2524 13688 2576
rect 15108 2524 15160 2576
rect 5448 2456 5500 2508
rect 5908 2499 5960 2508
rect 5908 2465 5917 2499
rect 5917 2465 5951 2499
rect 5951 2465 5960 2499
rect 6552 2499 6604 2508
rect 5908 2456 5960 2465
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 7380 2499 7432 2508
rect 7380 2465 7389 2499
rect 7389 2465 7423 2499
rect 7423 2465 7432 2499
rect 7380 2456 7432 2465
rect 8300 2456 8352 2508
rect 8576 2499 8628 2508
rect 8576 2465 8585 2499
rect 8585 2465 8619 2499
rect 8619 2465 8628 2499
rect 8576 2456 8628 2465
rect 2780 2388 2832 2440
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 3240 2388 3292 2440
rect 3516 2320 3568 2372
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 5172 2388 5224 2440
rect 7196 2388 7248 2440
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 10324 2456 10376 2508
rect 10784 2499 10836 2508
rect 10784 2465 10793 2499
rect 10793 2465 10827 2499
rect 10827 2465 10836 2499
rect 10784 2456 10836 2465
rect 13084 2499 13136 2508
rect 13084 2465 13093 2499
rect 13093 2465 13127 2499
rect 13127 2465 13136 2499
rect 13084 2456 13136 2465
rect 7564 2388 7616 2397
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 11704 2388 11756 2440
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 12164 2431 12216 2440
rect 12164 2397 12173 2431
rect 12173 2397 12207 2431
rect 12207 2397 12216 2431
rect 12900 2431 12952 2440
rect 12164 2388 12216 2397
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 14280 2456 14332 2508
rect 13360 2431 13412 2440
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 13728 2431 13780 2440
rect 13728 2397 13737 2431
rect 13737 2397 13771 2431
rect 13771 2397 13780 2431
rect 13728 2388 13780 2397
rect 13912 2388 13964 2440
rect 4988 2363 5040 2372
rect 4988 2329 4997 2363
rect 4997 2329 5031 2363
rect 5031 2329 5040 2363
rect 4988 2320 5040 2329
rect 5356 2320 5408 2372
rect 9588 2320 9640 2372
rect 5632 2295 5684 2304
rect 5632 2261 5641 2295
rect 5641 2261 5675 2295
rect 5675 2261 5684 2295
rect 5632 2252 5684 2261
rect 7748 2252 7800 2304
rect 7840 2252 7892 2304
rect 8208 2252 8260 2304
rect 9220 2252 9272 2304
rect 11244 2363 11296 2372
rect 11244 2329 11253 2363
rect 11253 2329 11287 2363
rect 11287 2329 11296 2363
rect 11244 2320 11296 2329
rect 12440 2320 12492 2372
rect 12532 2320 12584 2372
rect 15292 2456 15344 2508
rect 14740 2431 14792 2440
rect 14740 2397 14749 2431
rect 14749 2397 14783 2431
rect 14783 2397 14792 2431
rect 14740 2388 14792 2397
rect 15200 2431 15252 2440
rect 10232 2295 10284 2304
rect 10232 2261 10241 2295
rect 10241 2261 10275 2295
rect 10275 2261 10284 2295
rect 10600 2295 10652 2304
rect 10232 2252 10284 2261
rect 10600 2261 10609 2295
rect 10609 2261 10643 2295
rect 10643 2261 10652 2295
rect 10600 2252 10652 2261
rect 11152 2295 11204 2304
rect 11152 2261 11161 2295
rect 11161 2261 11195 2295
rect 11195 2261 11204 2295
rect 11152 2252 11204 2261
rect 11888 2295 11940 2304
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 12808 2252 12860 2304
rect 14648 2320 14700 2372
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 16212 2524 16264 2576
rect 17776 2592 17828 2644
rect 19616 2592 19668 2644
rect 19708 2635 19760 2644
rect 19708 2601 19717 2635
rect 19717 2601 19751 2635
rect 19751 2601 19760 2635
rect 19708 2592 19760 2601
rect 16948 2524 17000 2576
rect 18420 2524 18472 2576
rect 17132 2456 17184 2508
rect 15936 2431 15988 2440
rect 15936 2397 15945 2431
rect 15945 2397 15979 2431
rect 15979 2397 15988 2431
rect 15936 2388 15988 2397
rect 16304 2431 16356 2440
rect 16304 2397 16313 2431
rect 16313 2397 16347 2431
rect 16347 2397 16356 2431
rect 16304 2388 16356 2397
rect 16396 2388 16448 2440
rect 15108 2320 15160 2372
rect 17316 2388 17368 2440
rect 17684 2388 17736 2440
rect 18328 2456 18380 2508
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 18236 2388 18288 2440
rect 19156 2456 19208 2508
rect 20720 2499 20772 2508
rect 20720 2465 20729 2499
rect 20729 2465 20763 2499
rect 20763 2465 20772 2499
rect 20720 2456 20772 2465
rect 20904 2456 20956 2508
rect 22836 2456 22888 2508
rect 18972 2388 19024 2440
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 14556 2252 14608 2304
rect 15660 2252 15712 2304
rect 20536 2388 20588 2440
rect 16764 2252 16816 2304
rect 17592 2295 17644 2304
rect 17592 2261 17601 2295
rect 17601 2261 17635 2295
rect 17635 2261 17644 2295
rect 17592 2252 17644 2261
rect 17684 2252 17736 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 6552 2048 6604 2100
rect 10784 2048 10836 2100
rect 11888 2048 11940 2100
rect 14924 2048 14976 2100
rect 3516 1980 3568 2032
rect 6644 1980 6696 2032
rect 6736 1980 6788 2032
rect 10232 1980 10284 2032
rect 13544 1980 13596 2032
rect 16304 2048 16356 2100
rect 15384 1980 15436 2032
rect 19156 1980 19208 2032
rect 4988 1912 5040 1964
rect 7380 1912 7432 1964
rect 7748 1912 7800 1964
rect 11704 1912 11756 1964
rect 12164 1912 12216 1964
rect 13268 1912 13320 1964
rect 14280 1912 14332 1964
rect 14464 1912 14516 1964
rect 19800 1912 19852 1964
rect 5632 1844 5684 1896
rect 9404 1844 9456 1896
rect 9864 1844 9916 1896
rect 15752 1844 15804 1896
rect 4344 1776 4396 1828
rect 10876 1776 10928 1828
rect 14740 1776 14792 1828
rect 15660 1776 15712 1828
rect 3792 1708 3844 1760
rect 9772 1708 9824 1760
rect 2872 1640 2924 1692
rect 8208 1640 8260 1692
rect 11796 1640 11848 1692
rect 7932 1572 7984 1624
rect 9588 1572 9640 1624
rect 5816 1368 5868 1420
rect 6276 1368 6328 1420
rect 16580 1368 16632 1420
rect 17592 1368 17644 1420
rect 4620 1232 4672 1284
rect 15568 1232 15620 1284
rect 848 1164 900 1216
rect 11152 1164 11204 1216
rect 1676 1096 1728 1148
rect 13176 1096 13228 1148
<< metal2 >>
rect 18 22536 74 22545
rect 18 22471 74 22480
rect 32 8022 60 22471
rect 308 22222 520 22250
rect 112 19440 164 19446
rect 112 19382 164 19388
rect 124 16182 152 19382
rect 204 19372 256 19378
rect 204 19314 256 19320
rect 112 16176 164 16182
rect 112 16118 164 16124
rect 216 15570 244 19314
rect 204 15564 256 15570
rect 204 15506 256 15512
rect 308 15434 336 22222
rect 492 22114 520 22222
rect 570 22200 626 23000
rect 938 22200 994 23000
rect 1306 22200 1362 23000
rect 1582 22264 1638 22273
rect 584 22114 612 22200
rect 492 22086 612 22114
rect 952 19446 980 22200
rect 1032 21140 1084 21146
rect 1032 21082 1084 21088
rect 940 19440 992 19446
rect 940 19382 992 19388
rect 296 15428 348 15434
rect 296 15370 348 15376
rect 938 14376 994 14385
rect 124 14334 938 14362
rect 20 8016 72 8022
rect 20 7958 72 7964
rect 124 6798 152 14334
rect 938 14311 994 14320
rect 848 13252 900 13258
rect 848 13194 900 13200
rect 860 10554 888 13194
rect 1044 12434 1072 21082
rect 1320 19378 1348 22200
rect 1582 22199 1638 22208
rect 1674 22200 1730 23000
rect 2042 22200 2098 23000
rect 2410 22200 2466 23000
rect 2778 22200 2834 23000
rect 2884 22222 3096 22250
rect 1492 20256 1544 20262
rect 1490 20224 1492 20233
rect 1544 20224 1546 20233
rect 1490 20159 1546 20168
rect 1400 19780 1452 19786
rect 1400 19722 1452 19728
rect 1308 19372 1360 19378
rect 1308 19314 1360 19320
rect 1216 18352 1268 18358
rect 1216 18294 1268 18300
rect 1122 16280 1178 16289
rect 1122 16215 1178 16224
rect 676 10526 888 10554
rect 952 12406 1072 12434
rect 112 6792 164 6798
rect 112 6734 164 6740
rect 676 2774 704 10526
rect 952 10282 980 12406
rect 860 10254 980 10282
rect 860 2922 888 10254
rect 1136 10248 1164 16215
rect 1044 10220 1164 10248
rect 940 8016 992 8022
rect 938 7984 940 7993
rect 992 7984 994 7993
rect 938 7919 994 7928
rect 952 7478 980 7919
rect 940 7472 992 7478
rect 940 7414 992 7420
rect 940 6792 992 6798
rect 938 6760 940 6769
rect 992 6760 994 6769
rect 938 6695 994 6704
rect 952 5846 980 6695
rect 1044 6225 1072 10220
rect 1228 10146 1256 18294
rect 1412 16522 1440 19722
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1504 19417 1532 19654
rect 1596 19514 1624 22199
rect 1688 21162 1716 22200
rect 1950 21448 2006 21457
rect 1950 21383 2006 21392
rect 1688 21134 1808 21162
rect 1676 21072 1728 21078
rect 1676 21014 1728 21020
rect 1688 20466 1716 21014
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 1780 19938 1808 21134
rect 1858 20632 1914 20641
rect 1858 20567 1860 20576
rect 1912 20567 1914 20576
rect 1860 20538 1912 20544
rect 1964 20058 1992 21383
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 1780 19910 1992 19938
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1858 19816 1914 19825
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 19009 1532 19110
rect 1490 19000 1546 19009
rect 1688 18970 1716 19314
rect 1490 18935 1546 18944
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1780 18902 1808 19790
rect 1858 19751 1914 19760
rect 1872 19718 1900 19751
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1964 19530 1992 19910
rect 1872 19502 1992 19530
rect 1768 18896 1820 18902
rect 1768 18838 1820 18844
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1504 18193 1532 18566
rect 1490 18184 1546 18193
rect 1490 18119 1546 18128
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17785 1532 18022
rect 1688 17882 1716 18702
rect 1780 18426 1808 18702
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1490 17776 1546 17785
rect 1490 17711 1546 17720
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17377 1532 17478
rect 1490 17368 1546 17377
rect 1490 17303 1546 17312
rect 1492 16992 1544 16998
rect 1490 16960 1492 16969
rect 1544 16960 1546 16969
rect 1490 16895 1546 16904
rect 1688 16794 1716 17614
rect 1780 17338 1808 18226
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1400 16516 1452 16522
rect 1400 16458 1452 16464
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1504 16153 1532 16390
rect 1688 16250 1716 16526
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1490 16144 1546 16153
rect 1490 16079 1546 16088
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15745 1532 15846
rect 1490 15736 1546 15745
rect 1780 15706 1808 17138
rect 1872 16998 1900 19502
rect 1950 19408 2006 19417
rect 1950 19343 1952 19352
rect 2004 19343 2006 19352
rect 1952 19314 2004 19320
rect 1952 18624 2004 18630
rect 1950 18592 1952 18601
rect 2004 18592 2006 18601
rect 1950 18527 2006 18536
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1964 17338 1992 18226
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1858 16552 1914 16561
rect 1858 16487 1914 16496
rect 1872 16454 1900 16487
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1490 15671 1546 15680
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1872 15586 1900 15982
rect 1964 15706 1992 16050
rect 2056 15978 2084 22200
rect 2226 21040 2282 21049
rect 2226 20975 2282 20984
rect 2136 20868 2188 20874
rect 2136 20810 2188 20816
rect 2148 20466 2176 20810
rect 2240 20602 2268 20975
rect 2424 20618 2452 22200
rect 2792 22114 2820 22200
rect 2884 22114 2912 22222
rect 2792 22086 2912 22114
rect 2228 20596 2280 20602
rect 2424 20590 2544 20618
rect 2228 20538 2280 20544
rect 2410 20496 2466 20505
rect 2136 20460 2188 20466
rect 2410 20431 2412 20440
rect 2136 20402 2188 20408
rect 2464 20431 2466 20440
rect 2412 20402 2464 20408
rect 2410 19952 2466 19961
rect 2410 19887 2466 19896
rect 2424 19854 2452 19887
rect 2412 19848 2464 19854
rect 2412 19790 2464 19796
rect 2228 19780 2280 19786
rect 2228 19722 2280 19728
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 2148 17610 2176 18022
rect 2240 17626 2268 19722
rect 2516 18970 2544 20590
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 2608 18873 2636 19790
rect 2688 18964 2740 18970
rect 2688 18906 2740 18912
rect 2594 18864 2650 18873
rect 2594 18799 2650 18808
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2504 18692 2556 18698
rect 2504 18634 2556 18640
rect 2412 17876 2464 17882
rect 2412 17818 2464 17824
rect 2136 17604 2188 17610
rect 2240 17598 2360 17626
rect 2136 17546 2188 17552
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2044 15972 2096 15978
rect 2044 15914 2096 15920
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1872 15558 1992 15586
rect 1492 15360 1544 15366
rect 1490 15328 1492 15337
rect 1544 15328 1546 15337
rect 1490 15263 1546 15272
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1504 14521 1532 14758
rect 1688 14618 1716 14962
rect 1858 14920 1914 14929
rect 1858 14855 1860 14864
rect 1912 14855 1914 14864
rect 1860 14826 1912 14832
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1490 14512 1546 14521
rect 1490 14447 1546 14456
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 14113 1532 14214
rect 1490 14104 1546 14113
rect 1490 14039 1546 14048
rect 1964 13977 1992 15558
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2056 14550 2084 14962
rect 2044 14544 2096 14550
rect 2044 14486 2096 14492
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2056 14249 2084 14350
rect 2042 14240 2098 14249
rect 2042 14175 2098 14184
rect 1950 13968 2006 13977
rect 2148 13954 2176 17138
rect 2228 17128 2280 17134
rect 2226 17096 2228 17105
rect 2280 17096 2282 17105
rect 2226 17031 2282 17040
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2240 15706 2268 16526
rect 2332 16250 2360 17598
rect 2424 16250 2452 17818
rect 2516 16726 2544 18634
rect 2608 17649 2636 18702
rect 2594 17640 2650 17649
rect 2594 17575 2650 17584
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2608 17377 2636 17478
rect 2594 17368 2650 17377
rect 2594 17303 2650 17312
rect 2504 16720 2556 16726
rect 2504 16662 2556 16668
rect 2596 16584 2648 16590
rect 2596 16526 2648 16532
rect 2504 16516 2556 16522
rect 2504 16458 2556 16464
rect 2516 16425 2544 16458
rect 2502 16416 2558 16425
rect 2502 16351 2558 16360
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2608 16017 2636 16526
rect 2700 16114 2728 18906
rect 2792 18358 2820 20198
rect 2884 19990 2912 20266
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 2872 19984 2924 19990
rect 2872 19926 2924 19932
rect 2976 19689 3004 20198
rect 2962 19680 3018 19689
rect 2962 19615 3018 19624
rect 2962 19544 3018 19553
rect 2872 19508 2924 19514
rect 2962 19479 3018 19488
rect 2872 19450 2924 19456
rect 2884 18970 2912 19450
rect 2976 19378 3004 19479
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2964 18896 3016 18902
rect 2964 18838 3016 18844
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2780 17536 2832 17542
rect 2780 17478 2832 17484
rect 2792 16794 2820 17478
rect 2884 17338 2912 18566
rect 2976 18358 3004 18838
rect 2964 18352 3016 18358
rect 2964 18294 3016 18300
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2976 17218 3004 18294
rect 3068 17762 3096 22222
rect 3146 22200 3202 23000
rect 3514 22200 3570 23000
rect 3882 22200 3938 23000
rect 4250 22200 4306 23000
rect 4618 22200 4674 23000
rect 4986 22200 5042 23000
rect 5354 22200 5410 23000
rect 5722 22200 5778 23000
rect 6090 22200 6146 23000
rect 6196 22222 6408 22250
rect 3160 19446 3188 22200
rect 3238 21312 3294 21321
rect 3238 21247 3294 21256
rect 3252 19990 3280 21247
rect 3330 21040 3386 21049
rect 3330 20975 3386 20984
rect 3344 19990 3372 20975
rect 3528 20584 3556 22200
rect 3528 20556 3648 20584
rect 3620 20466 3648 20556
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3528 20369 3556 20402
rect 3514 20360 3570 20369
rect 3514 20295 3570 20304
rect 3424 20256 3476 20262
rect 3424 20198 3476 20204
rect 3240 19984 3292 19990
rect 3240 19926 3292 19932
rect 3332 19984 3384 19990
rect 3332 19926 3384 19932
rect 3332 19780 3384 19786
rect 3332 19722 3384 19728
rect 3344 19514 3372 19722
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3148 19440 3200 19446
rect 3200 19388 3280 19394
rect 3148 19382 3280 19388
rect 3160 19366 3280 19382
rect 3252 19281 3280 19366
rect 3332 19304 3384 19310
rect 3238 19272 3294 19281
rect 3332 19246 3384 19252
rect 3238 19207 3294 19216
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3160 18834 3188 19110
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3252 18766 3280 19110
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 3344 18630 3372 19246
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3332 18352 3384 18358
rect 3436 18329 3464 20198
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3896 20058 3924 22200
rect 4158 21856 4214 21865
rect 4158 21791 4214 21800
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 3988 20534 4016 20742
rect 3976 20528 4028 20534
rect 3976 20470 4028 20476
rect 4068 20460 4120 20466
rect 4068 20402 4120 20408
rect 3976 20324 4028 20330
rect 3976 20266 4028 20272
rect 3988 20233 4016 20266
rect 3974 20224 4030 20233
rect 3974 20159 4030 20168
rect 3884 20052 3936 20058
rect 3936 20012 4016 20040
rect 3884 19994 3936 20000
rect 3608 19780 3660 19786
rect 3608 19722 3660 19728
rect 3620 19281 3648 19722
rect 3792 19508 3844 19514
rect 3712 19468 3792 19496
rect 3712 19310 3740 19468
rect 3792 19450 3844 19456
rect 3700 19304 3752 19310
rect 3606 19272 3662 19281
rect 3700 19246 3752 19252
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3606 19207 3662 19216
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3896 18873 3924 19246
rect 3882 18864 3938 18873
rect 3700 18828 3752 18834
rect 3882 18799 3938 18808
rect 3700 18770 3752 18776
rect 3332 18294 3384 18300
rect 3422 18320 3478 18329
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3068 17734 3188 17762
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 2884 17190 3004 17218
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2884 16658 2912 17190
rect 3068 17134 3096 17546
rect 3160 17542 3188 17734
rect 3252 17678 3280 18022
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3252 17202 3280 17614
rect 3344 17338 3372 18294
rect 3712 18290 3740 18770
rect 3988 18290 4016 20012
rect 4080 18737 4108 20402
rect 4066 18728 4122 18737
rect 4066 18663 4122 18672
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 3422 18255 3478 18264
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3516 18216 3568 18222
rect 3436 18176 3516 18204
rect 3436 17882 3464 18176
rect 3516 18158 3568 18164
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3436 17270 3464 17818
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3606 17640 3662 17649
rect 3424 17264 3476 17270
rect 3424 17206 3476 17212
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2594 16008 2650 16017
rect 2594 15943 2650 15952
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2792 15638 2820 15846
rect 2780 15632 2832 15638
rect 2318 15600 2374 15609
rect 2780 15574 2832 15580
rect 2884 15570 2912 16594
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 2976 15706 3004 16458
rect 3068 16046 3096 17070
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 3160 15978 3188 17138
rect 3528 17082 3556 17614
rect 3606 17575 3662 17584
rect 3252 17054 3556 17082
rect 3252 16130 3280 17054
rect 3620 16980 3648 17575
rect 3436 16952 3648 16980
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3344 16250 3372 16390
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3252 16102 3372 16130
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3148 15972 3200 15978
rect 3148 15914 3200 15920
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2318 15535 2374 15544
rect 2872 15564 2924 15570
rect 2332 15502 2360 15535
rect 2872 15506 2924 15512
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2240 14618 2268 15438
rect 2412 15428 2464 15434
rect 2412 15370 2464 15376
rect 2424 15162 2452 15370
rect 2608 15201 2636 15438
rect 2594 15192 2650 15201
rect 2412 15156 2464 15162
rect 2594 15127 2650 15136
rect 2412 15098 2464 15104
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2792 14550 2820 15438
rect 2884 14890 2912 15506
rect 3068 15502 3096 15846
rect 3252 15706 3280 15982
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2872 14884 2924 14890
rect 2872 14826 2924 14832
rect 2976 14618 3004 15438
rect 3344 15366 3372 16102
rect 3056 15360 3108 15366
rect 3054 15328 3056 15337
rect 3332 15360 3384 15366
rect 3108 15328 3110 15337
rect 3332 15302 3384 15308
rect 3054 15263 3110 15272
rect 3238 15056 3294 15065
rect 3238 14991 3294 15000
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 3252 14482 3280 14991
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2424 14074 2452 14350
rect 3436 14074 3464 16952
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3896 16250 3924 18226
rect 4080 18170 4108 18566
rect 3988 18142 4108 18170
rect 3988 16590 4016 18142
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4080 17202 4108 17478
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3896 14346 3924 15914
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3240 14000 3292 14006
rect 2148 13926 2636 13954
rect 3240 13942 3292 13948
rect 1950 13903 2006 13912
rect 2504 13796 2556 13802
rect 2504 13738 2556 13744
rect 1492 13728 1544 13734
rect 1490 13696 1492 13705
rect 2320 13728 2372 13734
rect 1544 13696 1546 13705
rect 2320 13670 2372 13676
rect 1490 13631 1546 13640
rect 1676 13320 1728 13326
rect 1490 13288 1546 13297
rect 1676 13262 1728 13268
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 1490 13223 1546 13232
rect 1504 13190 1532 13223
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1688 12986 1716 13262
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1872 12889 1900 13126
rect 1858 12880 1914 12889
rect 1858 12815 1914 12824
rect 1490 12472 1546 12481
rect 1490 12407 1492 12416
rect 1544 12407 1546 12416
rect 1492 12378 1544 12384
rect 1306 12336 1362 12345
rect 1306 12271 1362 12280
rect 1136 10118 1256 10146
rect 1136 8022 1164 10118
rect 1214 9480 1270 9489
rect 1214 9415 1270 9424
rect 1228 8401 1256 9415
rect 1214 8392 1270 8401
rect 1214 8327 1270 8336
rect 1124 8016 1176 8022
rect 1124 7958 1176 7964
rect 1228 6798 1256 8327
rect 1216 6792 1268 6798
rect 1216 6734 1268 6740
rect 1030 6216 1086 6225
rect 1030 6151 1086 6160
rect 940 5840 992 5846
rect 940 5782 992 5788
rect 1044 5030 1072 6151
rect 1122 5944 1178 5953
rect 1122 5879 1178 5888
rect 1032 5024 1084 5030
rect 1032 4966 1084 4972
rect 1136 4622 1164 5879
rect 1214 5264 1270 5273
rect 1214 5199 1270 5208
rect 1124 4616 1176 4622
rect 1124 4558 1176 4564
rect 1228 4162 1256 5199
rect 1320 4865 1348 12271
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1492 12164 1544 12170
rect 1492 12106 1544 12112
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1412 9586 1440 11494
rect 1504 11257 1532 12106
rect 1860 12096 1912 12102
rect 1858 12064 1860 12073
rect 1912 12064 1914 12073
rect 1858 11999 1914 12008
rect 1860 11620 1912 11626
rect 1860 11562 1912 11568
rect 1674 11384 1730 11393
rect 1674 11319 1730 11328
rect 1688 11286 1716 11319
rect 1676 11280 1728 11286
rect 1490 11248 1546 11257
rect 1676 11222 1728 11228
rect 1490 11183 1546 11192
rect 1504 11150 1532 11183
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1872 11082 1900 11562
rect 1964 11354 1992 12174
rect 2056 11506 2084 13262
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12918 2268 13126
rect 2228 12912 2280 12918
rect 2228 12854 2280 12860
rect 2136 12232 2188 12238
rect 2332 12209 2360 13670
rect 2410 13152 2466 13161
rect 2410 13087 2466 13096
rect 2136 12174 2188 12180
rect 2318 12200 2374 12209
rect 2148 11778 2176 12174
rect 2318 12135 2374 12144
rect 2332 11898 2360 12135
rect 2424 11898 2452 13087
rect 2516 12646 2544 13738
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2516 12238 2544 12582
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2148 11750 2360 11778
rect 2228 11688 2280 11694
rect 2226 11656 2228 11665
rect 2280 11656 2282 11665
rect 2226 11591 2282 11600
rect 2056 11478 2268 11506
rect 2042 11384 2098 11393
rect 1952 11348 2004 11354
rect 2042 11319 2098 11328
rect 1952 11290 2004 11296
rect 2056 11200 2084 11319
rect 1964 11172 2084 11200
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1872 10849 1900 11018
rect 1858 10840 1914 10849
rect 1858 10775 1914 10784
rect 1768 10736 1820 10742
rect 1768 10678 1820 10684
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1504 10130 1532 10406
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1504 9625 1532 10066
rect 1582 10024 1638 10033
rect 1582 9959 1638 9968
rect 1490 9616 1546 9625
rect 1400 9580 1452 9586
rect 1490 9551 1546 9560
rect 1400 9522 1452 9528
rect 1596 9500 1624 9959
rect 1780 9722 1808 10678
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1872 9926 1900 10610
rect 1964 10441 1992 11172
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 2056 10713 2084 11018
rect 2042 10704 2098 10713
rect 2042 10639 2098 10648
rect 2240 10470 2268 11478
rect 2228 10464 2280 10470
rect 1950 10432 2006 10441
rect 2228 10406 2280 10412
rect 1950 10367 2006 10376
rect 1964 9994 1992 10367
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 2056 9926 2084 10066
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1872 9518 1900 9862
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2148 9602 2176 9658
rect 2044 9580 2096 9586
rect 2148 9574 2268 9602
rect 2044 9522 2096 9528
rect 1504 9472 1624 9500
rect 1860 9512 1912 9518
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1412 8498 1440 9143
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1412 7177 1440 8191
rect 1504 7886 1532 9472
rect 1860 9454 1912 9460
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 9042 1716 9318
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1582 8664 1638 8673
rect 1582 8599 1584 8608
rect 1636 8599 1638 8608
rect 1584 8570 1636 8576
rect 1688 7954 1716 8978
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1582 7848 1638 7857
rect 1582 7783 1638 7792
rect 1596 7750 1624 7783
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1780 7546 1808 8774
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1872 7954 1900 8230
rect 2056 8090 2084 9522
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2148 9178 2176 9454
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 1860 7948 1912 7954
rect 1860 7890 1912 7896
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1860 7336 1912 7342
rect 1674 7304 1730 7313
rect 1860 7278 1912 7284
rect 1674 7239 1676 7248
rect 1728 7239 1730 7248
rect 1676 7210 1728 7216
rect 1768 7200 1820 7206
rect 1398 7168 1454 7177
rect 1768 7142 1820 7148
rect 1398 7103 1454 7112
rect 1412 5778 1440 7103
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1596 6662 1624 6831
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1504 5914 1532 6054
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1504 5817 1532 5850
rect 1490 5808 1546 5817
rect 1400 5772 1452 5778
rect 1490 5743 1546 5752
rect 1676 5772 1728 5778
rect 1400 5714 1452 5720
rect 1676 5714 1728 5720
rect 1584 5296 1636 5302
rect 1584 5238 1636 5244
rect 1306 4856 1362 4865
rect 1596 4826 1624 5238
rect 1306 4791 1362 4800
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1228 4134 1440 4162
rect 1412 3233 1440 4134
rect 1688 4078 1716 5714
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1490 3768 1546 3777
rect 1490 3703 1546 3712
rect 1504 3534 1532 3703
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1398 3224 1454 3233
rect 1398 3159 1454 3168
rect 848 2916 900 2922
rect 848 2858 900 2864
rect 676 2746 888 2774
rect 860 1222 888 2746
rect 848 1216 900 1222
rect 848 1158 900 1164
rect 1688 1154 1716 3606
rect 1676 1148 1728 1154
rect 1676 1090 1728 1096
rect 1504 870 1624 898
rect 1504 800 1532 870
rect 1490 0 1546 800
rect 1596 762 1624 870
rect 1780 762 1808 7142
rect 1872 6866 1900 7278
rect 2056 7002 2084 7686
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 2042 6896 2098 6905
rect 1860 6860 1912 6866
rect 2042 6831 2098 6840
rect 1860 6802 1912 6808
rect 2056 6730 2084 6831
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 1872 4282 1900 6666
rect 2042 6488 2098 6497
rect 2042 6423 2098 6432
rect 1950 5400 2006 5409
rect 1950 5335 2006 5344
rect 1964 5234 1992 5335
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1950 4992 2006 5001
rect 1950 4927 2006 4936
rect 1964 4622 1992 4927
rect 2056 4758 2084 6423
rect 2148 5574 2176 8570
rect 2240 5642 2268 9574
rect 2332 6118 2360 11750
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2424 9450 2452 11698
rect 2504 11620 2556 11626
rect 2504 11562 2556 11568
rect 2516 11150 2544 11562
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2516 10810 2544 11086
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2424 8430 2452 8978
rect 2516 8838 2544 9046
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2516 8673 2544 8774
rect 2502 8664 2558 8673
rect 2502 8599 2558 8608
rect 2608 8430 2636 13926
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2700 9110 2728 11834
rect 2792 11830 2820 13126
rect 3252 12986 3280 13942
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3344 12986 3372 13806
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2884 12238 2912 12718
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2792 10810 2820 11630
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2884 10690 2912 11766
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2792 10662 2912 10690
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2424 7342 2452 8366
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2516 7546 2544 7754
rect 2594 7712 2650 7721
rect 2594 7647 2650 7656
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2608 7018 2636 7647
rect 2424 6990 2636 7018
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2228 5636 2280 5642
rect 2228 5578 2280 5584
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2044 4752 2096 4758
rect 2044 4694 2096 4700
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1872 800 1900 3538
rect 1964 2514 1992 4558
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 2056 3738 2084 4422
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 2148 3058 2176 5510
rect 2424 5352 2452 6990
rect 2700 6633 2728 8910
rect 2792 8514 2820 10662
rect 2976 10606 3004 11018
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2976 10266 3004 10542
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2976 9450 3004 9930
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2884 8945 2912 9318
rect 2870 8936 2926 8945
rect 2976 8906 3004 9386
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 8974 3096 9318
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2870 8871 2926 8880
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 3068 8809 3096 8910
rect 3054 8800 3110 8809
rect 3054 8735 3110 8744
rect 2870 8528 2926 8537
rect 2792 8486 2870 8514
rect 2870 8463 2872 8472
rect 2924 8463 2926 8472
rect 2872 8434 2924 8440
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2792 8242 2820 8366
rect 2872 8288 2924 8294
rect 2792 8236 2872 8242
rect 2792 8230 2924 8236
rect 2792 8214 2912 8230
rect 2792 7546 2820 8214
rect 2976 8090 3004 8366
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 3160 8022 3188 10950
rect 3252 9489 3280 12310
rect 3344 12306 3372 12786
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3436 11898 3464 13874
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3896 13274 3924 13874
rect 3988 13734 4016 16118
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4080 15570 4108 15982
rect 4172 15706 4200 21791
rect 4264 19718 4292 22200
rect 4528 20936 4580 20942
rect 4528 20878 4580 20884
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4264 19258 4292 19654
rect 4356 19378 4384 20538
rect 4540 20398 4568 20878
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 4632 19768 4660 22200
rect 4802 21176 4858 21185
rect 4802 21111 4858 21120
rect 4540 19740 4660 19768
rect 4712 19780 4764 19786
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4264 19230 4384 19258
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4264 17785 4292 19110
rect 4250 17776 4306 17785
rect 4250 17711 4306 17720
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4264 16590 4292 17614
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4066 15464 4122 15473
rect 4066 15399 4122 15408
rect 4080 15094 4108 15399
rect 4160 15360 4212 15366
rect 4158 15328 4160 15337
rect 4212 15328 4214 15337
rect 4158 15263 4214 15272
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 4264 15026 4292 16526
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4066 13968 4122 13977
rect 4264 13938 4292 14962
rect 4356 14822 4384 19230
rect 4448 17882 4476 19314
rect 4540 18465 4568 19740
rect 4712 19722 4764 19728
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 4526 18456 4582 18465
rect 4526 18391 4582 18400
rect 4632 18086 4660 19246
rect 4724 18630 4752 19722
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4724 18222 4752 18566
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4540 17921 4568 18022
rect 4526 17912 4582 17921
rect 4436 17876 4488 17882
rect 4816 17864 4844 21111
rect 4894 20904 4950 20913
rect 4894 20839 4950 20848
rect 4908 20330 4936 20839
rect 5000 20754 5028 22200
rect 5000 20726 5212 20754
rect 5184 20534 5212 20726
rect 5172 20528 5224 20534
rect 5172 20470 5224 20476
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 4896 20324 4948 20330
rect 4896 20266 4948 20272
rect 5092 19145 5120 20402
rect 5078 19136 5134 19145
rect 5078 19071 5134 19080
rect 5080 18352 5132 18358
rect 5080 18294 5132 18300
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4526 17847 4582 17856
rect 4436 17818 4488 17824
rect 4632 17836 4844 17864
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4448 17270 4476 17682
rect 4526 17640 4582 17649
rect 4526 17575 4582 17584
rect 4540 17542 4568 17575
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 4436 17264 4488 17270
rect 4436 17206 4488 17212
rect 4448 16590 4476 17206
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4448 14872 4476 16390
rect 4540 15881 4568 16730
rect 4526 15872 4582 15881
rect 4526 15807 4582 15816
rect 4632 15688 4660 17836
rect 4710 17776 4766 17785
rect 4710 17711 4766 17720
rect 4724 16590 4752 17711
rect 4908 17066 4936 18022
rect 5000 17338 5028 18226
rect 5092 17882 5120 18294
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 5078 17640 5134 17649
rect 5078 17575 5134 17584
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4896 17060 4948 17066
rect 4896 17002 4948 17008
rect 5092 16998 5120 17575
rect 5184 17241 5212 20470
rect 5276 19514 5304 20470
rect 5368 20466 5396 22200
rect 5736 20754 5764 22200
rect 6104 22114 6132 22200
rect 6196 22114 6224 22222
rect 6104 22086 6224 22114
rect 6380 20890 6408 22222
rect 6458 22200 6514 23000
rect 6564 22222 6776 22250
rect 6472 22114 6500 22200
rect 6564 22114 6592 22222
rect 6472 22086 6592 22114
rect 6380 20862 6592 20890
rect 5736 20726 5948 20754
rect 5816 20596 5868 20602
rect 5816 20538 5868 20544
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 5368 19825 5396 20266
rect 5460 20233 5488 20334
rect 5724 20256 5776 20262
rect 5446 20224 5502 20233
rect 5724 20198 5776 20204
rect 5446 20159 5502 20168
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 5354 19816 5410 19825
rect 5552 19786 5580 19994
rect 5736 19854 5764 20198
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5354 19751 5410 19760
rect 5540 19780 5592 19786
rect 5540 19722 5592 19728
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5552 19310 5580 19722
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5644 19242 5672 19654
rect 5632 19236 5684 19242
rect 5632 19178 5684 19184
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5460 18290 5488 18906
rect 5736 18902 5764 19790
rect 5724 18896 5776 18902
rect 5724 18838 5776 18844
rect 5828 18714 5856 20538
rect 5920 19281 5948 20726
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6092 19712 6144 19718
rect 6012 19672 6092 19700
rect 6012 19553 6040 19672
rect 6092 19654 6144 19660
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 5998 19544 6054 19553
rect 6148 19547 6456 19556
rect 5998 19479 6000 19488
rect 6052 19479 6054 19488
rect 6000 19450 6052 19456
rect 6012 19419 6040 19450
rect 5906 19272 5962 19281
rect 5906 19207 5962 19216
rect 5920 18970 5948 19207
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 5736 18686 5856 18714
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 5908 18692 5960 18698
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5644 18426 5672 18566
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5736 18306 5764 18686
rect 5908 18634 5960 18640
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5644 18278 5764 18306
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5354 17776 5410 17785
rect 5354 17711 5410 17720
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 5170 17232 5226 17241
rect 5170 17167 5226 17176
rect 5276 17066 5304 17614
rect 5368 17202 5396 17711
rect 5460 17678 5488 18090
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5552 17610 5580 18158
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5264 17060 5316 17066
rect 5264 17002 5316 17008
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 4816 16794 4844 16934
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 5368 16697 5396 17138
rect 5354 16688 5410 16697
rect 5354 16623 5410 16632
rect 5552 16640 5580 17546
rect 5644 16810 5672 18278
rect 5722 17368 5778 17377
rect 5722 17303 5778 17312
rect 5736 16969 5764 17303
rect 5722 16960 5778 16969
rect 5722 16895 5778 16904
rect 5644 16782 5764 16810
rect 5632 16652 5684 16658
rect 5552 16612 5632 16640
rect 5632 16594 5684 16600
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4988 16516 5040 16522
rect 4988 16458 5040 16464
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4540 15660 4660 15688
rect 4540 15201 4568 15660
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4526 15192 4582 15201
rect 4526 15127 4582 15136
rect 4540 15026 4568 15127
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4528 14884 4580 14890
rect 4448 14844 4528 14872
rect 4528 14826 4580 14832
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4436 14272 4488 14278
rect 4436 14214 4488 14220
rect 4066 13903 4068 13912
rect 4120 13903 4122 13912
rect 4252 13932 4304 13938
rect 4068 13874 4120 13880
rect 4252 13874 4304 13880
rect 4160 13864 4212 13870
rect 4158 13832 4160 13841
rect 4212 13832 4214 13841
rect 4158 13767 4214 13776
rect 4252 13796 4304 13802
rect 4252 13738 4304 13744
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3804 13246 3924 13274
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 3804 12646 3832 13246
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3896 12434 3924 13126
rect 3988 12866 4016 13262
rect 4080 13161 4108 13262
rect 4066 13152 4122 13161
rect 4066 13087 4122 13096
rect 4264 12918 4292 13738
rect 4356 13462 4384 14214
rect 4448 13530 4476 14214
rect 4540 13734 4568 14826
rect 4632 13841 4660 15506
rect 4618 13832 4674 13841
rect 4618 13767 4674 13776
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4344 13456 4396 13462
rect 4344 13398 4396 13404
rect 4540 13394 4568 13466
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 4356 13161 4384 13194
rect 4342 13152 4398 13161
rect 4342 13087 4398 13096
rect 4252 12912 4304 12918
rect 4158 12880 4214 12889
rect 3988 12838 4108 12866
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3988 12442 4016 12582
rect 3804 12406 3924 12434
rect 3976 12436 4028 12442
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3712 12073 3740 12242
rect 3698 12064 3754 12073
rect 3698 11999 3754 12008
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3344 9722 3372 11154
rect 3436 11082 3464 11698
rect 3804 11558 3832 12406
rect 3976 12378 4028 12384
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3896 11694 3924 12242
rect 4080 12238 4108 12838
rect 4252 12854 4304 12860
rect 4158 12815 4214 12824
rect 4172 12374 4200 12815
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4264 12442 4292 12650
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 4080 11626 4108 12174
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 4172 11370 4200 12038
rect 4356 11898 4384 12718
rect 4344 11892 4396 11898
rect 4448 11880 4476 13194
rect 4540 12306 4568 13330
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4632 12753 4660 12786
rect 4618 12744 4674 12753
rect 4724 12714 4752 16050
rect 5000 15706 5028 16458
rect 5078 16416 5134 16425
rect 5078 16351 5134 16360
rect 5092 16046 5120 16351
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 5092 15570 5120 15982
rect 5368 15706 5396 16050
rect 5644 16046 5672 16594
rect 5448 16040 5500 16046
rect 5632 16040 5684 16046
rect 5500 15988 5580 15994
rect 5448 15982 5580 15988
rect 5632 15982 5684 15988
rect 5460 15966 5580 15982
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 5354 15464 5410 15473
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4816 14618 4844 14962
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4908 13954 4936 15302
rect 5000 14346 5028 15438
rect 5354 15399 5356 15408
rect 5408 15399 5410 15408
rect 5356 15370 5408 15376
rect 5552 15094 5580 15966
rect 5736 15706 5764 16782
rect 5828 16454 5856 18566
rect 5920 17882 5948 18634
rect 6012 18426 6040 18702
rect 6288 18698 6316 19110
rect 6276 18692 6328 18698
rect 6276 18634 6328 18640
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6564 18358 6592 20862
rect 6748 20806 6776 22222
rect 6826 22200 6882 23000
rect 7194 22200 7250 23000
rect 7562 22200 7618 23000
rect 7668 22222 7880 22250
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6840 20602 6868 22200
rect 7208 20618 7236 22200
rect 7576 22114 7604 22200
rect 7668 22114 7696 22222
rect 7576 22086 7696 22114
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 7024 20590 7236 20618
rect 6644 20528 6696 20534
rect 6696 20476 6868 20482
rect 6644 20470 6868 20476
rect 6656 20466 6868 20470
rect 6656 20460 6880 20466
rect 6656 20454 6828 20460
rect 6828 20402 6880 20408
rect 6644 20392 6696 20398
rect 7024 20369 7052 20590
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 7472 20528 7524 20534
rect 7472 20470 7524 20476
rect 7104 20392 7156 20398
rect 6644 20334 6696 20340
rect 7010 20360 7066 20369
rect 6552 18352 6604 18358
rect 6552 18294 6604 18300
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 5908 17876 5960 17882
rect 5960 17836 6040 17864
rect 5908 17818 5960 17824
rect 5908 17604 5960 17610
rect 5908 17546 5960 17552
rect 5920 17338 5948 17546
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 5920 16250 5948 17138
rect 6012 17134 6040 17836
rect 6104 17542 6132 18158
rect 6380 17814 6408 18226
rect 6656 17882 6684 20334
rect 6828 20324 6880 20330
rect 7104 20334 7156 20340
rect 7010 20295 7066 20304
rect 6828 20266 6880 20272
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6748 18766 6776 19994
rect 6736 18760 6788 18766
rect 6736 18702 6788 18708
rect 6736 18148 6788 18154
rect 6736 18090 6788 18096
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6368 17808 6420 17814
rect 6368 17750 6420 17756
rect 6458 17776 6514 17785
rect 6458 17711 6514 17720
rect 6552 17740 6604 17746
rect 6472 17610 6500 17711
rect 6552 17682 6604 17688
rect 6460 17604 6512 17610
rect 6460 17546 6512 17552
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 6000 17128 6052 17134
rect 6000 17070 6052 17076
rect 6196 16590 6224 17274
rect 6564 16658 6592 17682
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6656 16794 6684 17478
rect 6748 17066 6776 18090
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6184 16584 6236 16590
rect 6840 16538 6868 20266
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 6184 16526 6236 16532
rect 6748 16510 6868 16538
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 5998 16280 6054 16289
rect 6148 16283 6456 16292
rect 5908 16244 5960 16250
rect 5998 16215 6054 16224
rect 5908 16186 5960 16192
rect 6012 16182 6040 16215
rect 6000 16176 6052 16182
rect 6000 16118 6052 16124
rect 5998 16008 6054 16017
rect 5998 15943 6054 15952
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5906 15600 5962 15609
rect 6012 15570 6040 15943
rect 6642 15600 6698 15609
rect 5906 15535 5962 15544
rect 6000 15564 6052 15570
rect 5920 15348 5948 15535
rect 6642 15535 6698 15544
rect 6000 15506 6052 15512
rect 6000 15360 6052 15366
rect 5920 15320 6000 15348
rect 6000 15302 6052 15308
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 5906 15192 5962 15201
rect 5906 15127 5962 15136
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5722 15056 5778 15065
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5276 14618 5304 14894
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 4988 14340 5040 14346
rect 4988 14282 5040 14288
rect 5000 14074 5028 14282
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4816 13394 4844 13942
rect 4908 13926 5212 13954
rect 4988 13728 5040 13734
rect 5040 13688 5120 13716
rect 4988 13670 5040 13676
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4618 12679 4674 12688
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4710 12608 4766 12617
rect 4710 12543 4766 12552
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4724 12238 4752 12543
rect 4908 12238 4936 12650
rect 4988 12640 5040 12646
rect 4986 12608 4988 12617
rect 5040 12608 5042 12617
rect 4986 12543 5042 12552
rect 4712 12232 4764 12238
rect 4896 12232 4948 12238
rect 4712 12174 4764 12180
rect 4816 12192 4896 12220
rect 4448 11852 4660 11880
rect 4344 11834 4396 11840
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4540 11506 4568 11698
rect 4080 11342 4200 11370
rect 4264 11478 4568 11506
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3620 10742 3648 11222
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 10169 3464 10406
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3422 10160 3478 10169
rect 3422 10095 3478 10104
rect 3606 10160 3662 10169
rect 3606 10095 3608 10104
rect 3660 10095 3662 10104
rect 3608 10066 3660 10072
rect 3792 10056 3844 10062
rect 3422 10024 3478 10033
rect 3792 9998 3844 10004
rect 3422 9959 3478 9968
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3238 9480 3294 9489
rect 3238 9415 3294 9424
rect 3436 9178 3464 9959
rect 3804 9654 3832 9998
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3896 9178 3924 10542
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3988 9110 4016 11086
rect 4080 10554 4108 11342
rect 4264 10606 4292 11478
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4252 10600 4304 10606
rect 4080 10526 4200 10554
rect 4252 10542 4304 10548
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 4080 9042 4108 9998
rect 4172 9178 4200 10526
rect 4356 9722 4384 10610
rect 4448 10062 4476 11290
rect 4540 11218 4568 11478
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4342 9616 4398 9625
rect 4342 9551 4398 9560
rect 4356 9518 4384 9551
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2884 7585 2912 7822
rect 2870 7576 2926 7585
rect 2780 7540 2832 7546
rect 2870 7511 2926 7520
rect 2976 7528 3004 7890
rect 3146 7576 3202 7585
rect 2976 7500 3096 7528
rect 3146 7511 3202 7520
rect 2780 7482 2832 7488
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2884 7290 2912 7414
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2792 7262 2912 7290
rect 2792 7206 2820 7262
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2780 6928 2832 6934
rect 2976 6916 3004 7346
rect 3068 7002 3096 7500
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 2832 6888 3004 6916
rect 2780 6870 2832 6876
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2792 6662 2820 6734
rect 2780 6656 2832 6662
rect 2686 6624 2742 6633
rect 2780 6598 2832 6604
rect 2686 6559 2742 6568
rect 3160 6474 3188 7511
rect 3252 6934 3280 8434
rect 3240 6928 3292 6934
rect 3344 6905 3372 8774
rect 3240 6870 3292 6876
rect 3330 6896 3386 6905
rect 3330 6831 3386 6840
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 2700 6446 3188 6474
rect 3252 6458 3280 6598
rect 3240 6452 3292 6458
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 2608 5778 2636 6326
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2332 5324 2452 5352
rect 2228 5160 2280 5166
rect 2226 5128 2228 5137
rect 2280 5128 2282 5137
rect 2226 5063 2282 5072
rect 2240 4185 2268 5063
rect 2226 4176 2282 4185
rect 2226 4111 2282 4120
rect 2332 3670 2360 5324
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2424 5137 2452 5170
rect 2410 5128 2466 5137
rect 2410 5063 2466 5072
rect 2608 4826 2636 5170
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2410 4584 2466 4593
rect 2410 4519 2466 4528
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 2424 3194 2452 4519
rect 2502 4448 2558 4457
rect 2502 4383 2558 4392
rect 2516 3534 2544 4383
rect 2608 3602 2636 4762
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2594 3496 2650 3505
rect 2594 3431 2650 3440
rect 2502 3224 2558 3233
rect 2412 3188 2464 3194
rect 2502 3159 2558 3168
rect 2412 3130 2464 3136
rect 2516 3058 2544 3159
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2226 2544 2282 2553
rect 1952 2508 2004 2514
rect 2226 2479 2282 2488
rect 1952 2450 2004 2456
rect 2240 800 2268 2479
rect 2608 800 2636 3431
rect 2700 3194 2728 6446
rect 3240 6394 3292 6400
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2792 4282 2820 5510
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2884 4010 2912 6258
rect 2976 4078 3004 6326
rect 3344 6322 3372 6598
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5846 3188 6054
rect 3148 5840 3200 5846
rect 3148 5782 3200 5788
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 3068 5370 3096 5578
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3160 4706 3188 5646
rect 3252 5030 3280 6190
rect 3436 5896 3464 8910
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3620 7410 3648 7890
rect 3896 7750 3924 8366
rect 4068 8288 4120 8294
rect 3974 8256 4030 8265
rect 4068 8230 4120 8236
rect 3974 8191 4030 8200
rect 3988 7886 4016 8191
rect 4080 7886 4108 8230
rect 4172 7954 4200 9114
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3712 7449 3740 7686
rect 3698 7440 3754 7449
rect 3608 7404 3660 7410
rect 3698 7375 3754 7384
rect 3608 7346 3660 7352
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3514 6896 3570 6905
rect 3514 6831 3570 6840
rect 3700 6860 3752 6866
rect 3528 6730 3556 6831
rect 3700 6802 3752 6808
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3528 6361 3556 6666
rect 3712 6390 3740 6802
rect 3700 6384 3752 6390
rect 3514 6352 3570 6361
rect 3700 6326 3752 6332
rect 3514 6287 3570 6296
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3516 5908 3568 5914
rect 3436 5868 3516 5896
rect 3516 5850 3568 5856
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3344 4826 3372 5782
rect 3792 5704 3844 5710
rect 3790 5672 3792 5681
rect 3844 5672 3846 5681
rect 3790 5607 3846 5616
rect 3792 5568 3844 5574
rect 3514 5536 3570 5545
rect 3792 5510 3844 5516
rect 3514 5471 3570 5480
rect 3424 5296 3476 5302
rect 3422 5264 3424 5273
rect 3476 5264 3478 5273
rect 3422 5199 3478 5208
rect 3528 5148 3556 5471
rect 3436 5120 3556 5148
rect 3804 5137 3832 5510
rect 3896 5302 3924 7686
rect 4264 7546 4292 9454
rect 4344 9376 4396 9382
rect 4448 9364 4476 9862
rect 4540 9586 4568 11018
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4396 9336 4476 9364
rect 4344 9318 4396 9324
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4264 7410 4292 7482
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 3974 7168 4030 7177
rect 3974 7103 4030 7112
rect 3988 6934 4016 7103
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 4080 6798 4108 7346
rect 4356 7206 4384 9318
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4448 7274 4476 7346
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4342 7032 4398 7041
rect 4342 6967 4398 6976
rect 4250 6896 4306 6905
rect 4250 6831 4306 6840
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4080 5658 4108 6326
rect 4172 6322 4200 6598
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4264 5817 4292 6831
rect 4356 6798 4384 6967
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4250 5808 4306 5817
rect 4250 5743 4306 5752
rect 3988 5630 4108 5658
rect 4160 5704 4212 5710
rect 4356 5658 4384 6598
rect 4448 5778 4476 7210
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4160 5646 4212 5652
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3884 5160 3936 5166
rect 3790 5128 3846 5137
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3160 4678 3372 4706
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 3068 4282 3096 4490
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 3068 3602 3096 4218
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3160 3482 3188 4150
rect 3344 4010 3372 4678
rect 3436 4321 3464 5120
rect 3884 5102 3936 5108
rect 3790 5063 3846 5072
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3896 4690 3924 5102
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3792 4616 3844 4622
rect 3988 4570 4016 5630
rect 4172 5556 4200 5646
rect 4264 5642 4384 5658
rect 4252 5636 4384 5642
rect 4304 5630 4384 5636
rect 4252 5578 4304 5584
rect 3792 4558 3844 4564
rect 3620 4486 3648 4558
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3422 4312 3478 4321
rect 3422 4247 3478 4256
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3804 3924 3832 4558
rect 3896 4542 4016 4570
rect 4080 5528 4200 5556
rect 3896 4282 3924 4542
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3330 3904 3386 3913
rect 3804 3896 3924 3924
rect 3330 3839 3386 3848
rect 2976 3454 3188 3482
rect 3344 3482 3372 3839
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3516 3596 3568 3602
rect 3896 3584 3924 3896
rect 3516 3538 3568 3544
rect 3804 3556 3924 3584
rect 3344 3454 3464 3482
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2688 2984 2740 2990
rect 2740 2932 2912 2938
rect 2688 2926 2912 2932
rect 2700 2910 2912 2926
rect 2884 2689 2912 2910
rect 2870 2680 2926 2689
rect 2870 2615 2926 2624
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2792 1193 2820 2382
rect 2884 1698 2912 2382
rect 2872 1692 2924 1698
rect 2872 1634 2924 1640
rect 2778 1184 2834 1193
rect 2778 1119 2834 1128
rect 2976 800 3004 3454
rect 3240 3392 3292 3398
rect 3146 3360 3202 3369
rect 3240 3334 3292 3340
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3146 3295 3202 3304
rect 3160 3194 3188 3295
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 3160 2650 3188 2790
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3146 2544 3202 2553
rect 3146 2479 3148 2488
rect 3200 2479 3202 2488
rect 3148 2450 3200 2456
rect 3252 2446 3280 3334
rect 3344 3194 3372 3334
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3436 3126 3464 3454
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3528 3058 3556 3538
rect 3804 3097 3832 3556
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 3790 3088 3846 3097
rect 3516 3052 3568 3058
rect 3896 3058 3924 3402
rect 3790 3023 3846 3032
rect 3884 3052 3936 3058
rect 3516 2994 3568 3000
rect 3884 2994 3936 3000
rect 3330 2952 3386 2961
rect 3514 2952 3570 2961
rect 3330 2887 3386 2896
rect 3436 2910 3514 2938
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3344 800 3372 2887
rect 3436 2417 3464 2910
rect 3514 2887 3570 2896
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3422 2408 3478 2417
rect 3422 2343 3478 2352
rect 3516 2372 3568 2378
rect 3516 2314 3568 2320
rect 3528 2038 3556 2314
rect 3712 2281 3740 2450
rect 3698 2272 3754 2281
rect 3698 2207 3754 2216
rect 3516 2032 3568 2038
rect 3516 1974 3568 1980
rect 3712 800 3740 2207
rect 3988 1873 4016 4422
rect 3790 1864 3846 1873
rect 3790 1799 3846 1808
rect 3974 1864 4030 1873
rect 3974 1799 4030 1808
rect 3804 1766 3832 1799
rect 3792 1760 3844 1766
rect 3792 1702 3844 1708
rect 4080 1170 4108 5528
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4172 4554 4200 4966
rect 4264 4729 4292 5238
rect 4342 4856 4398 4865
rect 4342 4791 4398 4800
rect 4436 4820 4488 4826
rect 4250 4720 4306 4729
rect 4250 4655 4306 4664
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4160 3052 4212 3058
rect 4264 3040 4292 4422
rect 4356 3398 4384 4791
rect 4436 4762 4488 4768
rect 4448 4622 4476 4762
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4212 3012 4292 3040
rect 4160 2994 4212 3000
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4356 1834 4384 2382
rect 4344 1828 4396 1834
rect 4344 1770 4396 1776
rect 3896 1142 4108 1170
rect 1596 734 1808 762
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 3896 105 3924 1142
rect 4080 800 4108 1142
rect 4448 800 4476 4558
rect 4540 2961 4568 9522
rect 4632 8566 4660 11852
rect 4816 11830 4844 12192
rect 4896 12174 4948 12180
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4724 7936 4752 11494
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4816 10810 4844 11018
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4802 10296 4858 10305
rect 4802 10231 4858 10240
rect 4816 9450 4844 10231
rect 4908 10146 4936 12038
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5000 10266 5028 11698
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4908 10118 5028 10146
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 4804 8832 4856 8838
rect 4908 8809 4936 9454
rect 4804 8774 4856 8780
rect 4894 8800 4950 8809
rect 4816 8498 4844 8774
rect 4894 8735 4950 8744
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4632 7908 4752 7936
rect 4632 5030 4660 7908
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4724 7546 4752 7754
rect 4816 7721 4844 8298
rect 4908 8090 4936 8570
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4802 7712 4858 7721
rect 4802 7647 4858 7656
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4712 7404 4764 7410
rect 4816 7392 4844 7647
rect 4764 7364 4844 7392
rect 4896 7404 4948 7410
rect 4712 7346 4764 7352
rect 4896 7346 4948 7352
rect 4712 7200 4764 7206
rect 4764 7148 4844 7154
rect 4712 7142 4844 7148
rect 4724 7126 4844 7142
rect 4712 6656 4764 6662
rect 4710 6624 4712 6633
rect 4764 6624 4766 6633
rect 4710 6559 4766 6568
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4724 5710 4752 6190
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4724 5098 4752 5646
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4816 4729 4844 7126
rect 4908 6100 4936 7346
rect 5000 6769 5028 10118
rect 5092 10033 5120 13688
rect 5184 11121 5212 13926
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5276 13190 5304 13806
rect 5368 13802 5396 14758
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5460 13394 5488 14214
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5552 13258 5580 15030
rect 5920 15026 5948 15127
rect 5722 14991 5778 15000
rect 5816 15020 5868 15026
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5644 14414 5672 14894
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5644 14074 5672 14350
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5264 13184 5316 13190
rect 5448 13184 5500 13190
rect 5264 13126 5316 13132
rect 5446 13152 5448 13161
rect 5500 13152 5502 13161
rect 5446 13087 5502 13096
rect 5644 12918 5672 13262
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5736 12850 5764 14991
rect 5816 14962 5868 14968
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5828 13734 5856 14962
rect 6012 14822 6040 15302
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6564 15162 6592 15302
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6460 14884 6512 14890
rect 6460 14826 6512 14832
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6472 14414 6500 14826
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5920 12850 5948 13942
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6184 13796 6236 13802
rect 6184 13738 6236 13744
rect 6104 13530 6132 13738
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 5356 12844 5408 12850
rect 5540 12844 5592 12850
rect 5356 12786 5408 12792
rect 5460 12804 5540 12832
rect 5368 12646 5396 12786
rect 5356 12640 5408 12646
rect 5276 12600 5356 12628
rect 5276 12073 5304 12600
rect 5356 12582 5408 12588
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5262 12064 5318 12073
rect 5262 11999 5318 12008
rect 5368 11898 5396 12106
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5170 11112 5226 11121
rect 5170 11047 5226 11056
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5184 10130 5212 10746
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5078 10024 5134 10033
rect 5078 9959 5134 9968
rect 5276 9674 5304 11290
rect 5460 10826 5488 12804
rect 5540 12786 5592 12792
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 6012 12782 6040 13194
rect 6196 13190 6224 13738
rect 6564 13705 6592 14826
rect 6656 13802 6684 15535
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6550 13696 6606 13705
rect 6550 13631 6606 13640
rect 6564 13326 6592 13631
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6552 13184 6604 13190
rect 6656 13161 6684 13194
rect 6552 13126 6604 13132
rect 6642 13152 6698 13161
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 5644 12434 5672 12718
rect 5644 12406 5764 12434
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5368 10798 5488 10826
rect 5368 10674 5396 10798
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5368 9722 5396 10610
rect 5552 10266 5580 11766
rect 5644 11694 5672 12038
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5644 11286 5672 11630
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5460 9994 5488 10066
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5092 9646 5304 9674
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5092 7857 5120 9646
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5184 9110 5212 9454
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5172 8968 5224 8974
rect 5264 8968 5316 8974
rect 5172 8910 5224 8916
rect 5262 8936 5264 8945
rect 5316 8936 5318 8945
rect 5184 8634 5212 8910
rect 5262 8871 5318 8880
rect 5262 8800 5318 8809
rect 5262 8735 5318 8744
rect 5276 8634 5304 8735
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7886 5212 8230
rect 5368 8022 5396 8978
rect 5460 8430 5488 9930
rect 5540 9920 5592 9926
rect 5538 9888 5540 9897
rect 5592 9888 5594 9897
rect 5538 9823 5594 9832
rect 5552 9654 5580 9823
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5538 9072 5594 9081
rect 5538 9007 5594 9016
rect 5552 8838 5580 9007
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5538 8528 5594 8537
rect 5538 8463 5594 8472
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5172 7880 5224 7886
rect 5078 7848 5134 7857
rect 5172 7822 5224 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5078 7783 5134 7792
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4986 6760 5042 6769
rect 4986 6695 5042 6704
rect 4986 6624 5042 6633
rect 4986 6559 5042 6568
rect 5000 6390 5028 6559
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 5092 6118 5120 7686
rect 5184 7206 5212 7822
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5264 6860 5316 6866
rect 5184 6820 5264 6848
rect 4988 6112 5040 6118
rect 4908 6072 4988 6100
rect 4988 6054 5040 6060
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4894 5944 4950 5953
rect 4894 5879 4950 5888
rect 4908 4826 4936 5879
rect 5000 5642 5028 6054
rect 5184 5817 5212 6820
rect 5264 6802 5316 6808
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 5276 6361 5304 6666
rect 5262 6352 5318 6361
rect 5262 6287 5318 6296
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5170 5808 5226 5817
rect 5170 5743 5226 5752
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 5276 5370 5304 6122
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 4988 5296 5040 5302
rect 4988 5238 5040 5244
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4802 4720 4858 4729
rect 4802 4655 4858 4664
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4632 4078 4660 4490
rect 4804 4480 4856 4486
rect 4802 4448 4804 4457
rect 4896 4480 4948 4486
rect 4856 4448 4858 4457
rect 4896 4422 4948 4428
rect 4802 4383 4858 4392
rect 4908 4321 4936 4422
rect 4894 4312 4950 4321
rect 4712 4276 4764 4282
rect 4894 4247 4950 4256
rect 4712 4218 4764 4224
rect 4724 4078 4752 4218
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4724 3670 4752 4014
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4526 2952 4582 2961
rect 4526 2887 4582 2896
rect 4632 1290 4660 3470
rect 4710 2680 4766 2689
rect 4710 2615 4766 2624
rect 4724 2582 4752 2615
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4620 1284 4672 1290
rect 4620 1226 4672 1232
rect 4816 800 4844 3878
rect 4908 2990 4936 4082
rect 5000 3346 5028 5238
rect 5080 5228 5132 5234
rect 5132 5188 5212 5216
rect 5080 5170 5132 5176
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5092 3534 5120 4626
rect 5184 4146 5212 5188
rect 5262 4992 5318 5001
rect 5262 4927 5318 4936
rect 5276 4826 5304 4927
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5262 4720 5318 4729
rect 5262 4655 5318 4664
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5000 3318 5120 3346
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4986 2952 5042 2961
rect 4986 2887 5042 2896
rect 5000 2650 5028 2887
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 5000 1970 5028 2314
rect 4988 1964 5040 1970
rect 4988 1906 5040 1912
rect 5092 1034 5120 3318
rect 5276 2774 5304 4655
rect 5368 2854 5396 7822
rect 5552 7562 5580 8463
rect 5644 7750 5672 11018
rect 5736 7886 5764 12406
rect 6196 12084 6224 12854
rect 6380 12646 6408 12922
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6288 12424 6316 12582
rect 6368 12436 6420 12442
rect 6288 12396 6368 12424
rect 6368 12378 6420 12384
rect 6012 12056 6224 12084
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5828 11354 5856 11698
rect 6012 11558 6040 12056
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6366 11792 6422 11801
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5906 11384 5962 11393
rect 5816 11348 5868 11354
rect 5906 11319 5962 11328
rect 6090 11384 6146 11393
rect 6090 11319 6146 11328
rect 5816 11290 5868 11296
rect 5920 11121 5948 11319
rect 6104 11218 6132 11319
rect 6092 11212 6144 11218
rect 6012 11172 6092 11200
rect 5906 11112 5962 11121
rect 5906 11047 5962 11056
rect 6012 10713 6040 11172
rect 6092 11154 6144 11160
rect 6196 11014 6224 11766
rect 6366 11727 6422 11736
rect 6380 11218 6408 11727
rect 6564 11336 6592 13126
rect 6642 13087 6698 13096
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6656 12374 6684 12786
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6748 12186 6776 16510
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6840 16250 6868 16390
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 14890 6868 15846
rect 6932 15706 6960 19722
rect 7024 19281 7052 20295
rect 7116 19718 7144 20334
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7102 19544 7158 19553
rect 7208 19514 7236 19654
rect 7102 19479 7158 19488
rect 7196 19508 7248 19514
rect 7116 19360 7144 19479
rect 7196 19450 7248 19456
rect 7196 19372 7248 19378
rect 7116 19332 7196 19360
rect 7300 19352 7328 20470
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 7392 19718 7420 20402
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7196 19314 7248 19320
rect 7288 19346 7340 19352
rect 7288 19288 7340 19294
rect 7010 19272 7066 19281
rect 7392 19258 7420 19654
rect 7116 19242 7420 19258
rect 7010 19207 7066 19216
rect 7104 19236 7420 19242
rect 7156 19230 7420 19236
rect 7104 19178 7156 19184
rect 7378 19136 7434 19145
rect 7378 19071 7434 19080
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 7024 18290 7052 18634
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7024 17610 7052 18226
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 17134 7144 17478
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7208 16794 7236 18226
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7024 16182 7052 16390
rect 7012 16176 7064 16182
rect 7012 16118 7064 16124
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6932 14618 6960 15302
rect 7024 15162 7052 15302
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6840 14006 6868 14554
rect 6918 14512 6974 14521
rect 6918 14447 6974 14456
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6932 13870 6960 14447
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 7024 13546 7052 14826
rect 7116 14278 7144 15506
rect 7208 14958 7236 16390
rect 7300 15144 7328 18362
rect 7392 16454 7420 19071
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7380 15156 7432 15162
rect 7300 15116 7380 15144
rect 7380 15098 7432 15104
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7286 14512 7342 14521
rect 7286 14447 7342 14456
rect 7300 14414 7328 14447
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 6656 12158 6776 12186
rect 6840 13518 7052 13546
rect 6656 11506 6684 12158
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11626 6776 12038
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6656 11478 6776 11506
rect 6564 11308 6684 11336
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6380 11082 6408 11154
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6564 10810 6592 11018
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 5998 10704 6054 10713
rect 5998 10639 6054 10648
rect 6182 10704 6238 10713
rect 6182 10639 6238 10648
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5828 9586 5856 9862
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 8090 5856 9522
rect 5920 9518 5948 10542
rect 6196 10538 6224 10639
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6460 10532 6512 10538
rect 6460 10474 6512 10480
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6368 10464 6420 10470
rect 6472 10441 6500 10474
rect 6368 10406 6420 10412
rect 6458 10432 6514 10441
rect 5908 9512 5960 9518
rect 5906 9480 5908 9489
rect 5960 9480 5962 9489
rect 5906 9415 5962 9424
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5814 7848 5870 7857
rect 5814 7783 5870 7792
rect 5828 7750 5856 7783
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5552 7534 5856 7562
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 4622 5488 7346
rect 5828 7206 5856 7534
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5460 4078 5488 4422
rect 5552 4282 5580 7142
rect 5920 7018 5948 9114
rect 6012 9058 6040 10406
rect 6274 10296 6330 10305
rect 6274 10231 6330 10240
rect 6288 9926 6316 10231
rect 6380 10130 6408 10406
rect 6458 10367 6514 10376
rect 6458 10296 6514 10305
rect 6458 10231 6514 10240
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6472 10010 6500 10231
rect 6564 10130 6592 10746
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6472 9982 6592 10010
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6090 9072 6146 9081
rect 6012 9030 6090 9058
rect 6090 9007 6146 9016
rect 6104 8974 6132 9007
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6196 8820 6224 9658
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6288 9042 6316 9454
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6564 8974 6592 9982
rect 6656 9178 6684 11308
rect 6748 10674 6776 11478
rect 6840 10810 6868 13518
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 7024 12753 7052 13398
rect 7116 13394 7144 14214
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 7010 12744 7066 12753
rect 7010 12679 7066 12688
rect 7102 12336 7158 12345
rect 7102 12271 7104 12280
rect 7156 12271 7158 12280
rect 7104 12242 7156 12248
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6932 11150 6960 12106
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11937 7052 12038
rect 7010 11928 7066 11937
rect 7010 11863 7066 11872
rect 7012 11688 7064 11694
rect 7116 11665 7144 12242
rect 7208 11898 7236 12854
rect 7300 12374 7328 14350
rect 7392 14113 7420 15098
rect 7378 14104 7434 14113
rect 7378 14039 7434 14048
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12986 7420 13126
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7012 11630 7064 11636
rect 7102 11656 7158 11665
rect 7024 11506 7052 11630
rect 7102 11591 7158 11600
rect 7024 11478 7144 11506
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 7024 11014 7052 11222
rect 7116 11218 7144 11478
rect 7300 11234 7328 12310
rect 7392 11393 7420 12378
rect 7378 11384 7434 11393
rect 7484 11354 7512 20470
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7576 19174 7604 19314
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7576 18970 7604 19110
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7576 18222 7604 18906
rect 7564 18216 7616 18222
rect 7668 18193 7696 20402
rect 7852 20233 7880 22222
rect 7930 22200 7986 23000
rect 8298 22200 8354 23000
rect 8666 22200 8722 23000
rect 9034 22200 9090 23000
rect 9140 22222 9352 22250
rect 7838 20224 7894 20233
rect 7838 20159 7894 20168
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7760 18834 7788 19858
rect 7852 18986 7880 20159
rect 7944 19145 7972 22200
rect 8208 20460 8260 20466
rect 8312 20448 8340 22200
rect 8260 20420 8340 20448
rect 8208 20402 8260 20408
rect 8312 19802 8340 20420
rect 8680 20398 8708 22200
rect 9048 22114 9076 22200
rect 9140 22114 9168 22222
rect 9048 22086 9168 22114
rect 9324 20466 9352 22222
rect 9402 22200 9458 23000
rect 9770 22200 9826 23000
rect 10138 22200 10194 23000
rect 10506 22200 10562 23000
rect 10874 22200 10930 23000
rect 11242 22200 11298 23000
rect 11610 22200 11666 23000
rect 11978 22200 12034 23000
rect 12346 22200 12402 23000
rect 12714 22200 12770 23000
rect 13082 22200 13138 23000
rect 13450 22200 13506 23000
rect 13818 22200 13874 23000
rect 14186 22200 14242 23000
rect 14554 22200 14610 23000
rect 14922 22200 14978 23000
rect 15290 22200 15346 23000
rect 15658 22200 15714 23000
rect 16026 22200 16082 23000
rect 16132 22222 16344 22250
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8404 19990 8432 20198
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8208 19780 8260 19786
rect 8312 19774 8432 19802
rect 8208 19722 8260 19728
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 7930 19136 7986 19145
rect 7930 19071 7986 19080
rect 7852 18958 8064 18986
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7564 18158 7616 18164
rect 7654 18184 7710 18193
rect 7654 18119 7710 18128
rect 7760 18086 7788 18770
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 7944 18426 7972 18566
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7656 17264 7708 17270
rect 7654 17232 7656 17241
rect 7708 17232 7710 17241
rect 7564 17196 7616 17202
rect 7654 17167 7710 17176
rect 7564 17138 7616 17144
rect 7576 16833 7604 17138
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7562 16824 7618 16833
rect 7562 16759 7618 16768
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7576 16561 7604 16594
rect 7668 16590 7696 17070
rect 7760 16794 7788 17818
rect 7852 17513 7880 18226
rect 7944 17542 7972 18226
rect 7932 17536 7984 17542
rect 7838 17504 7894 17513
rect 7932 17478 7984 17484
rect 7838 17439 7894 17448
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7852 16998 7880 17138
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7746 16688 7802 16697
rect 7746 16623 7802 16632
rect 7656 16584 7708 16590
rect 7562 16552 7618 16561
rect 7656 16526 7708 16532
rect 7562 16487 7618 16496
rect 7668 16046 7696 16526
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7760 15910 7788 16623
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7852 15745 7880 16934
rect 7838 15736 7894 15745
rect 7748 15700 7800 15706
rect 7838 15671 7894 15680
rect 7748 15642 7800 15648
rect 7760 15162 7788 15642
rect 7944 15586 7972 17478
rect 8036 16250 8064 18958
rect 8128 18306 8156 19654
rect 8220 18426 8248 19722
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8312 19553 8340 19654
rect 8298 19544 8354 19553
rect 8298 19479 8354 19488
rect 8300 18760 8352 18766
rect 8404 18748 8432 19774
rect 8352 18720 8432 18748
rect 8300 18702 8352 18708
rect 8300 18624 8352 18630
rect 8352 18584 8432 18612
rect 8300 18566 8352 18572
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8128 18278 8248 18306
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8128 17270 8156 17682
rect 8220 17649 8248 18278
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8312 17746 8340 18158
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8206 17640 8262 17649
rect 8404 17626 8432 18584
rect 8206 17575 8262 17584
rect 8312 17598 8432 17626
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8220 17338 8248 17478
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 8312 17066 8340 17598
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8404 16794 8432 17478
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8024 16244 8076 16250
rect 8024 16186 8076 16192
rect 8022 16008 8078 16017
rect 8022 15943 8024 15952
rect 8076 15943 8078 15952
rect 8024 15914 8076 15920
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 7944 15558 8064 15586
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7576 14414 7604 14894
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7852 14278 7880 14758
rect 7944 14414 7972 15438
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7852 13734 7880 14010
rect 7944 13938 7972 14350
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 8036 13025 8064 15558
rect 8220 15502 8248 15846
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8116 15360 8168 15366
rect 8312 15337 8340 16390
rect 8116 15302 8168 15308
rect 8298 15328 8354 15337
rect 8128 13938 8156 15302
rect 8298 15263 8354 15272
rect 8496 15162 8524 20198
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8576 19984 8628 19990
rect 8576 19926 8628 19932
rect 8588 18306 8616 19926
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8680 19514 8708 19858
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8772 19514 8800 19654
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8680 18834 8708 19450
rect 8864 19378 8892 19654
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8588 18278 8708 18306
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8588 17338 8616 18158
rect 8576 17332 8628 17338
rect 8680 17320 8708 18278
rect 9048 18154 9076 18566
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 8760 17536 8812 17542
rect 8758 17504 8760 17513
rect 8812 17504 8814 17513
rect 8758 17439 8814 17448
rect 8680 17292 8800 17320
rect 8576 17274 8628 17280
rect 8666 17232 8722 17241
rect 8666 17167 8668 17176
rect 8720 17167 8722 17176
rect 8668 17138 8720 17144
rect 8772 16980 8800 17292
rect 8574 16960 8630 16969
rect 8574 16895 8630 16904
rect 8680 16952 8800 16980
rect 8588 16658 8616 16895
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 8588 15881 8616 16390
rect 8574 15872 8630 15881
rect 8574 15807 8630 15816
rect 8680 15706 8708 16952
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 9048 16182 9076 16594
rect 9140 16250 9168 20334
rect 9416 18766 9444 22200
rect 9784 20482 9812 22200
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9600 20454 9812 20482
rect 9600 19786 9628 20454
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9600 19258 9628 19722
rect 9692 19553 9720 20334
rect 9678 19544 9734 19553
rect 9678 19479 9734 19488
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9600 19230 9720 19258
rect 9692 19174 9720 19230
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9784 18970 9812 19314
rect 10060 19145 10088 20742
rect 10152 20584 10180 22200
rect 10152 20556 10272 20584
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10046 19136 10102 19145
rect 10046 19071 10102 19080
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9494 18864 9550 18873
rect 9494 18799 9550 18808
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9218 17912 9274 17921
rect 9324 17882 9352 18566
rect 9416 18426 9444 18702
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9508 18290 9536 18799
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9588 18216 9640 18222
rect 9416 18164 9588 18170
rect 9640 18164 9720 18170
rect 9416 18142 9720 18164
rect 9218 17847 9274 17856
rect 9312 17876 9364 17882
rect 9232 17649 9260 17847
rect 9312 17818 9364 17824
rect 9218 17640 9274 17649
rect 9218 17575 9274 17584
rect 9416 17320 9444 18142
rect 9692 18086 9720 18142
rect 9680 18080 9732 18086
rect 9784 18057 9812 18634
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9680 18022 9732 18028
rect 9770 18048 9826 18057
rect 9770 17983 9826 17992
rect 9876 17746 9904 18090
rect 10152 17882 10180 20402
rect 10244 19446 10272 20556
rect 10520 20466 10548 22200
rect 10888 20602 10916 22200
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10612 20058 10640 20402
rect 11072 20369 11100 21082
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11058 20360 11114 20369
rect 10968 20324 11020 20330
rect 11058 20295 11114 20304
rect 10968 20266 11020 20272
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10232 19440 10284 19446
rect 10232 19382 10284 19388
rect 10244 18970 10272 19382
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10336 18850 10364 19790
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10876 19780 10928 19786
rect 10876 19722 10928 19728
rect 10428 19310 10456 19722
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10506 19000 10562 19009
rect 10506 18935 10562 18944
rect 10336 18822 10456 18850
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9864 17740 9916 17746
rect 10048 17740 10100 17746
rect 9864 17682 9916 17688
rect 9968 17700 10048 17728
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9232 17292 9444 17320
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8680 15434 8708 15642
rect 9232 15552 9260 17292
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9416 16658 9444 17138
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9324 16250 9352 16390
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9140 15524 9260 15552
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 9140 15337 9168 15524
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9126 15328 9182 15337
rect 9126 15263 9182 15272
rect 8666 15192 8722 15201
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8576 15156 8628 15162
rect 8666 15127 8722 15136
rect 8576 15098 8628 15104
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8220 14657 8248 14962
rect 8206 14648 8262 14657
rect 8206 14583 8262 14592
rect 8312 14414 8340 15098
rect 8588 14618 8616 15098
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8300 14408 8352 14414
rect 8352 14368 8432 14396
rect 8300 14350 8352 14356
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8404 13870 8432 14368
rect 8392 13864 8444 13870
rect 8298 13832 8354 13841
rect 8392 13806 8444 13812
rect 8298 13767 8354 13776
rect 8116 13184 8168 13190
rect 8312 13161 8340 13767
rect 8116 13126 8168 13132
rect 8298 13152 8354 13161
rect 8022 13016 8078 13025
rect 8022 12951 8078 12960
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 8024 12912 8076 12918
rect 8024 12854 8076 12860
rect 7668 12238 7696 12854
rect 8036 12753 8064 12854
rect 8022 12744 8078 12753
rect 8022 12679 8078 12688
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7746 12336 7802 12345
rect 7746 12271 7748 12280
rect 7800 12271 7802 12280
rect 7748 12242 7800 12248
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7760 11898 7788 12242
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7668 11665 7696 11766
rect 7654 11656 7710 11665
rect 7654 11591 7710 11600
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7378 11319 7434 11328
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7104 11212 7156 11218
rect 7300 11206 7420 11234
rect 7104 11154 7156 11160
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7392 10826 7420 11206
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 7300 10798 7420 10826
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6748 9976 6776 10610
rect 6840 10470 6868 10746
rect 7102 10704 7158 10713
rect 7012 10668 7064 10674
rect 6932 10628 7012 10656
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6932 10305 6960 10628
rect 7300 10674 7328 10798
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7102 10639 7158 10648
rect 7288 10668 7340 10674
rect 7012 10610 7064 10616
rect 7116 10470 7144 10639
rect 7288 10610 7340 10616
rect 7104 10464 7156 10470
rect 7010 10432 7066 10441
rect 7104 10406 7156 10412
rect 7194 10432 7250 10441
rect 7010 10367 7066 10376
rect 6918 10296 6974 10305
rect 6918 10231 6974 10240
rect 6828 10056 6880 10062
rect 6880 10016 6960 10044
rect 6828 9998 6880 10004
rect 6739 9948 6776 9976
rect 6739 9908 6767 9948
rect 6739 9880 6776 9908
rect 6644 9172 6696 9178
rect 6748 9160 6776 9880
rect 6826 9752 6882 9761
rect 6826 9687 6882 9696
rect 6840 9586 6868 9687
rect 6932 9586 6960 10016
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6748 9132 6868 9160
rect 6644 9114 6696 9120
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6012 8792 6224 8820
rect 6012 8566 6040 8792
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6550 8664 6606 8673
rect 6276 8628 6328 8634
rect 6328 8608 6550 8616
rect 6656 8634 6684 8978
rect 6328 8599 6606 8608
rect 6644 8628 6696 8634
rect 6328 8588 6592 8599
rect 6276 8570 6328 8576
rect 6644 8570 6696 8576
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 6748 8498 6776 8978
rect 6840 8838 6868 9132
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6090 8120 6146 8129
rect 6090 8055 6092 8064
rect 6144 8055 6146 8064
rect 6092 8026 6144 8032
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6564 7342 6592 8366
rect 6748 7546 6776 8434
rect 6840 7954 6868 8774
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 7024 7834 7052 10367
rect 7116 10198 7144 10406
rect 7194 10367 7250 10376
rect 7208 10266 7236 10367
rect 7392 10305 7420 10678
rect 7378 10296 7434 10305
rect 7196 10260 7248 10266
rect 7378 10231 7434 10240
rect 7196 10202 7248 10208
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7116 9722 7144 10134
rect 7380 9920 7432 9926
rect 7300 9880 7380 9908
rect 7104 9716 7156 9722
rect 7156 9676 7236 9704
rect 7104 9658 7156 9664
rect 7102 8528 7158 8537
rect 7102 8463 7158 8472
rect 7116 7886 7144 8463
rect 6932 7806 7052 7834
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6932 7426 6960 7806
rect 7012 7744 7064 7750
rect 7208 7732 7236 9676
rect 7300 8634 7328 9880
rect 7380 9862 7432 9868
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7392 9178 7420 9454
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7484 8974 7512 11290
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7576 10810 7604 11018
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7668 10538 7696 10950
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7656 10532 7708 10538
rect 7656 10474 7708 10480
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7576 9382 7604 9998
rect 7760 9722 7788 10746
rect 7852 10674 7880 11494
rect 7944 10810 7972 12378
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11937 8064 12038
rect 8022 11928 8078 11937
rect 8022 11863 8078 11872
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 8036 10674 8064 11698
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7838 10296 7894 10305
rect 7838 10231 7894 10240
rect 7852 9994 7880 10231
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7472 8968 7524 8974
rect 7392 8928 7472 8956
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7392 8090 7420 8928
rect 7472 8910 7524 8916
rect 7470 8528 7526 8537
rect 7470 8463 7526 8472
rect 7484 8294 7512 8463
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7012 7686 7064 7692
rect 7116 7704 7236 7732
rect 6748 7398 6960 7426
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 5644 6990 5948 7018
rect 5644 6474 5672 6990
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6633 5764 6734
rect 5722 6624 5778 6633
rect 5722 6559 5778 6568
rect 5644 6446 5764 6474
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5644 5778 5672 6190
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5644 5166 5672 5714
rect 5736 5710 5764 6446
rect 5828 5914 5856 6802
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5920 5914 5948 6598
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5736 5545 5764 5646
rect 5722 5536 5778 5545
rect 5828 5522 5856 5850
rect 6012 5846 6040 6598
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6564 6458 6592 6870
rect 6748 6780 6776 7398
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 7002 6960 7142
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6840 6882 6868 6938
rect 6840 6854 6960 6882
rect 6748 6752 6868 6780
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 6366 6352 6422 6361
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 6104 5692 6132 6258
rect 6196 6089 6224 6258
rect 6182 6080 6238 6089
rect 6182 6015 6238 6024
rect 6012 5664 6132 5692
rect 5828 5494 5948 5522
rect 5722 5471 5778 5480
rect 5814 5400 5870 5409
rect 5724 5364 5776 5370
rect 5814 5335 5816 5344
rect 5724 5306 5776 5312
rect 5868 5335 5870 5344
rect 5816 5306 5868 5312
rect 5736 5216 5764 5306
rect 5736 5188 5856 5216
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5552 3924 5580 4082
rect 5460 3896 5580 3924
rect 5460 3534 5488 3896
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5552 3398 5580 3674
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5184 2746 5304 2774
rect 5184 2446 5212 2746
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5276 2360 5304 2518
rect 5460 2514 5488 3334
rect 5538 3224 5594 3233
rect 5538 3159 5594 3168
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5356 2372 5408 2378
rect 5276 2332 5356 2360
rect 5356 2314 5408 2320
rect 5092 1006 5212 1034
rect 5184 800 5212 1006
rect 5552 800 5580 3159
rect 5644 2394 5672 4966
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5736 4593 5764 4694
rect 5828 4690 5856 5188
rect 5920 4690 5948 5494
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5722 4584 5778 4593
rect 6012 4570 6040 5664
rect 6288 5574 6316 6326
rect 6472 6338 6500 6394
rect 6550 6352 6606 6361
rect 6472 6310 6550 6338
rect 6366 6287 6422 6296
rect 6550 6287 6606 6296
rect 6380 5681 6408 6287
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6472 5710 6500 5850
rect 6460 5704 6512 5710
rect 6366 5672 6422 5681
rect 6460 5646 6512 5652
rect 6366 5607 6422 5616
rect 6380 5574 6408 5607
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6104 4729 6132 5170
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6090 4720 6146 4729
rect 6196 4690 6224 4966
rect 6288 4758 6316 5170
rect 6460 5160 6512 5166
rect 6458 5128 6460 5137
rect 6512 5128 6514 5137
rect 6458 5063 6514 5072
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6090 4655 6146 4664
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 5722 4519 5778 4528
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5920 4542 6040 4570
rect 6092 4616 6144 4622
rect 6380 4570 6408 4966
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6144 4564 6408 4570
rect 6092 4558 6408 4564
rect 6104 4542 6408 4558
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5736 3194 5764 3878
rect 5828 3194 5856 4490
rect 5920 4282 5948 4542
rect 6472 4468 6500 4626
rect 6012 4440 6500 4468
rect 5908 4276 5960 4282
rect 6012 4264 6040 4440
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6012 4236 6224 4264
rect 5908 4218 5960 4224
rect 6196 4078 6224 4236
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6012 3754 6040 4014
rect 5908 3732 5960 3738
rect 6012 3726 6132 3754
rect 5908 3674 5960 3680
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5920 2990 5948 3674
rect 6104 3505 6132 3726
rect 6090 3496 6146 3505
rect 6000 3460 6052 3466
rect 6196 3466 6224 4014
rect 6288 3777 6316 4150
rect 6368 4072 6420 4078
rect 6366 4040 6368 4049
rect 6420 4040 6422 4049
rect 6366 3975 6422 3984
rect 6274 3768 6330 3777
rect 6274 3703 6330 3712
rect 6472 3641 6500 4150
rect 6458 3632 6514 3641
rect 6458 3567 6514 3576
rect 6564 3534 6592 6054
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6090 3431 6146 3440
rect 6184 3460 6236 3466
rect 6000 3402 6052 3408
rect 6184 3402 6236 3408
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 5644 2366 5764 2394
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 5644 1902 5672 2246
rect 5632 1896 5684 1902
rect 5632 1838 5684 1844
rect 5736 1306 5764 2366
rect 5828 1426 5856 2858
rect 5920 2514 5948 2926
rect 6012 2854 6040 3402
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6656 2774 6684 6666
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6564 2746 6684 2774
rect 6564 2650 6592 2746
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6564 2106 6592 2450
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 6748 2038 6776 6598
rect 6840 6361 6868 6752
rect 6826 6352 6882 6361
rect 6826 6287 6882 6296
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6840 4826 6868 6190
rect 6932 5760 6960 6854
rect 7024 6390 7052 7686
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6932 5732 7052 5760
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6840 3534 6868 4762
rect 6932 4593 6960 5578
rect 7024 5574 7052 5732
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7024 5370 7052 5510
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6918 4584 6974 4593
rect 6918 4519 6974 4528
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6918 3632 6974 3641
rect 7024 3602 7052 4422
rect 7116 4214 7144 7704
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 6934 7236 7142
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7208 5710 7236 6734
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7300 5556 7328 7958
rect 7378 7712 7434 7721
rect 7378 7647 7434 7656
rect 7392 7410 7420 7647
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7392 7177 7420 7210
rect 7378 7168 7434 7177
rect 7378 7103 7434 7112
rect 7484 6914 7512 7958
rect 7576 7886 7604 8230
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 7546 7604 7686
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7668 7002 7696 9522
rect 7760 9178 7788 9658
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8430 7788 8910
rect 7852 8809 7880 9590
rect 7944 9586 7972 10406
rect 8036 10062 8064 10474
rect 8128 10180 8156 13126
rect 8298 13087 8354 13096
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8206 12608 8262 12617
rect 8206 12543 8262 12552
rect 8220 12374 8248 12543
rect 8312 12442 8340 12922
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11014 8248 12038
rect 8312 11150 8340 12106
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8404 10810 8432 13806
rect 8496 12782 8524 14418
rect 8680 13734 8708 15127
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 9140 14890 9168 15030
rect 9232 14958 9260 15370
rect 9324 15314 9352 16050
rect 9404 15360 9456 15366
rect 9324 15308 9404 15314
rect 9324 15302 9456 15308
rect 9324 15286 9444 15302
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9140 14793 9168 14826
rect 9126 14784 9182 14793
rect 8747 14716 9055 14725
rect 9126 14719 9182 14728
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9324 14521 9352 15286
rect 9508 15065 9536 17478
rect 9692 17134 9720 17682
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9692 16794 9720 17070
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9600 15162 9628 16390
rect 9692 16114 9720 16594
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9784 15994 9812 17070
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9692 15966 9812 15994
rect 9692 15910 9720 15966
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9692 15502 9720 15846
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9876 15162 9904 16390
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9494 15056 9550 15065
rect 9494 14991 9550 15000
rect 9680 14952 9732 14958
rect 9416 14900 9680 14906
rect 9416 14894 9732 14900
rect 9416 14878 9720 14894
rect 9416 14822 9444 14878
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9402 14648 9458 14657
rect 9402 14583 9458 14592
rect 8942 14512 8998 14521
rect 8942 14447 8944 14456
rect 8996 14447 8998 14456
rect 9310 14512 9366 14521
rect 9310 14447 9366 14456
rect 8944 14418 8996 14424
rect 9416 14396 9444 14583
rect 9508 14414 9536 14758
rect 9586 14512 9642 14521
rect 9586 14447 9642 14456
rect 9324 14368 9444 14396
rect 9496 14408 9548 14414
rect 9324 14278 9352 14368
rect 9496 14350 9548 14356
rect 9312 14272 9364 14278
rect 9034 14240 9090 14249
rect 9600 14226 9628 14447
rect 9312 14214 9364 14220
rect 9034 14175 9090 14184
rect 9048 13938 9076 14175
rect 9324 13954 9352 14214
rect 9416 14198 9628 14226
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9416 14074 9444 14198
rect 9770 14104 9826 14113
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9496 14068 9548 14074
rect 9876 14074 9904 14214
rect 9770 14039 9826 14048
rect 9864 14068 9916 14074
rect 9496 14010 9548 14016
rect 9036 13932 9088 13938
rect 9324 13926 9444 13954
rect 9036 13874 9088 13880
rect 8942 13832 8998 13841
rect 8942 13767 8944 13776
rect 8996 13767 8998 13776
rect 8944 13738 8996 13744
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 8574 13560 8630 13569
rect 8574 13495 8576 13504
rect 8628 13495 8630 13504
rect 8576 13466 8628 13472
rect 8680 12986 8708 13670
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 9140 12986 9168 13670
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 8576 12912 8628 12918
rect 8628 12860 8708 12866
rect 8576 12854 8708 12860
rect 8588 12838 8708 12854
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8576 12708 8628 12714
rect 8576 12650 8628 12656
rect 8588 12481 8616 12650
rect 8574 12472 8630 12481
rect 8574 12407 8630 12416
rect 8680 12424 8708 12838
rect 9232 12782 9260 13398
rect 9324 13190 9352 13670
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9218 12608 9274 12617
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8760 12436 8812 12442
rect 8680 12396 8760 12424
rect 8760 12378 8812 12384
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8588 11937 8616 12038
rect 8574 11928 8630 11937
rect 8574 11863 8630 11872
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8496 11082 8524 11562
rect 8574 11384 8630 11393
rect 8680 11370 8708 12038
rect 8864 11558 8892 12174
rect 9034 11928 9090 11937
rect 9034 11863 9036 11872
rect 9088 11863 9090 11872
rect 9036 11834 9088 11840
rect 8944 11824 8996 11830
rect 9140 11778 9168 12582
rect 9218 12543 9274 12552
rect 9232 12374 9260 12543
rect 9220 12368 9272 12374
rect 9220 12310 9272 12316
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 8996 11772 9168 11778
rect 8944 11766 9168 11772
rect 8956 11750 9168 11766
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8630 11342 8708 11370
rect 8760 11348 8812 11354
rect 8574 11319 8630 11328
rect 9140 11336 9168 11750
rect 9232 11336 9260 12174
rect 9312 11824 9364 11830
rect 9312 11766 9364 11772
rect 8760 11290 8812 11296
rect 8956 11308 9168 11336
rect 9223 11308 9260 11336
rect 8772 11257 8800 11290
rect 8574 11248 8630 11257
rect 8574 11183 8630 11192
rect 8758 11248 8814 11257
rect 8758 11183 8814 11192
rect 8588 11150 8616 11183
rect 8956 11150 8984 11308
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9128 11212 9180 11218
rect 9223 11200 9251 11308
rect 9324 11257 9352 11766
rect 9180 11172 9251 11200
rect 9310 11248 9366 11257
rect 9310 11183 9366 11192
rect 9128 11154 9180 11160
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8312 10690 8340 10746
rect 8496 10690 8524 11018
rect 8942 10840 8998 10849
rect 8668 10804 8720 10810
rect 8942 10775 8998 10784
rect 8668 10746 8720 10752
rect 8312 10662 8524 10690
rect 8574 10704 8630 10713
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8128 10152 8248 10180
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7944 9024 7972 9318
rect 7944 8996 8156 9024
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 7838 8800 7894 8809
rect 7838 8735 7894 8744
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7838 8120 7894 8129
rect 7838 8055 7894 8064
rect 7852 7886 7880 8055
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7840 7744 7892 7750
rect 7746 7712 7802 7721
rect 7840 7686 7892 7692
rect 7746 7647 7802 7656
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7392 6886 7512 6914
rect 7760 6905 7788 7647
rect 7852 7342 7880 7686
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7746 6896 7802 6905
rect 7392 6662 7420 6886
rect 7746 6831 7802 6840
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7208 5528 7328 5556
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 6918 3567 6974 3576
rect 7012 3596 7064 3602
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6840 3194 6868 3470
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6644 2032 6696 2038
rect 6644 1974 6696 1980
rect 6736 2032 6788 2038
rect 6736 1974 6788 1980
rect 6656 1737 6684 1974
rect 6642 1728 6698 1737
rect 6642 1663 6698 1672
rect 5816 1420 5868 1426
rect 5816 1362 5868 1368
rect 6276 1420 6328 1426
rect 6276 1362 6328 1368
rect 5736 1278 5948 1306
rect 5920 800 5948 1278
rect 6288 800 6316 1362
rect 6656 800 6684 1663
rect 6932 1442 6960 3567
rect 7012 3538 7064 3544
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 7024 3194 7052 3402
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7208 3126 7236 5528
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7300 5098 7328 5238
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 7286 4856 7342 4865
rect 7286 4791 7342 4800
rect 7300 4554 7328 4791
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7286 4312 7342 4321
rect 7286 4247 7342 4256
rect 7300 3398 7328 4247
rect 7288 3392 7340 3398
rect 7392 3369 7420 6394
rect 7484 6118 7512 6734
rect 7760 6610 7788 6831
rect 7576 6582 7788 6610
rect 7576 6390 7604 6582
rect 7654 6488 7710 6497
rect 7654 6423 7656 6432
rect 7708 6423 7710 6432
rect 7748 6452 7800 6458
rect 7656 6394 7708 6400
rect 7748 6394 7800 6400
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7472 6112 7524 6118
rect 7576 6089 7604 6190
rect 7472 6054 7524 6060
rect 7562 6080 7618 6089
rect 7288 3334 7340 3340
rect 7378 3360 7434 3369
rect 7378 3295 7434 3304
rect 7392 3126 7420 3295
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7484 2972 7512 6054
rect 7562 6015 7618 6024
rect 7668 5545 7696 6394
rect 7654 5536 7710 5545
rect 7654 5471 7710 5480
rect 7562 5400 7618 5409
rect 7562 5335 7564 5344
rect 7616 5335 7618 5344
rect 7564 5306 7616 5312
rect 7760 5234 7788 6394
rect 7852 6254 7880 7278
rect 7944 6361 7972 8842
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 7954 8064 8774
rect 8128 8634 8156 8996
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8220 8548 8248 10152
rect 8312 9217 8340 10542
rect 8404 10130 8432 10662
rect 8574 10639 8630 10648
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8404 9722 8432 9862
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8392 9580 8444 9586
rect 8444 9540 8524 9568
rect 8392 9522 8444 9528
rect 8298 9208 8354 9217
rect 8298 9143 8354 9152
rect 8298 8936 8354 8945
rect 8298 8871 8354 8880
rect 8312 8673 8340 8871
rect 8298 8664 8354 8673
rect 8298 8599 8354 8608
rect 8114 8528 8170 8537
rect 8220 8520 8432 8548
rect 8114 8463 8170 8472
rect 8128 8362 8156 8463
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 7546 8064 7686
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8128 7478 8156 7754
rect 8404 7562 8432 8520
rect 8496 8412 8524 9540
rect 8588 8786 8616 10639
rect 8680 10146 8708 10746
rect 8956 10742 8984 10775
rect 9048 10742 9076 11154
rect 9416 10962 9444 13926
rect 9508 13818 9536 14010
rect 9784 14006 9812 14039
rect 9864 14010 9916 14016
rect 9772 14000 9824 14006
rect 9678 13968 9734 13977
rect 9772 13942 9824 13948
rect 9678 13903 9734 13912
rect 9508 13790 9628 13818
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9508 12986 9536 13262
rect 9600 13258 9628 13790
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9692 12986 9720 13903
rect 9968 13734 9996 17700
rect 10048 17682 10100 17688
rect 10140 17536 10192 17542
rect 10138 17504 10140 17513
rect 10192 17504 10194 17513
rect 10138 17439 10194 17448
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9956 13728 10008 13734
rect 10060 13705 10088 16526
rect 9956 13670 10008 13676
rect 10046 13696 10102 13705
rect 10046 13631 10102 13640
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9494 12472 9550 12481
rect 9494 12407 9496 12416
rect 9548 12407 9550 12416
rect 9496 12378 9548 12384
rect 9784 12374 9812 13262
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9876 12850 9904 12922
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 10060 12782 10088 13194
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9772 12368 9824 12374
rect 9692 12328 9772 12356
rect 9416 10934 9536 10962
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 9312 10736 9364 10742
rect 9364 10696 9444 10724
rect 9312 10678 9364 10684
rect 9218 10432 9274 10441
rect 8747 10364 9055 10373
rect 9218 10367 9274 10376
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 9126 10296 9182 10305
rect 8864 10240 9126 10248
rect 9232 10282 9260 10367
rect 8864 10231 9182 10240
rect 9223 10254 9260 10282
rect 8864 10220 9168 10231
rect 8680 10118 8800 10146
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8680 8974 8708 9998
rect 8772 9364 8800 10118
rect 8864 9994 8892 10220
rect 9223 10180 9251 10254
rect 9416 10198 9444 10696
rect 9404 10192 9456 10198
rect 9223 10152 9260 10180
rect 9036 10056 9088 10062
rect 9232 10033 9260 10152
rect 9404 10134 9456 10140
rect 9508 10044 9536 10934
rect 9692 10690 9720 12328
rect 9864 12368 9916 12374
rect 9772 12310 9824 12316
rect 9862 12336 9864 12345
rect 9916 12336 9918 12345
rect 9862 12271 9918 12280
rect 9864 12096 9916 12102
rect 10048 12096 10100 12102
rect 9916 12056 9996 12084
rect 9864 12038 9916 12044
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9784 10810 9812 11698
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9600 10674 9720 10690
rect 9588 10668 9720 10674
rect 9640 10662 9720 10668
rect 9588 10610 9640 10616
rect 9672 10606 9700 10662
rect 9672 10600 9732 10606
rect 9672 10560 9680 10600
rect 9680 10542 9732 10548
rect 9770 10568 9826 10577
rect 9770 10503 9772 10512
rect 9824 10503 9826 10512
rect 9772 10474 9824 10480
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9770 10160 9826 10169
rect 9036 9998 9088 10004
rect 9218 10024 9274 10033
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 9048 9897 9076 9998
rect 9218 9959 9274 9968
rect 9416 10016 9536 10044
rect 9220 9920 9272 9926
rect 9034 9888 9090 9897
rect 9220 9862 9272 9868
rect 9034 9823 9090 9832
rect 8772 9336 9168 9364
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 9140 9178 9168 9336
rect 9128 9172 9180 9178
rect 8956 9132 9128 9160
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8588 8758 8708 8786
rect 8680 8616 8708 8758
rect 8852 8628 8904 8634
rect 8680 8588 8852 8616
rect 8852 8570 8904 8576
rect 8956 8566 8984 9132
rect 9128 9114 9180 9120
rect 9126 8800 9182 8809
rect 9126 8735 9182 8744
rect 8944 8560 8996 8566
rect 8944 8502 8996 8508
rect 8668 8424 8720 8430
rect 8496 8384 8668 8412
rect 8668 8366 8720 8372
rect 9036 8288 9088 8294
rect 8574 8256 8630 8265
rect 8680 8248 9036 8276
rect 8680 8242 8708 8248
rect 8630 8214 8708 8242
rect 9036 8230 9088 8236
rect 8574 8191 8630 8200
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8574 8120 8630 8129
rect 8747 8123 9055 8132
rect 8574 8055 8630 8064
rect 8588 7936 8616 8055
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 8668 7948 8720 7954
rect 8588 7908 8668 7936
rect 8668 7890 8720 7896
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8404 7534 8616 7562
rect 8116 7472 8168 7478
rect 8392 7472 8444 7478
rect 8116 7414 8168 7420
rect 8303 7432 8392 7460
rect 8303 7324 8331 7432
rect 8392 7414 8444 7420
rect 8303 7296 8340 7324
rect 8024 7268 8076 7274
rect 8076 7228 8248 7256
rect 8024 7210 8076 7216
rect 8114 7032 8170 7041
rect 8114 6967 8170 6976
rect 8022 6896 8078 6905
rect 8022 6831 8078 6840
rect 8036 6730 8064 6831
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 7930 6352 7986 6361
rect 7930 6287 7986 6296
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5846 7880 6054
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 8128 5760 8156 6967
rect 8220 6662 8248 7228
rect 8312 6916 8340 7296
rect 8312 6888 8432 6916
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8404 6458 8432 6888
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8482 6352 8538 6361
rect 8482 6287 8538 6296
rect 8300 6112 8352 6118
rect 8352 6072 8432 6100
rect 8300 6054 8352 6060
rect 7944 5732 8156 5760
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7392 2944 7512 2972
rect 7392 2774 7420 2944
rect 7576 2774 7604 5170
rect 7852 5030 7880 5510
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7668 2972 7696 4966
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7760 3097 7788 4558
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7746 3088 7802 3097
rect 7746 3023 7802 3032
rect 7748 2984 7800 2990
rect 7668 2944 7748 2972
rect 7748 2926 7800 2932
rect 7208 2746 7420 2774
rect 7484 2746 7604 2774
rect 7208 2446 7236 2746
rect 7378 2544 7434 2553
rect 7378 2479 7380 2488
rect 7432 2479 7434 2488
rect 7380 2450 7432 2456
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7378 2000 7434 2009
rect 7378 1935 7380 1944
rect 7432 1935 7434 1944
rect 7380 1906 7432 1912
rect 6932 1414 7052 1442
rect 7024 800 7052 1414
rect 7392 800 7420 1906
rect 3882 96 3938 105
rect 3882 31 3938 40
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7484 762 7512 2746
rect 7562 2544 7618 2553
rect 7562 2479 7618 2488
rect 7576 2446 7604 2479
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7852 2310 7880 3334
rect 7944 3126 7972 5732
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 8036 5012 8064 5238
rect 8128 5137 8156 5578
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8220 5370 8248 5510
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8114 5128 8170 5137
rect 8114 5063 8170 5072
rect 8036 4984 8248 5012
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 7760 1970 7788 2246
rect 7748 1964 7800 1970
rect 7748 1906 7800 1912
rect 7944 1630 7972 3062
rect 8036 2650 8064 4422
rect 8128 4146 8156 4626
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8128 3670 8156 3878
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8128 3126 8156 3606
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 8220 3058 8248 4984
rect 8312 4826 8340 5306
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8312 3738 8340 4218
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8404 3602 8432 6072
rect 8496 5710 8524 6287
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8496 5234 8524 5646
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8482 4992 8538 5001
rect 8482 4927 8538 4936
rect 8496 4604 8524 4927
rect 8588 4758 8616 7534
rect 8680 7478 8708 7686
rect 8864 7478 8892 7754
rect 9048 7546 9076 7958
rect 9140 7886 9168 8735
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9232 7818 9260 9862
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9324 7993 9352 9590
rect 9416 8673 9444 10016
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 8838 9536 9862
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9600 9217 9628 9522
rect 9692 9382 9720 10134
rect 9770 10095 9826 10104
rect 9784 9722 9812 10095
rect 9876 9926 9904 11494
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9586 9208 9642 9217
rect 9586 9143 9588 9152
rect 9640 9143 9642 9152
rect 9588 9114 9640 9120
rect 9600 8974 9628 9114
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9402 8664 9458 8673
rect 9692 8634 9720 8842
rect 9402 8599 9404 8608
rect 9456 8599 9458 8608
rect 9680 8628 9732 8634
rect 9404 8570 9456 8576
rect 9680 8570 9732 8576
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9310 7984 9366 7993
rect 9310 7919 9366 7928
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 9128 7268 9180 7274
rect 8680 7228 9128 7256
rect 8680 6458 8708 7228
rect 9128 7210 9180 7216
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8944 6656 8996 6662
rect 9048 6644 9076 6802
rect 9232 6798 9260 7754
rect 9416 7342 9444 7890
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9416 7206 9444 7278
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9310 7032 9366 7041
rect 9310 6967 9366 6976
rect 9324 6798 9352 6967
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9312 6792 9364 6798
rect 9508 6746 9536 8434
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9600 7834 9628 8298
rect 9692 7954 9720 8570
rect 9784 8106 9812 9522
rect 9862 9344 9918 9353
rect 9862 9279 9918 9288
rect 9876 8906 9904 9279
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9876 8401 9904 8842
rect 9862 8392 9918 8401
rect 9862 8327 9918 8336
rect 9968 8294 9996 12056
rect 10048 12038 10100 12044
rect 10060 11121 10088 12038
rect 10046 11112 10102 11121
rect 10046 11047 10102 11056
rect 10046 10568 10102 10577
rect 10046 10503 10102 10512
rect 10060 9897 10088 10503
rect 10152 10010 10180 17274
rect 10244 17270 10272 17750
rect 10232 17264 10284 17270
rect 10232 17206 10284 17212
rect 10336 16454 10364 18702
rect 10428 17882 10456 18822
rect 10520 18630 10548 18935
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10612 17678 10640 19450
rect 10888 18970 10916 19722
rect 10980 18970 11008 20266
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10704 18630 10732 18702
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10704 18222 10732 18566
rect 10784 18284 10836 18290
rect 10784 18226 10836 18232
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 17338 10732 17478
rect 10796 17338 10824 18226
rect 10876 18216 10928 18222
rect 10928 18176 11008 18204
rect 10876 18158 10928 18164
rect 10876 17536 10928 17542
rect 10874 17504 10876 17513
rect 10928 17504 10930 17513
rect 10874 17439 10930 17448
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10416 16720 10468 16726
rect 10416 16662 10468 16668
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10244 15502 10272 16186
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10428 15201 10456 16662
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10520 15570 10548 16050
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10414 15192 10470 15201
rect 10414 15127 10470 15136
rect 10416 15088 10468 15094
rect 10416 15030 10468 15036
rect 10428 14958 10456 15030
rect 10324 14952 10376 14958
rect 10322 14920 10324 14929
rect 10416 14952 10468 14958
rect 10376 14920 10378 14929
rect 10416 14894 10468 14900
rect 10322 14855 10378 14864
rect 10336 14482 10364 14855
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10336 13977 10364 14214
rect 10322 13968 10378 13977
rect 10232 13932 10284 13938
rect 10322 13903 10378 13912
rect 10232 13874 10284 13880
rect 10244 12345 10272 13874
rect 10428 13870 10456 14894
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10520 14074 10548 14554
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10416 13864 10468 13870
rect 10520 13841 10548 14010
rect 10416 13806 10468 13812
rect 10506 13832 10562 13841
rect 10506 13767 10562 13776
rect 10612 13682 10640 16934
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 14550 10732 16390
rect 10888 16250 10916 16594
rect 10980 16454 11008 18176
rect 11060 18080 11112 18086
rect 11164 18057 11192 20878
rect 11256 20058 11284 22200
rect 11624 20890 11652 22200
rect 11624 20862 11744 20890
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11716 20602 11744 20862
rect 11992 20602 12020 22200
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11980 20596 12032 20602
rect 12360 20584 12388 22200
rect 12728 20602 12756 22200
rect 12990 21448 13046 21457
rect 12990 21383 13046 21392
rect 12440 20596 12492 20602
rect 12360 20556 12440 20584
rect 11980 20538 12032 20544
rect 12440 20538 12492 20544
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 11900 19854 11928 20198
rect 12084 20058 12112 20402
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 11612 19848 11664 19854
rect 11610 19816 11612 19825
rect 11888 19848 11940 19854
rect 11664 19816 11666 19825
rect 11888 19790 11940 19796
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 11610 19751 11666 19760
rect 11796 19712 11848 19718
rect 11794 19680 11796 19689
rect 11848 19680 11850 19689
rect 11346 19612 11654 19621
rect 11794 19615 11850 19624
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11612 19372 11664 19378
rect 11808 19334 11836 19615
rect 11612 19314 11664 19320
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11060 18022 11112 18028
rect 11150 18048 11206 18057
rect 11072 17882 11100 18022
rect 11150 17983 11206 17992
rect 11060 17876 11112 17882
rect 11256 17864 11284 19110
rect 11624 18698 11652 19314
rect 11716 19306 11836 19334
rect 11612 18692 11664 18698
rect 11612 18634 11664 18640
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11612 18284 11664 18290
rect 11060 17818 11112 17824
rect 11164 17836 11284 17864
rect 11532 18244 11612 18272
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10796 14958 10824 15642
rect 10888 15434 10916 16186
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10692 14544 10744 14550
rect 10692 14486 10744 14492
rect 10796 14482 10824 14894
rect 10968 14816 11020 14822
rect 10966 14784 10968 14793
rect 11072 14804 11100 16730
rect 11020 14784 11100 14804
rect 11022 14776 11100 14784
rect 10966 14719 11022 14728
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10782 14376 10838 14385
rect 10428 13654 10640 13682
rect 10322 13288 10378 13297
rect 10322 13223 10378 13232
rect 10336 12782 10364 13223
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10230 12336 10286 12345
rect 10230 12271 10286 12280
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10244 11121 10272 12038
rect 10230 11112 10286 11121
rect 10230 11047 10286 11056
rect 10336 10690 10364 12038
rect 10244 10662 10364 10690
rect 10244 10470 10272 10662
rect 10324 10600 10376 10606
rect 10428 10588 10456 13654
rect 10704 13546 10732 14350
rect 11058 14376 11114 14385
rect 10782 14311 10838 14320
rect 10876 14340 10928 14346
rect 10796 13841 10824 14311
rect 11058 14311 11114 14320
rect 10876 14282 10928 14288
rect 10888 13870 10916 14282
rect 11072 14074 11100 14311
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11164 13954 11192 17836
rect 11532 17746 11560 18244
rect 11612 18226 11664 18232
rect 11716 18170 11744 19306
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11624 18142 11744 18170
rect 11624 18086 11652 18142
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11704 18080 11756 18086
rect 11808 18068 11836 18294
rect 11756 18040 11836 18068
rect 11704 18022 11756 18028
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11256 17066 11284 17682
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11716 17320 11744 18022
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11624 17292 11744 17320
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11624 16538 11652 17292
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11716 16658 11744 17002
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11244 16516 11296 16522
rect 11624 16510 11744 16538
rect 11244 16458 11296 16464
rect 11256 15910 11284 16458
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 10980 13926 11192 13954
rect 10876 13864 10928 13870
rect 10782 13832 10838 13841
rect 10876 13806 10928 13812
rect 10782 13767 10838 13776
rect 10782 13696 10838 13705
rect 10782 13631 10838 13640
rect 10520 13518 10732 13546
rect 10520 11880 10548 13518
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10612 13297 10640 13398
rect 10796 13326 10824 13631
rect 10784 13320 10836 13326
rect 10598 13288 10654 13297
rect 10784 13262 10836 13268
rect 10598 13223 10654 13232
rect 10692 13252 10744 13258
rect 10612 13190 10640 13223
rect 10692 13194 10744 13200
rect 10600 13184 10652 13190
rect 10704 13161 10732 13194
rect 10600 13126 10652 13132
rect 10690 13152 10746 13161
rect 10690 13087 10746 13096
rect 10796 12782 10824 13262
rect 10784 12776 10836 12782
rect 10704 12736 10784 12764
rect 10598 12472 10654 12481
rect 10598 12407 10600 12416
rect 10652 12407 10654 12416
rect 10600 12378 10652 12384
rect 10520 11852 10640 11880
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10520 11014 10548 11698
rect 10612 11098 10640 11852
rect 10704 11354 10732 12736
rect 10784 12718 10836 12724
rect 10888 12646 10916 13806
rect 10980 12986 11008 13926
rect 11058 13288 11114 13297
rect 11058 13223 11114 13232
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 11072 12918 11100 13223
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10782 12472 10838 12481
rect 10782 12407 10838 12416
rect 10968 12436 11020 12442
rect 10796 12306 10824 12407
rect 10968 12378 11020 12384
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10874 12200 10930 12209
rect 10874 12135 10930 12144
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10612 11070 10732 11098
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10520 10690 10548 10950
rect 10612 10810 10640 10950
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10520 10662 10640 10690
rect 10612 10588 10640 10662
rect 10376 10560 10456 10588
rect 10324 10542 10376 10548
rect 10428 10470 10456 10560
rect 10520 10560 10640 10588
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10152 9982 10272 10010
rect 10140 9920 10192 9926
rect 10046 9888 10102 9897
rect 10140 9862 10192 9868
rect 10046 9823 10102 9832
rect 10152 9761 10180 9862
rect 10138 9752 10194 9761
rect 10138 9687 10194 9696
rect 10138 9072 10194 9081
rect 10138 9007 10194 9016
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9784 8078 9996 8106
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9600 7806 9720 7834
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9312 6734 9364 6740
rect 8996 6616 9076 6644
rect 8944 6598 8996 6604
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8680 5234 8708 6258
rect 8772 6186 8800 6598
rect 8956 6322 8984 6598
rect 9232 6338 9260 6734
rect 9416 6718 9536 6746
rect 9312 6656 9364 6662
rect 9310 6624 9312 6633
rect 9364 6624 9366 6633
rect 9310 6559 9366 6568
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9140 6310 9260 6338
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 9140 5896 9168 6310
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 8956 5868 9168 5896
rect 8956 5778 8984 5868
rect 9126 5808 9182 5817
rect 8944 5772 8996 5778
rect 9126 5743 9182 5752
rect 8944 5714 8996 5720
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8758 5536 8814 5545
rect 8758 5471 8814 5480
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8772 5098 8800 5471
rect 9048 5234 9076 5646
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 9140 4690 9168 5743
rect 9232 4826 9260 6190
rect 9312 6180 9364 6186
rect 9416 6168 9444 6718
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6322 9536 6598
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9364 6140 9444 6168
rect 9312 6122 9364 6128
rect 9324 5953 9352 6122
rect 9310 5944 9366 5953
rect 9310 5879 9366 5888
rect 9600 5642 9628 6938
rect 9692 6798 9720 7806
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9784 6497 9812 7958
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9876 7002 9904 7210
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9770 6488 9826 6497
rect 9770 6423 9826 6432
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9324 4758 9352 5170
rect 9312 4752 9364 4758
rect 9312 4694 9364 4700
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 8576 4616 8628 4622
rect 8496 4576 8576 4604
rect 8576 4558 8628 4564
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8114 2952 8170 2961
rect 8114 2887 8170 2896
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 7932 1624 7984 1630
rect 7932 1566 7984 1572
rect 7668 870 7788 898
rect 7668 762 7696 870
rect 7760 800 7788 870
rect 8128 800 8156 2887
rect 8206 2680 8262 2689
rect 8206 2615 8208 2624
rect 8260 2615 8262 2624
rect 8208 2586 8260 2592
rect 8312 2514 8340 3334
rect 8496 2582 8524 4082
rect 8760 4004 8812 4010
rect 8680 3964 8760 3992
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 3097 8616 3878
rect 8680 3738 8708 3964
rect 8760 3946 8812 3952
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8574 3088 8630 3097
rect 8574 3023 8630 3032
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8220 1698 8248 2246
rect 8208 1692 8260 1698
rect 8208 1634 8260 1640
rect 8496 800 8524 2518
rect 8588 2514 8616 2790
rect 8680 2530 8708 3538
rect 9140 3534 9168 4626
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 8772 3194 8800 3470
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 9232 3126 9260 4422
rect 9310 4312 9366 4321
rect 9508 4282 9536 5170
rect 9310 4247 9366 4256
rect 9496 4276 9548 4282
rect 9324 4146 9352 4247
rect 9496 4218 9548 4224
rect 9600 4162 9628 5578
rect 9678 5400 9734 5409
rect 9678 5335 9734 5344
rect 9772 5364 9824 5370
rect 9692 5001 9720 5335
rect 9772 5306 9824 5312
rect 9678 4992 9734 5001
rect 9678 4927 9734 4936
rect 9784 4622 9812 5306
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9312 4140 9364 4146
rect 9600 4134 9812 4162
rect 9312 4082 9364 4088
rect 9324 3670 9352 4082
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9312 3664 9364 3670
rect 9312 3606 9364 3612
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9324 2990 9352 3470
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9508 2774 9536 3402
rect 9600 2922 9628 4014
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3466 9720 3878
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9784 3194 9812 4134
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9876 3074 9904 5578
rect 9968 4554 9996 8078
rect 10060 7954 10088 8570
rect 10152 8022 10180 9007
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 10244 7750 10272 9982
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7546 10272 7686
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10060 7177 10088 7414
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10152 7206 10180 7346
rect 10140 7200 10192 7206
rect 10046 7168 10102 7177
rect 10244 7177 10272 7482
rect 10140 7142 10192 7148
rect 10230 7168 10286 7177
rect 10046 7103 10102 7112
rect 10230 7103 10286 7112
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9968 3534 9996 4014
rect 10060 3670 10088 5850
rect 10152 5710 10180 6122
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10152 5370 10180 5646
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10152 4536 10180 4966
rect 10244 4690 10272 6598
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10232 4548 10284 4554
rect 10152 4508 10232 4536
rect 10232 4490 10284 4496
rect 10138 4040 10194 4049
rect 10138 3975 10194 3984
rect 10152 3738 10180 3975
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 9956 3528 10008 3534
rect 10152 3505 10180 3674
rect 9956 3470 10008 3476
rect 10138 3496 10194 3505
rect 10138 3431 10194 3440
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9784 3046 9904 3074
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 9508 2746 9628 2774
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 9404 2576 9456 2582
rect 8576 2508 8628 2514
rect 8680 2502 8892 2530
rect 9404 2518 9456 2524
rect 8576 2450 8628 2456
rect 8864 800 8892 2502
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 800 9260 2246
rect 9416 1902 9444 2518
rect 9600 2378 9628 2746
rect 9588 2372 9640 2378
rect 9588 2314 9640 2320
rect 9404 1896 9456 1902
rect 9404 1838 9456 1844
rect 9784 1766 9812 3046
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9876 1902 9904 2382
rect 9864 1896 9916 1902
rect 9864 1838 9916 1844
rect 9772 1760 9824 1766
rect 9772 1702 9824 1708
rect 9588 1624 9640 1630
rect 9588 1566 9640 1572
rect 9600 800 9628 1566
rect 9968 800 9996 3334
rect 10138 3224 10194 3233
rect 10138 3159 10140 3168
rect 10192 3159 10194 3168
rect 10140 3130 10192 3136
rect 10138 2544 10194 2553
rect 10336 2514 10364 10406
rect 10520 10130 10548 10560
rect 10704 10554 10732 11070
rect 10796 10985 10824 12038
rect 10888 11286 10916 12135
rect 10980 11937 11008 12378
rect 11072 12306 11100 12582
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10966 11928 11022 11937
rect 10966 11863 11022 11872
rect 11072 11830 11100 12242
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 11164 11642 11192 13126
rect 11256 12442 11284 15846
rect 11440 15434 11468 16118
rect 11716 15609 11744 16510
rect 11808 16250 11836 17478
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11900 16182 11928 19790
rect 12084 19514 12112 19790
rect 12176 19786 12204 20402
rect 12440 19984 12492 19990
rect 12492 19944 12572 19972
rect 12440 19926 12492 19932
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12268 19446 12296 19858
rect 12544 19514 12572 19944
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12624 19712 12676 19718
rect 12820 19689 12848 19722
rect 12624 19654 12676 19660
rect 12806 19680 12862 19689
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 12072 19372 12124 19378
rect 12268 19334 12296 19382
rect 12072 19314 12124 19320
rect 12084 18834 12112 19314
rect 12176 19306 12296 19334
rect 12452 19334 12480 19450
rect 12452 19306 12572 19334
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12176 18714 12204 19306
rect 12544 18902 12572 19306
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 12084 18686 12204 18714
rect 11992 18222 12020 18634
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11992 16998 12020 17138
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11992 15994 12020 16934
rect 12084 16697 12112 18686
rect 12360 18630 12388 18838
rect 12440 18760 12492 18766
rect 12636 18714 12664 19654
rect 12806 19615 12862 19624
rect 12912 19446 12940 19790
rect 12900 19440 12952 19446
rect 12900 19382 12952 19388
rect 12900 19168 12952 19174
rect 12806 19136 12862 19145
rect 12900 19110 12952 19116
rect 12806 19071 12862 19080
rect 12440 18702 12492 18708
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12176 17882 12204 18158
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12176 16998 12204 17682
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12360 16794 12388 17818
rect 12452 17542 12480 18702
rect 12544 18686 12664 18714
rect 12544 18154 12572 18686
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12636 18426 12664 18566
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 17354 12572 17478
rect 12452 17326 12572 17354
rect 12728 17338 12756 18158
rect 12820 17796 12848 19071
rect 12912 18766 12940 19110
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12912 18358 12940 18702
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 13004 18034 13032 21383
rect 13096 20602 13124 22200
rect 13464 20602 13492 22200
rect 13832 20602 13860 22200
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13452 20596 13504 20602
rect 13452 20538 13504 20544
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13096 20058 13124 20402
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13188 19990 13216 20402
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 13372 20058 13400 20334
rect 13544 20324 13596 20330
rect 13544 20266 13596 20272
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13176 19984 13228 19990
rect 13176 19926 13228 19932
rect 13268 19848 13320 19854
rect 13188 19796 13268 19802
rect 13188 19790 13320 19796
rect 13188 19774 13308 19790
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 13096 18222 13124 19246
rect 13188 19174 13216 19774
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13004 18006 13124 18034
rect 12990 17912 13046 17921
rect 12990 17847 13046 17856
rect 12900 17808 12952 17814
rect 12820 17768 12900 17796
rect 12900 17750 12952 17756
rect 13004 17338 13032 17847
rect 12716 17332 12768 17338
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12452 16726 12480 17326
rect 12716 17274 12768 17280
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12440 16720 12492 16726
rect 12070 16688 12126 16697
rect 12440 16662 12492 16668
rect 12070 16623 12126 16632
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12360 16153 12388 16390
rect 12162 16144 12218 16153
rect 12162 16079 12218 16088
rect 12346 16144 12402 16153
rect 12346 16079 12402 16088
rect 11992 15966 12112 15994
rect 12084 15910 12112 15966
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 11702 15600 11758 15609
rect 11702 15535 11758 15544
rect 11992 15502 12020 15846
rect 12084 15706 12112 15846
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11428 15428 11480 15434
rect 11428 15370 11480 15376
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11716 15026 11744 15438
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11888 14408 11940 14414
rect 11992 14396 12020 15438
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11940 14368 12020 14396
rect 11888 14350 11940 14356
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11348 13190 11376 13806
rect 11532 13705 11560 13942
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 11518 13696 11574 13705
rect 11518 13631 11574 13640
rect 11624 13258 11652 13738
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11336 12164 11388 12170
rect 11256 12124 11336 12152
rect 11256 11898 11284 12124
rect 11336 12106 11388 12112
rect 11440 12084 11468 12922
rect 11716 12866 11744 14282
rect 11886 14240 11942 14249
rect 11886 14175 11942 14184
rect 11794 14104 11850 14113
rect 11794 14039 11796 14048
rect 11848 14039 11850 14048
rect 11796 14010 11848 14016
rect 11796 13864 11848 13870
rect 11794 13832 11796 13841
rect 11848 13832 11850 13841
rect 11794 13767 11850 13776
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11808 12889 11836 13262
rect 11532 12850 11744 12866
rect 11520 12844 11744 12850
rect 11572 12838 11744 12844
rect 11794 12880 11850 12889
rect 11794 12815 11850 12824
rect 11520 12786 11572 12792
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11440 12056 11744 12084
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 10980 11614 11192 11642
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10782 10976 10838 10985
rect 10782 10911 10838 10920
rect 10874 10840 10930 10849
rect 10874 10775 10930 10784
rect 10704 10526 10824 10554
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10428 8090 10456 9318
rect 10520 9042 10548 9454
rect 10612 9110 10640 10066
rect 10704 10033 10732 10406
rect 10690 10024 10746 10033
rect 10690 9959 10746 9968
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10612 8566 10640 9046
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10612 7954 10640 8502
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10704 7886 10732 9862
rect 10796 9722 10824 10526
rect 10888 10266 10916 10775
rect 10980 10452 11008 11614
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11072 10713 11100 11494
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11058 10704 11114 10713
rect 11164 10674 11192 10950
rect 11058 10639 11114 10648
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11256 10606 11284 11834
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11440 11626 11468 11766
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11612 11552 11664 11558
rect 11610 11520 11612 11529
rect 11664 11520 11666 11529
rect 11610 11455 11666 11464
rect 11716 11354 11744 12056
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11440 11132 11468 11290
rect 11808 11218 11836 12106
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11704 11144 11756 11150
rect 11440 11104 11704 11132
rect 11704 11086 11756 11092
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11716 10742 11744 10950
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11704 10464 11756 10470
rect 10980 10424 11284 10452
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11072 9722 11100 9862
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 11164 9194 11192 9862
rect 11072 9178 11192 9194
rect 11060 9172 11192 9178
rect 11112 9166 11192 9172
rect 11060 9114 11112 9120
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 10874 8664 10930 8673
rect 10874 8599 10930 8608
rect 10888 8566 10916 8599
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 11164 8362 11192 8910
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11164 8090 11192 8298
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10796 7478 10824 8026
rect 10876 8016 10928 8022
rect 11256 7993 11284 10424
rect 11704 10406 11756 10412
rect 11518 10024 11574 10033
rect 11518 9959 11520 9968
rect 11572 9959 11574 9968
rect 11520 9930 11572 9936
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11716 9722 11744 10406
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11716 9110 11744 9522
rect 11808 9518 11836 11154
rect 11900 10810 11928 14175
rect 11992 13938 12020 14368
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 12084 13530 12112 15370
rect 12176 14074 12204 16079
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12268 15094 12296 15642
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12268 14074 12296 15030
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12256 13864 12308 13870
rect 12254 13832 12256 13841
rect 12308 13832 12310 13841
rect 12254 13767 12310 13776
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12256 13456 12308 13462
rect 11978 13424 12034 13433
rect 12254 13424 12256 13433
rect 12308 13424 12310 13433
rect 11978 13359 12034 13368
rect 12164 13388 12216 13394
rect 11992 12889 12020 13359
rect 12254 13359 12310 13368
rect 12164 13330 12216 13336
rect 12176 13274 12204 13330
rect 12084 13246 12204 13274
rect 11978 12880 12034 12889
rect 11978 12815 12034 12824
rect 11978 12472 12034 12481
rect 11978 12407 11980 12416
rect 12032 12407 12034 12416
rect 11980 12378 12032 12384
rect 11978 12200 12034 12209
rect 11978 12135 12034 12144
rect 11992 11014 12020 12135
rect 12084 11150 12112 13246
rect 12164 13184 12216 13190
rect 12162 13152 12164 13161
rect 12216 13152 12218 13161
rect 12162 13087 12218 13096
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12176 11626 12204 12922
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12268 11801 12296 12378
rect 12360 12238 12388 16079
rect 12544 15502 12572 17070
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12636 15570 12664 16934
rect 13096 16289 13124 18006
rect 13082 16280 13138 16289
rect 13082 16215 13138 16224
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12544 15065 12572 15438
rect 12530 15056 12586 15065
rect 12530 14991 12586 15000
rect 12728 14958 12756 15574
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12438 13696 12494 13705
rect 12438 13631 12494 13640
rect 12452 13530 12480 13631
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12544 12889 12572 13398
rect 12530 12880 12586 12889
rect 12530 12815 12586 12824
rect 12532 12776 12584 12782
rect 12452 12736 12532 12764
rect 12452 12306 12480 12736
rect 12532 12718 12584 12724
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12348 12232 12400 12238
rect 12544 12186 12572 12310
rect 12348 12174 12400 12180
rect 12452 12158 12572 12186
rect 12254 11792 12310 11801
rect 12254 11727 12310 11736
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11900 10062 11928 10746
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11794 9344 11850 9353
rect 11794 9279 11850 9288
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11334 8528 11390 8537
rect 11334 8463 11336 8472
rect 11388 8463 11390 8472
rect 11336 8434 11388 8440
rect 11716 8430 11744 8910
rect 11808 8634 11836 9279
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11716 8090 11744 8366
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 10876 7958 10928 7964
rect 11242 7984 11298 7993
rect 10600 7472 10652 7478
rect 10506 7440 10562 7449
rect 10600 7414 10652 7420
rect 10784 7472 10836 7478
rect 10784 7414 10836 7420
rect 10506 7375 10562 7384
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10428 6254 10456 6666
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10428 5914 10456 6190
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10428 4690 10456 5850
rect 10520 5370 10548 7375
rect 10612 6780 10640 7414
rect 10784 6792 10836 6798
rect 10612 6752 10784 6780
rect 10784 6734 10836 6740
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10506 4856 10562 4865
rect 10506 4791 10562 4800
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10138 2479 10194 2488
rect 10324 2508 10376 2514
rect 10152 2446 10180 2479
rect 10324 2450 10376 2456
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10244 2038 10272 2246
rect 10232 2032 10284 2038
rect 10232 1974 10284 1980
rect 10336 800 10364 2450
rect 10520 1748 10548 4791
rect 10612 4622 10640 6054
rect 10796 5778 10824 6054
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10690 5672 10746 5681
rect 10690 5607 10746 5616
rect 10784 5636 10836 5642
rect 10704 5098 10732 5607
rect 10784 5578 10836 5584
rect 10796 5166 10824 5578
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10796 4758 10824 5102
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10796 4146 10824 4422
rect 10888 4162 10916 7958
rect 11242 7919 11298 7928
rect 11808 7886 11836 8230
rect 11796 7880 11848 7886
rect 11702 7848 11758 7857
rect 11796 7822 11848 7828
rect 11702 7783 11758 7792
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10980 7392 11008 7686
rect 11072 7585 11100 7686
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11058 7576 11114 7585
rect 11346 7579 11654 7588
rect 11058 7511 11114 7520
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11428 7472 11480 7478
rect 11716 7449 11744 7783
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11808 7585 11836 7686
rect 11794 7576 11850 7585
rect 11794 7511 11796 7520
rect 11848 7511 11850 7520
rect 11796 7482 11848 7488
rect 11808 7451 11836 7482
rect 11428 7414 11480 7420
rect 11702 7440 11758 7449
rect 11060 7404 11112 7410
rect 10980 7364 11060 7392
rect 11060 7346 11112 7352
rect 11164 7274 11192 7414
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11164 7002 11192 7210
rect 11440 7206 11468 7414
rect 11702 7375 11758 7384
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11716 7041 11744 7142
rect 11702 7032 11758 7041
rect 11152 6996 11204 7002
rect 11808 7002 11836 7278
rect 11900 7018 11928 9658
rect 11992 7410 12020 10678
rect 12084 10606 12112 10746
rect 12176 10742 12204 11562
rect 12268 11200 12296 11562
rect 12360 11354 12388 11698
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12348 11212 12400 11218
rect 12268 11172 12348 11200
rect 12348 11154 12400 11160
rect 12360 10810 12388 11154
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12164 10736 12216 10742
rect 12164 10678 12216 10684
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 12176 10198 12204 10678
rect 12452 10674 12480 12158
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 11898 12572 12038
rect 12636 11898 12664 14758
rect 12728 14346 12756 14894
rect 12820 14657 12848 15574
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12806 14648 12862 14657
rect 12806 14583 12862 14592
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12530 11792 12586 11801
rect 12636 11762 12664 11834
rect 12530 11727 12586 11736
rect 12624 11756 12676 11762
rect 12544 11608 12572 11727
rect 12624 11698 12676 11704
rect 12544 11580 12664 11608
rect 12530 10976 12586 10985
rect 12530 10911 12586 10920
rect 12256 10668 12308 10674
rect 12440 10668 12492 10674
rect 12308 10628 12388 10656
rect 12256 10610 12308 10616
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12176 9450 12204 9862
rect 12268 9722 12296 10406
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12070 8664 12126 8673
rect 12070 8599 12126 8608
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11702 6967 11758 6976
rect 11796 6996 11848 7002
rect 11152 6938 11204 6944
rect 11900 6990 12020 7018
rect 11796 6938 11848 6944
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10980 6361 11008 6394
rect 10966 6352 11022 6361
rect 10966 6287 11022 6296
rect 10980 5914 11008 6287
rect 11072 5914 11100 6394
rect 11164 6254 11192 6802
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11060 5568 11112 5574
rect 11058 5536 11060 5545
rect 11112 5536 11114 5545
rect 11058 5471 11114 5480
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10980 4758 11008 5170
rect 11072 5098 11100 5306
rect 11164 5250 11192 5714
rect 11256 5352 11284 6598
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11518 6080 11574 6089
rect 11518 6015 11574 6024
rect 11334 5944 11390 5953
rect 11334 5879 11336 5888
rect 11388 5879 11390 5888
rect 11336 5850 11388 5856
rect 11532 5574 11560 6015
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11336 5364 11388 5370
rect 11256 5324 11336 5352
rect 11336 5306 11388 5312
rect 11164 5222 11284 5250
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 11256 4690 11284 5222
rect 11612 5160 11664 5166
rect 11334 5128 11390 5137
rect 11612 5102 11664 5108
rect 11334 5063 11390 5072
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 10784 4140 10836 4146
rect 10888 4134 11008 4162
rect 10784 4082 10836 4088
rect 10980 4078 11008 4134
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10874 3904 10930 3913
rect 10874 3839 10930 3848
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10704 3058 10732 3674
rect 10888 3194 10916 3839
rect 11256 3738 11284 4626
rect 11348 4554 11376 5063
rect 11624 5030 11652 5102
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11440 4622 11468 4966
rect 11716 4826 11744 6598
rect 11808 5846 11836 6598
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 5234 11836 5510
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11808 4865 11836 5170
rect 11794 4856 11850 4865
rect 11704 4820 11756 4826
rect 11794 4791 11850 4800
rect 11704 4762 11756 4768
rect 11900 4706 11928 6802
rect 11992 5953 12020 6990
rect 11978 5944 12034 5953
rect 11978 5879 12034 5888
rect 11978 5400 12034 5409
rect 11978 5335 12034 5344
rect 11716 4678 11928 4706
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11716 4282 11744 4678
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4321 11928 4422
rect 11886 4312 11942 4321
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11796 4276 11848 4282
rect 11886 4247 11942 4256
rect 11796 4218 11848 4224
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10692 2440 10744 2446
rect 10690 2408 10692 2417
rect 10744 2408 10746 2417
rect 10690 2343 10746 2352
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10612 1873 10640 2246
rect 10796 2106 10824 2450
rect 10784 2100 10836 2106
rect 10784 2042 10836 2048
rect 10598 1864 10654 1873
rect 10888 1834 10916 3130
rect 10598 1799 10654 1808
rect 10876 1828 10928 1834
rect 10876 1770 10928 1776
rect 10520 1720 10732 1748
rect 10704 800 10732 1720
rect 10980 1612 11008 3334
rect 11150 3224 11206 3233
rect 11150 3159 11206 3168
rect 11164 3126 11192 3159
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 11256 2922 11284 3402
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11716 2854 11744 3878
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11164 2582 11192 2790
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 10980 1584 11100 1612
rect 11072 800 11100 1584
rect 11164 1222 11192 2246
rect 11256 2088 11284 2314
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11256 2060 11468 2088
rect 11152 1216 11204 1222
rect 11152 1158 11204 1164
rect 11440 800 11468 2060
rect 11716 1970 11744 2382
rect 11704 1964 11756 1970
rect 11704 1906 11756 1912
rect 11808 1698 11836 4218
rect 11886 4040 11942 4049
rect 11886 3975 11942 3984
rect 11900 3738 11928 3975
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11900 2650 11928 3130
rect 11992 2990 12020 5335
rect 12084 3194 12112 8599
rect 12268 8566 12296 8842
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12176 7546 12204 8434
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12268 7750 12296 8366
rect 12360 7970 12388 10628
rect 12440 10610 12492 10616
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12452 8430 12480 9590
rect 12544 9586 12572 10911
rect 12636 9926 12664 11580
rect 12728 11150 12756 14010
rect 12820 13394 12848 14214
rect 12912 14074 12940 14758
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13004 13394 13032 15302
rect 13096 13530 13124 16215
rect 13188 15706 13216 19110
rect 13372 18834 13400 19110
rect 13450 19000 13506 19009
rect 13450 18935 13506 18944
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13464 18698 13492 18935
rect 13452 18692 13504 18698
rect 13452 18634 13504 18640
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13280 18426 13308 18566
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13266 18184 13322 18193
rect 13266 18119 13322 18128
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12820 12084 12848 12718
rect 13004 12374 13032 12854
rect 13188 12850 13216 15506
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12900 12368 12952 12374
rect 12900 12310 12952 12316
rect 12992 12368 13044 12374
rect 12992 12310 13044 12316
rect 12912 12220 12940 12310
rect 13096 12220 13124 12582
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 12912 12192 13124 12220
rect 12900 12096 12952 12102
rect 12820 12056 12900 12084
rect 12900 12038 12952 12044
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12912 11830 12940 12038
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 12900 11824 12952 11830
rect 12900 11766 12952 11772
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12806 11248 12862 11257
rect 12806 11183 12862 11192
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12728 10742 12756 11086
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12820 10130 12848 11183
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12912 10062 12940 11494
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12898 9888 12954 9897
rect 12898 9823 12954 9832
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12622 9616 12678 9625
rect 12532 9580 12584 9586
rect 12622 9551 12678 9560
rect 12716 9580 12768 9586
rect 12532 9522 12584 9528
rect 12636 9042 12664 9551
rect 12716 9522 12768 9528
rect 12728 9382 12756 9522
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12360 7942 12480 7970
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12268 7002 12296 7414
rect 12360 7274 12388 7754
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12360 6866 12388 7210
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12164 6792 12216 6798
rect 12452 6746 12480 7942
rect 12544 7041 12572 8910
rect 12728 8634 12756 9318
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12622 7848 12678 7857
rect 12622 7783 12678 7792
rect 12636 7546 12664 7783
rect 12624 7540 12676 7546
rect 12820 7528 12848 9658
rect 12912 8974 12940 9823
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12912 7834 12940 8910
rect 13004 8809 13032 11834
rect 13096 10985 13124 12038
rect 13188 11830 13216 12242
rect 13280 11937 13308 18119
rect 13450 17640 13506 17649
rect 13450 17575 13452 17584
rect 13504 17575 13506 17584
rect 13452 17546 13504 17552
rect 13556 17490 13584 20266
rect 13648 20058 13676 20402
rect 14200 20330 14228 22200
rect 14568 20602 14596 22200
rect 14936 20618 14964 22200
rect 14936 20602 15240 20618
rect 14556 20596 14608 20602
rect 14936 20596 15252 20602
rect 14936 20590 15200 20596
rect 14556 20538 14608 20544
rect 15200 20538 15252 20544
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 14188 20324 14240 20330
rect 14188 20266 14240 20272
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13740 19825 13768 19926
rect 13726 19816 13782 19825
rect 13726 19751 13782 19760
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13740 17678 13768 19110
rect 13832 18766 13860 20198
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 14292 20058 14320 20402
rect 14660 20058 14688 20402
rect 14936 20058 14964 20402
rect 15304 20330 15332 22200
rect 15672 20602 15700 22200
rect 16040 22114 16068 22200
rect 16132 22114 16160 22222
rect 16040 22086 16160 22114
rect 16316 20618 16344 22222
rect 16394 22200 16450 23000
rect 16762 22200 16818 23000
rect 16868 22222 17080 22250
rect 16408 20924 16436 22200
rect 16776 22114 16804 22200
rect 16868 22114 16896 22222
rect 16776 22086 16896 22114
rect 16408 20896 16528 20924
rect 16500 20890 16528 20896
rect 16500 20862 16988 20890
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 15660 20596 15712 20602
rect 16316 20590 16436 20618
rect 16960 20602 16988 20862
rect 16408 20584 16436 20590
rect 16580 20596 16632 20602
rect 16408 20556 16580 20584
rect 15660 20538 15712 20544
rect 16580 20538 16632 20544
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 15752 20528 15804 20534
rect 15752 20470 15804 20476
rect 16854 20496 16910 20505
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15580 20058 15608 20402
rect 15764 20058 15792 20470
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 16672 20460 16724 20466
rect 16854 20431 16910 20440
rect 16948 20460 17000 20466
rect 16672 20402 16724 20408
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15948 19990 15976 20402
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 15936 19984 15988 19990
rect 15936 19926 15988 19932
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 15016 19848 15068 19854
rect 15016 19790 15068 19796
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 14108 19514 14136 19790
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 14108 19174 14136 19450
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14096 19168 14148 19174
rect 14096 19110 14148 19116
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 14292 18086 14320 18770
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 13464 17462 13584 17490
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 13372 16590 13400 16934
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13372 16114 13400 16526
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13464 15994 13492 17462
rect 13648 17202 13676 17546
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13740 16998 13768 17478
rect 14200 17202 14228 17614
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13832 16454 13860 17070
rect 14384 17066 14412 19314
rect 14476 19174 14504 19790
rect 14752 19446 14780 19790
rect 15028 19514 15056 19790
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 14556 19372 14608 19378
rect 14608 19332 14688 19360
rect 14556 19314 14608 19320
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14476 17678 14504 18022
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14568 17490 14596 18226
rect 14476 17462 14596 17490
rect 14476 17202 14504 17462
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 14476 16794 14504 17138
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 16250 13860 16390
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 13728 16040 13780 16046
rect 13464 15966 13584 15994
rect 13728 15982 13780 15988
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13372 13326 13400 14758
rect 13464 14074 13492 15370
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13556 13954 13584 15966
rect 13740 15638 13768 15982
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13832 15706 13860 15846
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 13820 15700 13872 15706
rect 14292 15688 14320 16050
rect 14384 15706 14412 16118
rect 13820 15642 13872 15648
rect 14200 15660 14320 15688
rect 14372 15700 14424 15706
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13648 15094 13676 15302
rect 13832 15162 13860 15642
rect 14200 15366 14228 15660
rect 14372 15642 14424 15648
rect 14384 15570 14412 15642
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14188 15360 14240 15366
rect 14186 15328 14188 15337
rect 14240 15328 14242 15337
rect 14186 15263 14242 15272
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 14002 15056 14058 15065
rect 13648 14414 13676 15030
rect 13820 15020 13872 15026
rect 14002 14991 14058 15000
rect 14292 15042 14320 15438
rect 14476 15162 14504 16730
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14568 15366 14596 15914
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14292 15026 14412 15042
rect 14292 15020 14424 15026
rect 14292 15014 14372 15020
rect 13820 14962 13872 14968
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13740 14074 13768 14894
rect 13832 14482 13860 14962
rect 14016 14958 14044 14991
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 14188 14408 14240 14414
rect 14292 14396 14320 15014
rect 14372 14962 14424 14968
rect 14240 14368 14320 14396
rect 14188 14350 14240 14356
rect 13818 14240 13874 14249
rect 13818 14175 13874 14184
rect 14370 14240 14426 14249
rect 14370 14175 14426 14184
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13452 13932 13504 13938
rect 13556 13926 13768 13954
rect 13832 13938 13860 14175
rect 14384 13938 14412 14175
rect 13452 13874 13504 13880
rect 13464 13841 13492 13874
rect 13450 13832 13506 13841
rect 13450 13767 13506 13776
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13358 13016 13414 13025
rect 13358 12951 13360 12960
rect 13412 12951 13414 12960
rect 13360 12922 13412 12928
rect 13556 12442 13584 13466
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13648 12889 13676 13262
rect 13634 12880 13690 12889
rect 13634 12815 13690 12824
rect 13544 12436 13596 12442
rect 13740 12434 13768 13926
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14004 13864 14056 13870
rect 14188 13864 14240 13870
rect 14056 13824 14188 13852
rect 14004 13806 14056 13812
rect 14188 13806 14240 13812
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 13530 13860 13670
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 14292 13433 14320 13874
rect 14384 13734 14412 13874
rect 14568 13841 14596 15302
rect 14554 13832 14610 13841
rect 14554 13767 14610 13776
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14372 13456 14424 13462
rect 14278 13424 14334 13433
rect 14660 13444 14688 19332
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14424 13416 14688 13444
rect 14372 13398 14424 13404
rect 14278 13359 14334 13368
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13832 12850 13860 13262
rect 14292 13002 14320 13359
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14292 12974 14412 13002
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13818 12608 13874 12617
rect 13818 12543 13874 12552
rect 13544 12378 13596 12384
rect 13648 12406 13768 12434
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 13266 11928 13322 11937
rect 13266 11863 13322 11872
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13372 11762 13400 12310
rect 13450 12200 13506 12209
rect 13450 12135 13452 12144
rect 13504 12135 13506 12144
rect 13452 12106 13504 12112
rect 13648 12050 13676 12406
rect 13832 12238 13860 12543
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 14292 12442 14320 12854
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13820 12096 13872 12102
rect 13464 12022 13676 12050
rect 13726 12064 13782 12073
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13188 11354 13216 11630
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13280 11257 13308 11494
rect 13358 11384 13414 11393
rect 13358 11319 13360 11328
rect 13412 11319 13414 11328
rect 13360 11290 13412 11296
rect 13266 11248 13322 11257
rect 13266 11183 13322 11192
rect 13176 11008 13228 11014
rect 13082 10976 13138 10985
rect 13176 10950 13228 10956
rect 13082 10911 13138 10920
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 13096 9722 13124 10746
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13188 9586 13216 10950
rect 13266 10840 13322 10849
rect 13266 10775 13322 10784
rect 13280 10441 13308 10775
rect 13266 10432 13322 10441
rect 13266 10367 13322 10376
rect 13464 9602 13492 12022
rect 13820 12038 13872 12044
rect 13726 11999 13782 12008
rect 13542 11792 13598 11801
rect 13542 11727 13598 11736
rect 13636 11756 13688 11762
rect 13556 10810 13584 11727
rect 13636 11698 13688 11704
rect 13648 11121 13676 11698
rect 13740 11234 13768 11999
rect 13832 11937 13860 12038
rect 13818 11928 13874 11937
rect 13818 11863 13874 11872
rect 14292 11694 14320 12378
rect 14280 11688 14332 11694
rect 13818 11656 13874 11665
rect 14280 11630 14332 11636
rect 14384 11626 14412 12974
rect 14476 11830 14504 13194
rect 14554 12744 14610 12753
rect 14554 12679 14610 12688
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 13818 11591 13874 11600
rect 14372 11620 14424 11626
rect 13832 11354 13860 11591
rect 14372 11562 14424 11568
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 14476 11354 14504 11766
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 13740 11206 13860 11234
rect 13634 11112 13690 11121
rect 13634 11047 13636 11056
rect 13688 11047 13690 11056
rect 13636 11018 13688 11024
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10130 13768 10406
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13740 9654 13768 10066
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13280 9574 13492 9602
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13174 9480 13230 9489
rect 13096 9178 13124 9454
rect 13174 9415 13230 9424
rect 13188 9178 13216 9415
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13176 8832 13228 8838
rect 12990 8800 13046 8809
rect 13176 8774 13228 8780
rect 12990 8735 13046 8744
rect 13188 8634 13216 8774
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13004 8294 13032 8434
rect 13176 8424 13228 8430
rect 13082 8392 13138 8401
rect 13176 8366 13228 8372
rect 13082 8327 13084 8336
rect 13136 8327 13138 8336
rect 13084 8298 13136 8304
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13004 8090 13032 8230
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13082 7984 13138 7993
rect 13082 7919 13138 7928
rect 12912 7806 13032 7834
rect 12624 7482 12676 7488
rect 12728 7500 12848 7528
rect 12898 7576 12954 7585
rect 12898 7511 12954 7520
rect 12530 7032 12586 7041
rect 12530 6967 12586 6976
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12164 6734 12216 6740
rect 12176 5692 12204 6734
rect 12360 6718 12480 6746
rect 12256 5704 12308 5710
rect 12176 5664 12256 5692
rect 12256 5646 12308 5652
rect 12360 5370 12388 6718
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12452 5914 12480 6190
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12438 5672 12494 5681
rect 12438 5607 12494 5616
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12176 4282 12204 5306
rect 12452 5137 12480 5607
rect 12438 5128 12494 5137
rect 12256 5092 12308 5098
rect 12438 5063 12494 5072
rect 12256 5034 12308 5040
rect 12268 4622 12296 5034
rect 12346 4992 12402 5001
rect 12346 4927 12402 4936
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12360 4554 12388 4927
rect 12544 4554 12572 6870
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12636 6118 12664 6394
rect 12728 6322 12756 7500
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12820 6780 12848 7346
rect 12912 7342 12940 7511
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12900 6792 12952 6798
rect 12820 6752 12900 6780
rect 12900 6734 12952 6740
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12636 5681 12664 5850
rect 12912 5681 12940 6054
rect 12622 5672 12678 5681
rect 12622 5607 12678 5616
rect 12898 5672 12954 5681
rect 12898 5607 12954 5616
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12636 5370 12664 5510
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12728 5250 12756 5306
rect 12636 5222 12756 5250
rect 12900 5228 12952 5234
rect 12636 4758 12664 5222
rect 12900 5170 12952 5176
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12162 3496 12218 3505
rect 12162 3431 12218 3440
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12176 3126 12204 3431
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 12070 2952 12126 2961
rect 12070 2887 12126 2896
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12084 2446 12112 2887
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 12176 2446 12204 2790
rect 12268 2582 12296 4422
rect 12636 4282 12664 4422
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12360 3738 12388 3878
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12452 3534 12480 3878
rect 12544 3602 12572 3946
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12438 3224 12494 3233
rect 12438 3159 12494 3168
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11900 2106 11928 2246
rect 11888 2100 11940 2106
rect 11888 2042 11940 2048
rect 11796 1692 11848 1698
rect 11796 1634 11848 1640
rect 11808 870 11928 898
rect 11808 800 11836 870
rect 7484 734 7696 762
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 11900 762 11928 870
rect 12084 762 12112 2382
rect 12452 2378 12480 3159
rect 12636 2650 12664 4082
rect 12728 3641 12756 4966
rect 12912 4826 12940 5170
rect 13004 5137 13032 7806
rect 13096 7750 13124 7919
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13096 7206 13124 7686
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12990 5128 13046 5137
rect 12990 5063 13046 5072
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 13004 4604 13032 4966
rect 13096 4826 13124 7142
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12912 4576 13032 4604
rect 12912 4298 12940 4576
rect 13188 4554 13216 8366
rect 13280 6905 13308 9574
rect 13452 9512 13504 9518
rect 13832 9466 13860 11206
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14476 10849 14504 11154
rect 14462 10840 14518 10849
rect 14372 10804 14424 10810
rect 14424 10784 14462 10792
rect 14424 10775 14518 10784
rect 14424 10764 14504 10775
rect 14372 10746 14424 10752
rect 14476 10715 14504 10764
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14200 9994 14228 10066
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13452 9454 13504 9460
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 9042 13400 9386
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13464 8838 13492 9454
rect 13648 9438 13860 9466
rect 13648 8922 13676 9438
rect 13924 9364 13952 9862
rect 14200 9586 14228 9930
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 13740 9336 13952 9364
rect 13740 9058 13768 9336
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13818 9208 13874 9217
rect 13945 9211 14253 9220
rect 13818 9143 13820 9152
rect 13872 9143 13874 9152
rect 13820 9114 13872 9120
rect 13740 9030 13952 9058
rect 14292 9042 14320 10610
rect 14464 10532 14516 10538
rect 14464 10474 14516 10480
rect 14476 10441 14504 10474
rect 14462 10432 14518 10441
rect 14462 10367 14518 10376
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 13728 8968 13780 8974
rect 13556 8894 13676 8922
rect 13726 8936 13728 8945
rect 13780 8936 13782 8945
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13358 7848 13414 7857
rect 13358 7783 13414 7792
rect 13372 7206 13400 7783
rect 13464 7342 13492 8774
rect 13556 8430 13584 8894
rect 13726 8871 13782 8880
rect 13634 8800 13690 8809
rect 13634 8735 13690 8744
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13450 7032 13506 7041
rect 13450 6967 13506 6976
rect 13266 6896 13322 6905
rect 13322 6840 13400 6848
rect 13266 6831 13400 6840
rect 13280 6820 13400 6831
rect 13266 6760 13322 6769
rect 13266 6695 13322 6704
rect 13280 6458 13308 6695
rect 13372 6458 13400 6820
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13372 6118 13400 6258
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13372 5545 13400 6054
rect 13358 5536 13414 5545
rect 13358 5471 13414 5480
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 12820 4270 12940 4298
rect 12992 4276 13044 4282
rect 12820 4146 12848 4270
rect 12992 4218 13044 4224
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12714 3632 12770 3641
rect 12714 3567 12770 3576
rect 12820 3466 12848 4082
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 12820 3194 12848 3402
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12912 2446 12940 3878
rect 13004 3618 13032 4218
rect 13096 4146 13124 4422
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13188 3913 13216 4490
rect 13174 3904 13230 3913
rect 13174 3839 13230 3848
rect 13280 3738 13308 5034
rect 13372 5001 13400 5471
rect 13358 4992 13414 5001
rect 13358 4927 13414 4936
rect 13358 4584 13414 4593
rect 13358 4519 13414 4528
rect 13372 4486 13400 4519
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13464 4298 13492 6967
rect 13372 4270 13492 4298
rect 13372 3890 13400 4270
rect 13556 4214 13584 8366
rect 13648 6866 13676 8735
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13740 7886 13768 8570
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13740 7041 13768 7142
rect 13726 7032 13782 7041
rect 13726 6967 13782 6976
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13832 6746 13860 8298
rect 13924 8276 13952 9030
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14002 8664 14058 8673
rect 14002 8599 14004 8608
rect 14056 8599 14058 8608
rect 14004 8570 14056 8576
rect 14108 8498 14136 8774
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 13924 8248 14320 8276
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 14016 7546 14044 8026
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14292 7410 14320 8248
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 14188 6860 14240 6866
rect 14292 6848 14320 7142
rect 14240 6820 14320 6848
rect 14188 6802 14240 6808
rect 13832 6718 13952 6746
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 6390 13860 6598
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13924 6322 13952 6718
rect 14200 6390 14228 6802
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13924 6202 13952 6258
rect 13832 6174 13952 6202
rect 14278 6216 14334 6225
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 13648 4026 13676 5510
rect 13740 5216 13768 5714
rect 13832 5710 13860 6174
rect 14278 6151 14334 6160
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 14292 5846 14320 6151
rect 14280 5840 14332 5846
rect 14280 5782 14332 5788
rect 14384 5794 14412 10202
rect 14568 10062 14596 12679
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14660 11937 14688 12106
rect 14646 11928 14702 11937
rect 14646 11863 14702 11872
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14660 11354 14688 11630
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14476 9110 14504 9590
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14568 9178 14596 9522
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14568 8294 14596 8774
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7750 14596 8230
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14476 6798 14504 7686
rect 14568 7449 14596 7686
rect 14554 7440 14610 7449
rect 14554 7375 14610 7384
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14568 5817 14596 6666
rect 14554 5808 14610 5817
rect 14384 5766 14504 5794
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14108 5409 14136 5510
rect 14094 5400 14150 5409
rect 14094 5335 14150 5344
rect 14384 5234 14412 5646
rect 13820 5228 13872 5234
rect 13740 5188 13820 5216
rect 13820 5170 13872 5176
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 13832 4758 13860 5170
rect 14476 5166 14504 5766
rect 14554 5743 14610 5752
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14372 5092 14424 5098
rect 14292 5052 14372 5080
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13740 4282 13768 4626
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13464 4010 13676 4026
rect 13452 4004 13676 4010
rect 13504 3998 13676 4004
rect 13452 3946 13504 3952
rect 13372 3862 13584 3890
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13004 3590 13124 3618
rect 13096 2938 13124 3590
rect 13188 3058 13216 3674
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13096 2910 13216 2938
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 13096 2514 13124 2790
rect 13084 2508 13136 2514
rect 13084 2450 13136 2456
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12532 2372 12584 2378
rect 12532 2314 12584 2320
rect 12164 1964 12216 1970
rect 12164 1906 12216 1912
rect 12176 800 12204 1906
rect 12544 800 12572 2314
rect 12808 2304 12860 2310
rect 12860 2264 12940 2292
rect 12808 2246 12860 2252
rect 12912 800 12940 2264
rect 13188 1154 13216 2910
rect 13372 2446 13400 3334
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13464 2854 13492 3130
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13556 2038 13584 3862
rect 13648 2938 13676 3998
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13740 3398 13768 3946
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 3194 13768 3334
rect 13832 3194 13860 4082
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13820 2984 13872 2990
rect 13648 2932 13820 2938
rect 13924 2961 13952 3606
rect 14292 3482 14320 5052
rect 14372 5034 14424 5040
rect 14370 4992 14426 5001
rect 14370 4927 14426 4936
rect 14384 4690 14412 4927
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14200 3454 14320 3482
rect 14200 3233 14228 3454
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14186 3224 14242 3233
rect 14186 3159 14242 3168
rect 13648 2926 13872 2932
rect 13910 2952 13966 2961
rect 13648 2910 13860 2926
rect 13910 2887 13966 2896
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13726 2680 13782 2689
rect 13945 2683 14253 2692
rect 13726 2615 13782 2624
rect 13912 2644 13964 2650
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13544 2032 13596 2038
rect 13544 1974 13596 1980
rect 13268 1964 13320 1970
rect 13268 1906 13320 1912
rect 13176 1148 13228 1154
rect 13176 1090 13228 1096
rect 13280 800 13308 1906
rect 13648 800 13676 2518
rect 13740 2446 13768 2615
rect 13912 2586 13964 2592
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 13924 2446 13952 2586
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14016 800 14044 2586
rect 14292 2514 14320 3334
rect 14384 3194 14412 4422
rect 14476 3913 14504 4490
rect 14556 3936 14608 3942
rect 14462 3904 14518 3913
rect 14556 3878 14608 3884
rect 14462 3839 14518 3848
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14476 3398 14504 3674
rect 14568 3602 14596 3878
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14660 3210 14688 10542
rect 14752 9926 14780 17478
rect 14844 17338 14872 18566
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14832 15088 14884 15094
rect 14832 15030 14884 15036
rect 14844 14464 14872 15030
rect 14936 14906 14964 19382
rect 15212 19174 15240 19790
rect 15580 19378 15608 19790
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15290 19272 15346 19281
rect 15290 19207 15292 19216
rect 15344 19207 15346 19216
rect 15292 19178 15344 19184
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15028 18086 15056 19110
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 15212 17542 15240 19110
rect 15488 18737 15516 19110
rect 15474 18728 15530 18737
rect 15474 18663 15530 18672
rect 15672 18329 15700 19110
rect 15658 18320 15714 18329
rect 15658 18255 15714 18264
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15120 16250 15148 17070
rect 15212 16454 15240 17070
rect 15304 17066 15332 17478
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 15304 16522 15332 17002
rect 15580 16794 15608 17206
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15120 15502 15148 16050
rect 15304 16046 15332 16458
rect 15672 16250 15700 17478
rect 15764 16561 15792 19790
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16132 19174 16160 19314
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16132 18873 16160 19110
rect 16118 18864 16174 18873
rect 16118 18799 16174 18808
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16040 17542 16068 18022
rect 16316 17921 16344 19654
rect 16408 19446 16436 20198
rect 16684 20058 16712 20402
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16868 19990 16896 20431
rect 16948 20402 17000 20408
rect 16856 19984 16908 19990
rect 16856 19926 16908 19932
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16960 19514 16988 20402
rect 17052 20330 17080 22222
rect 17130 22200 17186 23000
rect 17498 22200 17554 23000
rect 17866 22200 17922 23000
rect 18234 22200 18290 23000
rect 18602 22200 18658 23000
rect 18970 22200 19026 23000
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 20074 22200 20130 23000
rect 20442 22200 20498 23000
rect 20810 22200 20866 23000
rect 21178 22200 21234 23000
rect 21546 22200 21602 23000
rect 21652 22222 21864 22250
rect 17144 20534 17172 22200
rect 17224 20868 17276 20874
rect 17224 20810 17276 20816
rect 17132 20528 17184 20534
rect 17132 20470 17184 20476
rect 17040 20324 17092 20330
rect 17040 20266 17092 20272
rect 17236 20058 17264 20810
rect 17512 20262 17540 22200
rect 17776 21072 17828 21078
rect 17776 21014 17828 21020
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17420 20058 17448 20198
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 17328 19446 17356 19790
rect 17604 19786 17632 20402
rect 17788 19990 17816 21014
rect 17880 20330 17908 22200
rect 18248 20618 18276 22200
rect 18248 20590 18368 20618
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 17868 20324 17920 20330
rect 17868 20266 17920 20272
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 16396 19440 16448 19446
rect 16396 19382 16448 19388
rect 17316 19440 17368 19446
rect 17512 19417 17540 19654
rect 17316 19382 17368 19388
rect 17498 19408 17554 19417
rect 16856 19372 16908 19378
rect 17880 19394 17908 19790
rect 17972 19514 18000 20402
rect 18050 20360 18106 20369
rect 18050 20295 18106 20304
rect 18064 20058 18092 20295
rect 18248 20058 18276 20402
rect 18340 20058 18368 20590
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17880 19378 18000 19394
rect 17880 19372 18012 19378
rect 17880 19366 17960 19372
rect 17498 19343 17554 19352
rect 16856 19314 16908 19320
rect 17960 19314 18012 19320
rect 16868 19174 16896 19314
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16408 18358 16436 19110
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 17972 18426 18000 19314
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 16396 18352 16448 18358
rect 16396 18294 16448 18300
rect 16302 17912 16358 17921
rect 16302 17847 16304 17856
rect 16356 17847 16358 17856
rect 16304 17818 16356 17824
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15856 16794 15884 17138
rect 16040 17082 16068 17478
rect 16040 17054 16252 17082
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 16040 16658 16068 16934
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 15750 16552 15806 16561
rect 15750 16487 15806 16496
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15856 16250 15884 16390
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 15028 15026 15056 15302
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 14936 14878 15056 14906
rect 14844 14436 14964 14464
rect 14832 14340 14884 14346
rect 14832 14282 14884 14288
rect 14844 12238 14872 14282
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14752 7954 14780 9318
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14752 7478 14780 7890
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14752 6934 14780 7414
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14844 6746 14872 12174
rect 14936 11778 14964 14436
rect 15028 13870 15056 14878
rect 15120 14346 15148 15438
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15028 12209 15056 13806
rect 15212 13410 15240 14758
rect 15120 13382 15240 13410
rect 15120 13326 15148 13382
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15212 12986 15240 13194
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 15014 12200 15070 12209
rect 15014 12135 15070 12144
rect 15120 11898 15148 12650
rect 15304 12186 15332 15846
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15764 14958 15792 15370
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15764 14618 15792 14894
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15396 12238 15424 13262
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15212 12158 15332 12186
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 14936 11750 15056 11778
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14936 10010 14964 11630
rect 15028 11218 15056 11750
rect 15212 11694 15240 12158
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 11218 15240 11494
rect 15304 11218 15332 12038
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 15028 10305 15056 11018
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15014 10296 15070 10305
rect 15014 10231 15070 10240
rect 15212 10146 15240 10678
rect 15028 10130 15240 10146
rect 15016 10124 15240 10130
rect 15068 10118 15240 10124
rect 15290 10160 15346 10169
rect 15290 10095 15346 10104
rect 15016 10066 15068 10072
rect 15304 10062 15332 10095
rect 15292 10056 15344 10062
rect 14936 9982 15148 10010
rect 15292 9998 15344 10004
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14936 8634 14964 9386
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15028 8514 15056 9862
rect 15120 9602 15148 9982
rect 15120 9574 15240 9602
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15120 8906 15148 9454
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 14752 6718 14872 6746
rect 14936 8486 15056 8514
rect 14752 6202 14780 6718
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14844 6390 14872 6598
rect 14832 6384 14884 6390
rect 14832 6326 14884 6332
rect 14752 6174 14872 6202
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14752 3942 14780 4694
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14738 3768 14794 3777
rect 14738 3703 14794 3712
rect 14752 3505 14780 3703
rect 14738 3496 14794 3505
rect 14738 3431 14794 3440
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14476 3182 14688 3210
rect 14372 2984 14424 2990
rect 14370 2952 14372 2961
rect 14424 2952 14426 2961
rect 14370 2887 14426 2896
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14292 1970 14320 2246
rect 14476 1970 14504 3182
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14660 2378 14688 2994
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14752 2446 14780 2790
rect 14844 2666 14872 6174
rect 14936 5370 14964 8486
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 15028 7886 15056 8366
rect 15120 8362 15148 8842
rect 15212 8362 15240 9574
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 8634 15332 9318
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 15396 8129 15424 12038
rect 15488 11914 15516 12854
rect 15580 12050 15608 14214
rect 15764 14006 15792 14554
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15752 13864 15804 13870
rect 15856 13852 15884 14282
rect 15948 14074 15976 14894
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15804 13824 15884 13852
rect 15752 13806 15804 13812
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15672 12442 15700 12786
rect 15660 12436 15712 12442
rect 15764 12434 15792 13670
rect 15856 13394 15884 13824
rect 15948 13530 15976 13874
rect 16040 13530 16068 14962
rect 16224 14521 16252 17054
rect 16316 16658 16344 17682
rect 16408 16776 16436 18294
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 16488 16788 16540 16794
rect 16408 16748 16488 16776
rect 16488 16730 16540 16736
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16396 16516 16448 16522
rect 16396 16458 16448 16464
rect 16302 16280 16358 16289
rect 16302 16215 16304 16224
rect 16356 16215 16358 16224
rect 16304 16186 16356 16192
rect 16316 16046 16344 16186
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16210 14512 16266 14521
rect 16210 14447 16266 14456
rect 16118 13968 16174 13977
rect 16118 13903 16174 13912
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15764 12406 15884 12434
rect 15660 12378 15712 12384
rect 15580 12022 15700 12050
rect 15488 11886 15608 11914
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15488 11354 15516 11698
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15474 10024 15530 10033
rect 15474 9959 15530 9968
rect 15488 9926 15516 9959
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15488 8974 15516 9454
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15488 8566 15516 8910
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15382 8120 15438 8129
rect 15200 8084 15252 8090
rect 15382 8055 15438 8064
rect 15200 8026 15252 8032
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15028 7546 15056 7686
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15028 5370 15056 7346
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 14936 4554 14964 5306
rect 15028 5030 15056 5306
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 14924 4548 14976 4554
rect 14924 4490 14976 4496
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 14936 3738 14964 4014
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14936 3058 14964 3334
rect 15028 3194 15056 4014
rect 15016 3188 15068 3194
rect 15016 3130 15068 3136
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14936 2774 14964 2994
rect 14936 2746 15056 2774
rect 14844 2638 14964 2666
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 14280 1964 14332 1970
rect 14280 1906 14332 1912
rect 14464 1964 14516 1970
rect 14464 1906 14516 1912
rect 14568 1170 14596 2246
rect 14936 2106 14964 2638
rect 14924 2100 14976 2106
rect 14924 2042 14976 2048
rect 14740 1828 14792 1834
rect 14740 1770 14792 1776
rect 14384 1142 14596 1170
rect 14384 800 14412 1142
rect 14752 800 14780 1770
rect 15028 1057 15056 2746
rect 15120 2582 15148 7958
rect 15212 7449 15240 8026
rect 15488 7886 15516 8502
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15396 7585 15424 7686
rect 15382 7576 15438 7585
rect 15382 7511 15438 7520
rect 15198 7440 15254 7449
rect 15198 7375 15254 7384
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15198 6896 15254 6905
rect 15198 6831 15200 6840
rect 15252 6831 15254 6840
rect 15200 6802 15252 6808
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15212 5710 15240 6122
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15198 5400 15254 5409
rect 15198 5335 15200 5344
rect 15252 5335 15254 5344
rect 15200 5306 15252 5312
rect 15198 5264 15254 5273
rect 15198 5199 15254 5208
rect 15212 4865 15240 5199
rect 15304 5001 15332 7278
rect 15396 7002 15424 7346
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15290 4992 15346 5001
rect 15290 4927 15346 4936
rect 15198 4856 15254 4865
rect 15198 4791 15254 4800
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15198 4312 15254 4321
rect 15198 4247 15254 4256
rect 15212 3126 15240 4247
rect 15304 3194 15332 4762
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15212 2446 15240 2790
rect 15304 2514 15332 2994
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15108 2372 15160 2378
rect 15108 2314 15160 2320
rect 15014 1048 15070 1057
rect 15014 983 15070 992
rect 15120 800 15148 2314
rect 15396 2038 15424 6802
rect 15488 3924 15516 7822
rect 15580 6866 15608 11886
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15580 6089 15608 6666
rect 15566 6080 15622 6089
rect 15566 6015 15622 6024
rect 15566 5944 15622 5953
rect 15566 5879 15622 5888
rect 15580 5846 15608 5879
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15580 5574 15608 5782
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15672 5370 15700 12022
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15764 10062 15792 10610
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15856 8265 15884 12406
rect 16132 12170 16160 13903
rect 16224 13802 16252 14447
rect 16408 14385 16436 16458
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16960 16250 16988 17070
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17130 16552 17186 16561
rect 17130 16487 17186 16496
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17144 16046 17172 16487
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17328 15706 17356 16594
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16960 15162 16988 15438
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16868 14550 16896 14758
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 17144 14482 17172 15302
rect 17328 15094 17356 15642
rect 17316 15088 17368 15094
rect 17316 15030 17368 15036
rect 17314 14920 17370 14929
rect 17420 14906 17448 17614
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17682 17232 17738 17241
rect 17682 17167 17738 17176
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17370 14878 17448 14906
rect 17314 14855 17370 14864
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 16394 14376 16450 14385
rect 16394 14311 16450 14320
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16224 12238 16252 12786
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15948 11354 15976 12038
rect 16040 11898 16068 12038
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16224 11778 16252 12174
rect 16040 11750 16252 11778
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16040 11150 16068 11750
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16132 11218 16160 11562
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 15948 10810 15976 10950
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 15948 10606 15976 10746
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 16040 10266 16068 10950
rect 16132 10810 16160 11154
rect 16224 11014 16252 11630
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16224 10742 16252 10950
rect 16212 10736 16264 10742
rect 16212 10678 16264 10684
rect 16210 10568 16266 10577
rect 16210 10503 16266 10512
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16026 10160 16082 10169
rect 16026 10095 16082 10104
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15948 9178 15976 9454
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15948 8430 15976 9114
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15842 8256 15898 8265
rect 15842 8191 15898 8200
rect 15856 7818 15884 8191
rect 15934 8120 15990 8129
rect 15934 8055 15990 8064
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15948 7698 15976 8055
rect 15856 7670 15976 7698
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15764 6458 15792 7142
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15672 4554 15700 5306
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 15568 4072 15620 4078
rect 15566 4040 15568 4049
rect 15620 4040 15622 4049
rect 15566 3975 15622 3984
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15488 3896 15608 3924
rect 15580 2922 15608 3896
rect 15672 3534 15700 3946
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15568 2916 15620 2922
rect 15568 2858 15620 2864
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15566 2816 15622 2825
rect 15384 2032 15436 2038
rect 15384 1974 15436 1980
rect 15488 800 15516 2790
rect 15566 2751 15622 2760
rect 15580 1290 15608 2751
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 15672 1834 15700 2246
rect 15764 1902 15792 5646
rect 15856 5302 15884 7670
rect 16040 7342 16068 10095
rect 16132 9761 16160 10406
rect 16224 10266 16252 10503
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16224 10062 16252 10202
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16316 10010 16344 13126
rect 16408 12442 16436 13806
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16592 12186 16620 12650
rect 16764 12640 16816 12646
rect 16762 12608 16764 12617
rect 16816 12608 16818 12617
rect 16762 12543 16818 12552
rect 16960 12306 16988 13330
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16592 12164 16988 12186
rect 17052 12170 17080 12582
rect 16592 12158 16764 12164
rect 16816 12158 16988 12164
rect 16764 12106 16816 12112
rect 16776 12075 16804 12106
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16408 11558 16436 11698
rect 16592 11665 16620 11698
rect 16764 11688 16816 11694
rect 16578 11656 16634 11665
rect 16764 11630 16816 11636
rect 16960 11642 16988 12158
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 17052 11801 17080 12106
rect 17144 11898 17172 14282
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17236 12753 17264 13126
rect 17222 12744 17278 12753
rect 17222 12679 17278 12688
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17038 11792 17094 11801
rect 17038 11727 17094 11736
rect 16578 11591 16634 11600
rect 16396 11552 16448 11558
rect 16394 11520 16396 11529
rect 16448 11520 16450 11529
rect 16394 11455 16450 11464
rect 16592 11098 16620 11591
rect 16776 11150 16804 11630
rect 16960 11614 17080 11642
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16868 11150 16896 11494
rect 16408 11070 16620 11098
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16948 11076 17000 11082
rect 16408 10470 16436 11070
rect 16948 11018 17000 11024
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16960 10810 16988 11018
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 17052 10713 17080 11614
rect 17144 11354 17172 11834
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17038 10704 17094 10713
rect 16948 10668 17000 10674
rect 17038 10639 17094 10648
rect 16948 10610 17000 10616
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16396 10464 16448 10470
rect 16868 10441 16896 10542
rect 16396 10406 16448 10412
rect 16854 10432 16910 10441
rect 16854 10367 16910 10376
rect 16316 9982 16436 10010
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16118 9752 16174 9761
rect 16118 9687 16174 9696
rect 16210 9616 16266 9625
rect 16210 9551 16266 9560
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16028 6928 16080 6934
rect 16028 6870 16080 6876
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15856 3534 15884 5102
rect 15948 4078 15976 6598
rect 16040 6236 16068 6870
rect 16132 6390 16160 8434
rect 16224 8090 16252 9551
rect 16316 8974 16344 9862
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16316 8430 16344 8910
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16408 7478 16436 9982
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16684 9382 16712 9454
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16684 9081 16712 9318
rect 16776 9217 16804 9318
rect 16762 9208 16818 9217
rect 16762 9143 16818 9152
rect 16670 9072 16726 9081
rect 16670 9007 16726 9016
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16120 6384 16172 6390
rect 16120 6326 16172 6332
rect 16040 6208 16160 6236
rect 16132 6118 16160 6208
rect 16224 6186 16252 6734
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15948 3670 15976 4014
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 16040 3534 16068 6054
rect 16118 5808 16174 5817
rect 16118 5743 16120 5752
rect 16172 5743 16174 5752
rect 16120 5714 16172 5720
rect 16120 4208 16172 4214
rect 16120 4150 16172 4156
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15948 3126 15976 3334
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 15936 2848 15988 2854
rect 16132 2825 16160 4150
rect 16224 3058 16252 6122
rect 16316 5817 16344 7210
rect 16408 7002 16436 7414
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16500 6882 16528 7142
rect 16408 6854 16528 6882
rect 16408 6322 16436 6854
rect 16684 6798 16712 7278
rect 16960 6882 16988 10610
rect 17144 9926 17172 11154
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17144 9586 17172 9862
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17052 9178 17080 9522
rect 17236 9466 17264 12038
rect 17328 11558 17356 14855
rect 17512 14618 17540 16594
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17604 16250 17632 16390
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17696 14634 17724 17167
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17788 15434 17816 15982
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17500 14612 17552 14618
rect 17696 14606 17816 14634
rect 17500 14554 17552 14560
rect 17788 14482 17816 14606
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17420 14074 17448 14214
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17408 13796 17460 13802
rect 17408 13738 17460 13744
rect 17420 12646 17448 13738
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17512 13326 17540 13670
rect 17604 13394 17632 13874
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17500 13320 17552 13326
rect 17552 13268 17632 13274
rect 17500 13262 17632 13268
rect 17512 13246 17632 13262
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 11898 17448 12582
rect 17604 12306 17632 13246
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17420 11665 17448 11834
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17406 11656 17462 11665
rect 17406 11591 17462 11600
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17328 11354 17356 11494
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 11014 17356 11086
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17328 10606 17356 10950
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 9586 17356 10066
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17132 9444 17184 9450
rect 17236 9438 17356 9466
rect 17132 9386 17184 9392
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17052 8514 17080 8910
rect 17144 8634 17172 9386
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17052 8486 17172 8514
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 17052 7342 17080 8366
rect 17144 8362 17172 8486
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17236 8294 17264 9318
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17144 7206 17172 7890
rect 17236 7410 17264 8230
rect 17328 7886 17356 9438
rect 17420 8634 17448 11494
rect 17512 9110 17540 11698
rect 17604 11694 17632 12242
rect 17696 11762 17724 13194
rect 17788 11778 17816 14418
rect 17880 12345 17908 17478
rect 18064 15026 18092 19654
rect 18156 16810 18184 19790
rect 18234 19408 18290 19417
rect 18340 19378 18368 19858
rect 18432 19514 18460 20198
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18524 19961 18552 19994
rect 18616 19990 18644 22200
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18604 19984 18656 19990
rect 18510 19952 18566 19961
rect 18604 19926 18656 19932
rect 18510 19887 18566 19896
rect 18420 19508 18472 19514
rect 18420 19450 18472 19456
rect 18234 19343 18236 19352
rect 18288 19343 18290 19352
rect 18328 19372 18380 19378
rect 18236 19314 18288 19320
rect 18328 19314 18380 19320
rect 18340 19174 18368 19314
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18616 18970 18644 19926
rect 18708 19786 18736 20402
rect 18880 20324 18932 20330
rect 18880 20266 18932 20272
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 18800 19514 18828 19790
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18156 16782 18368 16810
rect 18236 16720 18288 16726
rect 18234 16688 18236 16697
rect 18288 16688 18290 16697
rect 18234 16623 18290 16632
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17972 13938 18000 14758
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17972 12374 18000 13874
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18064 12442 18092 12718
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 17960 12368 18012 12374
rect 17866 12336 17922 12345
rect 17960 12310 18012 12316
rect 17866 12271 17922 12280
rect 17684 11756 17736 11762
rect 17788 11750 17908 11778
rect 17684 11698 17736 11704
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 17684 11620 17736 11626
rect 17684 11562 17736 11568
rect 17696 11218 17724 11562
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17604 10810 17632 11018
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17696 10266 17724 11154
rect 17788 10538 17816 11630
rect 17880 11354 17908 11750
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17866 10976 17922 10985
rect 17866 10911 17922 10920
rect 17880 10742 17908 10911
rect 17972 10742 18000 12310
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18064 11354 18092 11698
rect 18156 11558 18184 16526
rect 18340 14278 18368 16782
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18524 16182 18552 16390
rect 18512 16176 18564 16182
rect 18510 16144 18512 16153
rect 18564 16144 18566 16153
rect 18510 16079 18566 16088
rect 18604 16108 18656 16114
rect 18524 15638 18552 16079
rect 18604 16050 18656 16056
rect 18616 15706 18644 16050
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 18248 12986 18276 13194
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 18340 12850 18368 13126
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18248 11898 18276 12786
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18340 11830 18368 12786
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18328 11824 18380 11830
rect 18234 11792 18290 11801
rect 18328 11766 18380 11772
rect 18234 11727 18290 11736
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18248 11098 18276 11727
rect 18248 11070 18368 11098
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17958 10568 18014 10577
rect 17776 10532 17828 10538
rect 17958 10503 18014 10512
rect 17776 10474 17828 10480
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17696 9654 17724 9930
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17512 8294 17540 8434
rect 17604 8362 17632 9590
rect 17788 9489 17816 9930
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17880 9654 17908 9862
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17774 9480 17830 9489
rect 17972 9466 18000 10503
rect 17774 9415 17830 9424
rect 17880 9438 18000 9466
rect 17880 9330 17908 9438
rect 17788 9302 17908 9330
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 17696 8430 17724 8774
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17328 7528 17356 7822
rect 17420 7721 17448 8026
rect 17512 7954 17540 8230
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17406 7712 17462 7721
rect 17406 7647 17462 7656
rect 17328 7500 17540 7528
rect 17224 7404 17276 7410
rect 17408 7404 17460 7410
rect 17224 7346 17276 7352
rect 17328 7364 17408 7392
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 16960 6854 17080 6882
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16960 6458 16988 6598
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17052 6338 17080 6854
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16960 6310 17080 6338
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16578 6216 16634 6225
rect 16302 5808 16358 5817
rect 16500 5778 16528 6190
rect 16578 6151 16634 6160
rect 16592 5914 16620 6151
rect 16960 5953 16988 6310
rect 16946 5944 17002 5953
rect 16580 5908 16632 5914
rect 17144 5930 17172 6938
rect 17236 6798 17264 7346
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17328 6633 17356 7364
rect 17408 7346 17460 7352
rect 17406 7168 17462 7177
rect 17406 7103 17462 7112
rect 17314 6624 17370 6633
rect 17314 6559 17370 6568
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 16946 5879 17002 5888
rect 17052 5902 17172 5930
rect 16580 5850 16632 5856
rect 16302 5743 16358 5752
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16316 5545 16344 5578
rect 16960 5574 16988 5879
rect 16580 5568 16632 5574
rect 16302 5536 16358 5545
rect 16302 5471 16358 5480
rect 16408 5528 16580 5556
rect 16408 5302 16436 5528
rect 16580 5510 16632 5516
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16396 5296 16448 5302
rect 16302 5264 16358 5273
rect 16396 5238 16448 5244
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 16946 5264 17002 5273
rect 16302 5199 16358 5208
rect 16316 4282 16344 5199
rect 16592 5030 16620 5238
rect 16946 5199 17002 5208
rect 16960 5166 16988 5199
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 16408 4146 16436 4966
rect 16776 4826 16804 5102
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16868 4622 16896 4966
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16960 4282 16988 4422
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16868 3738 16896 4218
rect 16946 4176 17002 4185
rect 16946 4111 16948 4120
rect 17000 4111 17002 4120
rect 16948 4082 17000 4088
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 16868 3466 16896 3674
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16408 3194 16436 3334
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 16488 3052 16540 3058
rect 16960 3040 16988 3946
rect 17052 3534 17080 5902
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17144 5302 17172 5714
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17144 3670 17172 5238
rect 17236 4146 17264 6258
rect 17328 6254 17356 6559
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17328 5574 17356 6054
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 17314 5128 17370 5137
rect 17314 5063 17370 5072
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17236 3602 17264 3878
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17040 3052 17092 3058
rect 16960 3012 17040 3040
rect 16488 2994 16540 3000
rect 17040 2994 17092 3000
rect 16500 2922 16528 2994
rect 17236 2961 17264 3538
rect 17328 3534 17356 5063
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17420 3097 17448 7103
rect 17512 7002 17540 7500
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17512 6361 17540 6734
rect 17498 6352 17554 6361
rect 17498 6287 17554 6296
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17512 5642 17540 6190
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 17406 3088 17462 3097
rect 17406 3023 17462 3032
rect 17512 3040 17540 5578
rect 17604 5370 17632 7958
rect 17696 7546 17724 8230
rect 17788 7993 17816 9302
rect 18064 9217 18092 10746
rect 18050 9208 18106 9217
rect 18050 9143 18106 9152
rect 18052 9104 18104 9110
rect 17866 9072 17922 9081
rect 18052 9046 18104 9052
rect 17866 9007 17922 9016
rect 17774 7984 17830 7993
rect 17774 7919 17830 7928
rect 17776 7880 17828 7886
rect 17774 7848 17776 7857
rect 17828 7848 17830 7857
rect 17774 7783 17830 7792
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17682 6896 17738 6905
rect 17682 6831 17738 6840
rect 17696 6730 17724 6831
rect 17880 6746 17908 9007
rect 17958 8664 18014 8673
rect 17958 8599 18014 8608
rect 17972 8566 18000 8599
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 17958 7984 18014 7993
rect 17958 7919 18014 7928
rect 17972 7721 18000 7919
rect 17958 7712 18014 7721
rect 17958 7647 18014 7656
rect 17684 6724 17736 6730
rect 17880 6718 18000 6746
rect 17684 6666 17736 6672
rect 17696 6497 17724 6666
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17682 6488 17738 6497
rect 17682 6423 17738 6432
rect 17684 6316 17736 6322
rect 17788 6304 17816 6598
rect 17736 6276 17816 6304
rect 17684 6258 17736 6264
rect 17880 6202 17908 6598
rect 17788 6174 17908 6202
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17696 5914 17724 6054
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17788 5778 17816 6174
rect 17972 6066 18000 6718
rect 18064 6322 18092 9046
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18156 8634 18184 8774
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18156 6497 18184 6802
rect 18142 6488 18198 6497
rect 18142 6423 18198 6432
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17880 6038 18000 6066
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17590 4992 17646 5001
rect 17590 4927 17646 4936
rect 17604 4282 17632 4927
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17592 3052 17644 3058
rect 17512 3012 17592 3040
rect 17592 2994 17644 3000
rect 17408 2984 17460 2990
rect 17222 2952 17278 2961
rect 16488 2916 16540 2922
rect 17406 2952 17408 2961
rect 17460 2952 17462 2961
rect 17222 2887 17278 2896
rect 17316 2916 17368 2922
rect 16488 2858 16540 2864
rect 17406 2887 17462 2896
rect 17316 2858 17368 2864
rect 16396 2848 16448 2854
rect 15936 2790 15988 2796
rect 16118 2816 16174 2825
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15752 1896 15804 1902
rect 15752 1838 15804 1844
rect 15660 1828 15712 1834
rect 15660 1770 15712 1776
rect 15568 1284 15620 1290
rect 15568 1226 15620 1232
rect 15856 800 15884 2586
rect 15948 2446 15976 2790
rect 16396 2790 16448 2796
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 16118 2751 16174 2760
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 16224 800 16252 2518
rect 16408 2446 16436 2790
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 16316 2106 16344 2382
rect 16776 2310 16804 2586
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16304 2100 16356 2106
rect 16304 2042 16356 2048
rect 16580 1420 16632 1426
rect 16580 1362 16632 1368
rect 16592 800 16620 1362
rect 16960 800 16988 2518
rect 17144 2514 17172 2790
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 17328 2446 17356 2858
rect 17696 2446 17724 5646
rect 17880 5352 17908 6038
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17788 5324 17908 5352
rect 17788 4010 17816 5324
rect 17972 5302 18000 5714
rect 18064 5710 18092 6258
rect 18156 6254 18184 6423
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18156 5846 18184 6190
rect 18144 5840 18196 5846
rect 18144 5782 18196 5788
rect 18052 5704 18104 5710
rect 18248 5658 18276 10950
rect 18340 10606 18368 11070
rect 18432 10810 18460 12038
rect 18524 11014 18552 14282
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18420 10804 18472 10810
rect 18616 10792 18644 14894
rect 18708 11257 18736 19314
rect 18892 19242 18920 20266
rect 18984 20058 19012 22200
rect 19062 21856 19118 21865
rect 19062 21791 19118 21800
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 18984 19514 19012 19722
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18970 19408 19026 19417
rect 18970 19343 19026 19352
rect 18880 19236 18932 19242
rect 18880 19178 18932 19184
rect 18984 19122 19012 19343
rect 18892 19094 19012 19122
rect 18892 18766 18920 19094
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18892 17746 18920 18702
rect 19076 17882 19104 21791
rect 19352 20346 19380 22200
rect 19522 21448 19578 21457
rect 19522 21383 19578 21392
rect 19536 20602 19564 21383
rect 19524 20596 19576 20602
rect 19720 20584 19748 22200
rect 19984 20596 20036 20602
rect 19720 20556 19932 20584
rect 19524 20538 19576 20544
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19352 20318 19564 20346
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 19260 19378 19288 19926
rect 19352 19378 19380 19994
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 19444 19417 19472 19450
rect 19430 19408 19486 19417
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19340 19372 19392 19378
rect 19536 19378 19564 20318
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19628 19922 19656 20266
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 19430 19343 19486 19352
rect 19524 19372 19576 19378
rect 19340 19314 19392 19320
rect 19524 19314 19576 19320
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19432 18896 19484 18902
rect 19430 18864 19432 18873
rect 19484 18864 19486 18873
rect 19340 18828 19392 18834
rect 19430 18799 19486 18808
rect 19340 18770 19392 18776
rect 19352 18737 19380 18770
rect 19432 18760 19484 18766
rect 19338 18728 19394 18737
rect 19432 18702 19484 18708
rect 19338 18663 19394 18672
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19352 18222 19380 18566
rect 19444 18465 19472 18702
rect 19536 18630 19564 19314
rect 19628 18970 19656 19722
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19628 18737 19656 18906
rect 19720 18902 19748 20402
rect 19904 19938 19932 20556
rect 19984 20538 20036 20544
rect 19996 20505 20024 20538
rect 19982 20496 20038 20505
rect 19982 20431 20038 20440
rect 20088 19938 20116 22200
rect 20352 20596 20404 20602
rect 20352 20538 20404 20544
rect 20364 20233 20392 20538
rect 20350 20224 20406 20233
rect 20350 20159 20406 20168
rect 19904 19910 20024 19938
rect 20088 19910 20208 19938
rect 20456 19922 20484 22200
rect 20626 22128 20682 22137
rect 20626 22063 20682 22072
rect 20534 21040 20590 21049
rect 20534 20975 20590 20984
rect 20548 20058 20576 20975
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20640 19938 20668 22063
rect 20824 20369 20852 22200
rect 21192 20602 21220 22200
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 20810 20360 20866 20369
rect 20810 20295 20866 20304
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19812 19009 19840 19790
rect 19892 19780 19944 19786
rect 19892 19722 19944 19728
rect 19904 19417 19932 19722
rect 19996 19553 20024 19910
rect 20076 19780 20128 19786
rect 20076 19722 20128 19728
rect 19982 19544 20038 19553
rect 19982 19479 20038 19488
rect 19890 19408 19946 19417
rect 19890 19343 19946 19352
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19798 19000 19854 19009
rect 19798 18935 19854 18944
rect 19708 18896 19760 18902
rect 19708 18838 19760 18844
rect 19614 18728 19670 18737
rect 19614 18663 19670 18672
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19904 18465 19932 19110
rect 19430 18456 19486 18465
rect 19890 18456 19946 18465
rect 19430 18391 19486 18400
rect 19524 18420 19576 18426
rect 19576 18380 19748 18408
rect 19890 18391 19946 18400
rect 19524 18362 19576 18368
rect 19720 18290 19748 18380
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19614 18184 19670 18193
rect 19614 18119 19670 18128
rect 19628 18086 19656 18119
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19064 17876 19116 17882
rect 19064 17818 19116 17824
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 19524 17604 19576 17610
rect 19524 17546 19576 17552
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18800 16250 18828 16730
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 19076 15688 19104 15982
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19432 15700 19484 15706
rect 19076 15660 19288 15688
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18800 14006 18828 15302
rect 19076 14550 19104 15660
rect 19260 15570 19288 15660
rect 19432 15642 19484 15648
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19444 15502 19472 15642
rect 19536 15502 19564 17546
rect 19628 16561 19656 18022
rect 19720 17814 19748 18226
rect 19996 18086 20024 19314
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19708 17808 19760 17814
rect 19708 17750 19760 17756
rect 20088 17678 20116 19722
rect 20180 19174 20208 19910
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 20548 19910 20668 19938
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20260 19236 20312 19242
rect 20260 19178 20312 19184
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20272 18986 20300 19178
rect 20180 18958 20300 18986
rect 20180 18873 20208 18958
rect 20364 18873 20392 19790
rect 20456 19378 20484 19858
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 20442 19272 20498 19281
rect 20548 19242 20576 19910
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20442 19207 20498 19216
rect 20536 19236 20588 19242
rect 20166 18864 20222 18873
rect 20166 18799 20222 18808
rect 20350 18864 20406 18873
rect 20350 18799 20406 18808
rect 20180 18290 20208 18799
rect 20456 18766 20484 19207
rect 20536 19178 20588 19184
rect 20534 19000 20590 19009
rect 20534 18935 20590 18944
rect 20548 18902 20576 18935
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 20640 18766 20668 19314
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20444 18760 20496 18766
rect 20350 18728 20406 18737
rect 20260 18692 20312 18698
rect 20444 18702 20496 18708
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20350 18663 20406 18672
rect 20260 18634 20312 18640
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20168 18080 20220 18086
rect 20166 18048 20168 18057
rect 20220 18048 20222 18057
rect 20166 17983 20222 17992
rect 19708 17672 19760 17678
rect 19708 17614 19760 17620
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19720 17270 19748 17614
rect 20272 17338 20300 18634
rect 20364 18630 20392 18663
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20364 18193 20392 18226
rect 20456 18222 20484 18702
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20444 18216 20496 18222
rect 20350 18184 20406 18193
rect 20444 18158 20496 18164
rect 20350 18119 20406 18128
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 19708 17264 19760 17270
rect 19708 17206 19760 17212
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19812 16794 19840 17138
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19904 16574 19932 16934
rect 20364 16697 20392 17478
rect 20548 17338 20576 18226
rect 20640 18154 20668 18702
rect 20824 18358 20852 19246
rect 21008 18970 21036 20402
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 21100 19825 21128 20198
rect 21272 19848 21324 19854
rect 21086 19816 21142 19825
rect 21272 19790 21324 19796
rect 21086 19751 21142 19760
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20628 18148 20680 18154
rect 20628 18090 20680 18096
rect 20732 17338 20760 18226
rect 20810 17776 20866 17785
rect 20810 17711 20866 17720
rect 20536 17332 20588 17338
rect 20536 17274 20588 17280
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20824 17202 20852 17711
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20350 16688 20406 16697
rect 20168 16652 20220 16658
rect 20350 16623 20406 16632
rect 20168 16594 20220 16600
rect 19614 16552 19670 16561
rect 19614 16487 19670 16496
rect 19812 16546 19932 16574
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19444 14804 19472 15438
rect 19536 15162 19564 15438
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19444 14776 19564 14804
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19536 14618 19564 14776
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19064 14544 19116 14550
rect 19064 14486 19116 14492
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 18892 13818 18920 14214
rect 19536 14113 19564 14554
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19522 14104 19578 14113
rect 19522 14039 19578 14048
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 18800 13790 18920 13818
rect 18972 13796 19024 13802
rect 18800 13190 18828 13790
rect 18972 13738 19024 13744
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18892 13394 18920 13670
rect 18984 13530 19012 13738
rect 19076 13530 19104 13874
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 18880 13388 18932 13394
rect 18880 13330 18932 13336
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18892 12850 18920 13330
rect 18984 12918 19012 13466
rect 19536 12986 19564 13874
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18970 12744 19026 12753
rect 18970 12679 19026 12688
rect 19524 12708 19576 12714
rect 18984 12434 19012 12679
rect 19524 12650 19576 12656
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 18984 12406 19196 12434
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18788 11824 18840 11830
rect 18788 11766 18840 11772
rect 18800 11354 18828 11766
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18694 11248 18750 11257
rect 18694 11183 18750 11192
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18420 10746 18472 10752
rect 18524 10764 18644 10792
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18326 9208 18382 9217
rect 18326 9143 18382 9152
rect 18340 6225 18368 9143
rect 18524 7970 18552 10764
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18432 7942 18552 7970
rect 18326 6216 18382 6225
rect 18326 6151 18382 6160
rect 18328 6112 18380 6118
rect 18326 6080 18328 6089
rect 18380 6080 18382 6089
rect 18326 6015 18382 6024
rect 18326 5944 18382 5953
rect 18326 5879 18382 5888
rect 18340 5846 18368 5879
rect 18328 5840 18380 5846
rect 18328 5782 18380 5788
rect 18052 5646 18104 5652
rect 18156 5630 18276 5658
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17880 4826 17908 5170
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17972 4078 18000 4558
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 18064 4010 18092 5510
rect 18156 4282 18184 5630
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18248 4010 18276 5510
rect 18340 5166 18368 5646
rect 18432 5545 18460 7942
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18524 7274 18552 7754
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 18512 6928 18564 6934
rect 18512 6870 18564 6876
rect 18524 6633 18552 6870
rect 18510 6624 18566 6633
rect 18510 6559 18566 6568
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18524 6361 18552 6394
rect 18510 6352 18566 6361
rect 18510 6287 18566 6296
rect 18616 6118 18644 10610
rect 18708 10266 18736 11018
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18694 10024 18750 10033
rect 18694 9959 18750 9968
rect 18708 7818 18736 9959
rect 18800 9897 18828 10542
rect 18786 9888 18842 9897
rect 18786 9823 18842 9832
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18800 8129 18828 9318
rect 18892 9178 18920 12174
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18984 11132 19012 11494
rect 19076 11286 19104 11698
rect 19168 11558 19196 12406
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19352 11830 19380 12038
rect 19340 11824 19392 11830
rect 19340 11766 19392 11772
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 18984 11104 19104 11132
rect 18970 10704 19026 10713
rect 18970 10639 18972 10648
rect 19024 10639 19026 10648
rect 18972 10610 19024 10616
rect 18972 9988 19024 9994
rect 18972 9930 19024 9936
rect 18984 9625 19012 9930
rect 18970 9616 19026 9625
rect 18970 9551 19026 9560
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 19076 8974 19104 11104
rect 19260 10606 19288 11222
rect 19248 10600 19300 10606
rect 19248 10542 19300 10548
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19168 9722 19196 9862
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 19352 9586 19380 10134
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19444 9489 19472 9522
rect 19430 9480 19486 9489
rect 19430 9415 19486 9424
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19536 8974 19564 12650
rect 19628 10266 19656 14214
rect 19720 13530 19748 14962
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19708 13320 19760 13326
rect 19706 13288 19708 13297
rect 19760 13288 19762 13297
rect 19706 13223 19762 13232
rect 19812 11014 19840 16546
rect 20076 16516 20128 16522
rect 20076 16458 20128 16464
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19996 15094 20024 16390
rect 20088 15502 20116 16458
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 20180 15042 20208 16594
rect 20350 16552 20406 16561
rect 20350 16487 20406 16496
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20272 15162 20300 16050
rect 20364 15314 20392 16487
rect 20456 16250 20484 17070
rect 20548 16998 20576 17138
rect 20824 17066 20852 17138
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20812 17060 20864 17066
rect 20812 17002 20864 17008
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20548 15706 20576 16050
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20364 15286 20484 15314
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20180 15014 20300 15042
rect 20076 14340 20128 14346
rect 20076 14282 20128 14288
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19904 13326 19932 13670
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19904 10810 19932 12038
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19628 9450 19656 10066
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19720 9586 19748 9998
rect 19812 9722 19840 10610
rect 19892 10260 19944 10266
rect 19892 10202 19944 10208
rect 19800 9716 19852 9722
rect 19800 9658 19852 9664
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19616 9444 19668 9450
rect 19812 9432 19840 9522
rect 19616 9386 19668 9392
rect 19720 9404 19840 9432
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 18786 8120 18842 8129
rect 18892 8090 18920 8910
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 18786 8055 18842 8064
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18984 8022 19012 8502
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18800 6798 18828 7686
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18892 7002 18920 7278
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 18878 6896 18934 6905
rect 18878 6831 18934 6840
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18786 6352 18842 6361
rect 18786 6287 18788 6296
rect 18840 6287 18842 6296
rect 18788 6258 18840 6264
rect 18694 6216 18750 6225
rect 18694 6151 18750 6160
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18512 5568 18564 5574
rect 18418 5536 18474 5545
rect 18512 5510 18564 5516
rect 18418 5471 18474 5480
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18432 4758 18460 5170
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 17776 4004 17828 4010
rect 17776 3946 17828 3952
rect 18052 4004 18104 4010
rect 18052 3946 18104 3952
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18050 3088 18106 3097
rect 18050 3023 18052 3032
rect 18104 3023 18106 3032
rect 18052 2994 18104 3000
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17604 1426 17632 2246
rect 17592 1420 17644 1426
rect 17592 1362 17644 1368
rect 17696 1170 17724 2246
rect 17604 1142 17724 1170
rect 17328 870 17448 898
rect 17328 800 17356 870
rect 11900 734 12112 762
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17420 762 17448 870
rect 17604 762 17632 1142
rect 17788 898 17816 2586
rect 17696 870 17816 898
rect 17696 800 17724 870
rect 18064 800 18092 2858
rect 18156 2446 18184 3130
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 18248 2446 18276 2790
rect 18340 2514 18368 4558
rect 18524 4554 18552 5510
rect 18512 4548 18564 4554
rect 18512 4490 18564 4496
rect 18510 4448 18566 4457
rect 18510 4383 18566 4392
rect 18524 3058 18552 4383
rect 18616 3670 18644 6054
rect 18708 4622 18736 6151
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18800 4570 18828 6258
rect 18892 6168 18920 6831
rect 18984 6458 19012 7346
rect 19076 6798 19104 8910
rect 19352 8838 19380 8910
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19154 8664 19210 8673
rect 19444 8634 19472 8842
rect 19720 8634 19748 9404
rect 19904 9330 19932 10202
rect 19812 9302 19932 9330
rect 19154 8599 19210 8608
rect 19432 8628 19484 8634
rect 19168 8566 19196 8599
rect 19432 8570 19484 8576
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19156 8560 19208 8566
rect 19156 8502 19208 8508
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19340 8424 19392 8430
rect 19338 8392 19340 8401
rect 19392 8392 19394 8401
rect 19338 8327 19394 8336
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19628 7857 19656 8434
rect 19614 7848 19670 7857
rect 19614 7783 19670 7792
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 7546 19380 7686
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19260 6820 19380 6848
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 19076 6390 19104 6734
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 19168 6497 19196 6666
rect 19260 6633 19288 6820
rect 19246 6624 19302 6633
rect 19246 6559 19302 6568
rect 19154 6488 19210 6497
rect 19154 6423 19210 6432
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 19352 6322 19380 6820
rect 19432 6724 19484 6730
rect 19432 6666 19484 6672
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19444 6254 19472 6666
rect 19536 6458 19564 7414
rect 19628 7177 19656 7783
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19720 7546 19748 7686
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19614 7168 19670 7177
rect 19614 7103 19670 7112
rect 19812 6848 19840 9302
rect 19892 8492 19944 8498
rect 19892 8434 19944 8440
rect 19904 7993 19932 8434
rect 19890 7984 19946 7993
rect 19890 7919 19946 7928
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19628 6820 19840 6848
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19064 6180 19116 6186
rect 18892 6140 19012 6168
rect 18878 6080 18934 6089
rect 18878 6015 18934 6024
rect 18892 5710 18920 6015
rect 18984 5914 19012 6140
rect 19064 6122 19116 6128
rect 18972 5908 19024 5914
rect 18972 5850 19024 5856
rect 19076 5846 19104 6122
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19064 5840 19116 5846
rect 18970 5808 19026 5817
rect 19064 5782 19116 5788
rect 18970 5743 19026 5752
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18984 5642 19012 5743
rect 18972 5636 19024 5642
rect 18972 5578 19024 5584
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19536 4622 19564 4966
rect 19524 4616 19576 4622
rect 18800 4542 18920 4570
rect 19524 4558 19576 4564
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18708 3738 18736 4422
rect 18800 3738 18828 4422
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18892 3670 18920 4542
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18984 3913 19012 4082
rect 19430 4040 19486 4049
rect 19430 3975 19486 3984
rect 19444 3942 19472 3975
rect 19432 3936 19484 3942
rect 18970 3904 19026 3913
rect 19432 3878 19484 3884
rect 18970 3839 19026 3848
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 18984 3505 19012 3839
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 18970 3496 19026 3505
rect 18970 3431 19026 3440
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 19168 3058 19196 3402
rect 19260 3194 19288 3538
rect 19628 3534 19656 6820
rect 19800 6724 19852 6730
rect 19800 6666 19852 6672
rect 19812 5681 19840 6666
rect 19904 6186 19932 7278
rect 19892 6180 19944 6186
rect 19892 6122 19944 6128
rect 19798 5672 19854 5681
rect 19708 5636 19760 5642
rect 19798 5607 19854 5616
rect 19708 5578 19760 5584
rect 19720 5030 19748 5578
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 19720 4690 19748 4966
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 19812 4298 19840 5607
rect 19720 4270 19840 4298
rect 19720 4010 19748 4270
rect 19996 4146 20024 14214
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 19708 4004 19760 4010
rect 19708 3946 19760 3952
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19628 3210 19656 3470
rect 19248 3188 19300 3194
rect 19628 3182 19748 3210
rect 19248 3130 19300 3136
rect 19720 3097 19748 3182
rect 19706 3088 19762 3097
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 19616 3052 19668 3058
rect 19706 3023 19762 3032
rect 19616 2994 19668 3000
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 18432 800 18460 2518
rect 18800 800 18828 2790
rect 18984 2446 19012 2926
rect 19156 2848 19208 2854
rect 19076 2808 19156 2836
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 19076 1442 19104 2808
rect 19156 2790 19208 2796
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 19168 2038 19196 2450
rect 19156 2032 19208 2038
rect 19156 1974 19208 1980
rect 19076 1414 19196 1442
rect 19168 800 19196 1414
rect 19536 800 19564 2790
rect 19628 2650 19656 2994
rect 19706 2952 19762 2961
rect 19706 2887 19762 2896
rect 19720 2650 19748 2887
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 19812 1970 19840 4082
rect 19890 3768 19946 3777
rect 19890 3703 19892 3712
rect 19944 3703 19946 3712
rect 19892 3674 19944 3680
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19800 1964 19852 1970
rect 19800 1906 19852 1912
rect 19812 1873 19840 1906
rect 19798 1864 19854 1873
rect 19798 1799 19854 1808
rect 19904 800 19932 3470
rect 19996 2774 20024 4082
rect 20088 3534 20116 14282
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20180 12986 20208 13806
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20272 12374 20300 15014
rect 20352 13864 20404 13870
rect 20350 13832 20352 13841
rect 20404 13832 20406 13841
rect 20350 13767 20406 13776
rect 20456 12986 20484 15286
rect 20640 13569 20668 17002
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20732 16250 20760 16458
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20732 14618 20760 14962
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20810 13968 20866 13977
rect 20720 13932 20772 13938
rect 20810 13903 20866 13912
rect 20720 13874 20772 13880
rect 20626 13560 20682 13569
rect 20626 13495 20682 13504
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20548 12714 20576 13330
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 20536 12708 20588 12714
rect 20536 12650 20588 12656
rect 20444 12640 20496 12646
rect 20496 12588 20576 12594
rect 20444 12582 20576 12588
rect 20456 12566 20576 12582
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20180 10792 20208 12106
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20272 11762 20300 12038
rect 20364 11898 20392 12242
rect 20548 12238 20576 12566
rect 20640 12442 20668 13194
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20456 11898 20484 12106
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20364 11150 20392 11834
rect 20732 11665 20760 13874
rect 20824 12986 20852 13903
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 20824 12442 20852 12786
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20810 12336 20866 12345
rect 20810 12271 20866 12280
rect 20824 11694 20852 12271
rect 20812 11688 20864 11694
rect 20718 11656 20774 11665
rect 20812 11630 20864 11636
rect 20718 11591 20774 11600
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20352 11008 20404 11014
rect 20732 10985 20760 11086
rect 20812 11008 20864 11014
rect 20352 10950 20404 10956
rect 20718 10976 20774 10985
rect 20260 10804 20312 10810
rect 20180 10764 20260 10792
rect 20260 10746 20312 10752
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20180 9722 20208 10542
rect 20272 10266 20300 10542
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20364 10146 20392 10950
rect 20812 10950 20864 10956
rect 20718 10911 20774 10920
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20272 10118 20392 10146
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20166 9616 20222 9625
rect 20166 9551 20222 9560
rect 20180 8090 20208 9551
rect 20272 9518 20300 10118
rect 20456 9994 20484 10134
rect 20640 10062 20668 10406
rect 20628 10056 20680 10062
rect 20626 10024 20628 10033
rect 20680 10024 20682 10033
rect 20352 9988 20404 9994
rect 20352 9930 20404 9936
rect 20444 9988 20496 9994
rect 20626 9959 20682 9968
rect 20444 9930 20496 9936
rect 20260 9512 20312 9518
rect 20260 9454 20312 9460
rect 20258 9344 20314 9353
rect 20258 9279 20314 9288
rect 20272 8378 20300 9279
rect 20364 8634 20392 9930
rect 20456 9654 20484 9930
rect 20534 9888 20590 9897
rect 20534 9823 20590 9832
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20456 8430 20484 9454
rect 20548 8922 20576 9823
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20640 9042 20668 9386
rect 20732 9178 20760 10678
rect 20824 10130 20852 10950
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20718 9072 20774 9081
rect 20628 9036 20680 9042
rect 20718 9007 20774 9016
rect 20628 8978 20680 8984
rect 20548 8894 20668 8922
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20444 8424 20496 8430
rect 20350 8392 20406 8401
rect 20272 8350 20350 8378
rect 20444 8366 20496 8372
rect 20350 8327 20406 8336
rect 20258 8256 20314 8265
rect 20258 8191 20314 8200
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20272 8022 20300 8191
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 20180 7041 20208 7890
rect 20364 7546 20392 8327
rect 20456 8022 20484 8366
rect 20444 8016 20496 8022
rect 20444 7958 20496 7964
rect 20444 7880 20496 7886
rect 20442 7848 20444 7857
rect 20496 7848 20498 7857
rect 20442 7783 20498 7792
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20166 7032 20222 7041
rect 20166 6967 20222 6976
rect 20180 6186 20208 6967
rect 20272 6798 20300 7210
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20272 6458 20300 6598
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20168 6180 20220 6186
rect 20168 6122 20220 6128
rect 20272 4298 20300 6394
rect 20364 5098 20392 7346
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20456 6322 20484 6598
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20456 5166 20484 6258
rect 20548 6254 20576 8774
rect 20640 7478 20668 8894
rect 20732 8634 20760 9007
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20732 7954 20760 8366
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20628 7472 20680 7478
rect 20628 7414 20680 7420
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20352 5092 20404 5098
rect 20352 5034 20404 5040
rect 20442 4720 20498 4729
rect 20442 4655 20498 4664
rect 20180 4270 20300 4298
rect 20456 4282 20484 4655
rect 20444 4276 20496 4282
rect 20180 4010 20208 4270
rect 20444 4218 20496 4224
rect 20536 4072 20588 4078
rect 20258 4040 20314 4049
rect 20168 4004 20220 4010
rect 20258 3975 20314 3984
rect 20456 4020 20536 4026
rect 20456 4014 20588 4020
rect 20456 3998 20576 4014
rect 20168 3946 20220 3952
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20180 3398 20208 3674
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 20272 3058 20300 3975
rect 20456 3942 20484 3998
rect 20444 3936 20496 3942
rect 20350 3904 20406 3913
rect 20640 3890 20668 7414
rect 20732 6254 20760 7890
rect 20824 7546 20852 9454
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20824 6390 20852 7346
rect 20812 6384 20864 6390
rect 20812 6326 20864 6332
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20824 5846 20852 6326
rect 20812 5840 20864 5846
rect 20812 5782 20864 5788
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20732 5370 20760 5510
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20732 4146 20760 4422
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20444 3878 20496 3884
rect 20350 3839 20406 3848
rect 20548 3862 20668 3890
rect 20364 3058 20392 3839
rect 20548 3738 20576 3862
rect 20626 3768 20682 3777
rect 20536 3732 20588 3738
rect 20626 3703 20682 3712
rect 20720 3732 20772 3738
rect 20536 3674 20588 3680
rect 20640 3534 20668 3703
rect 20720 3674 20772 3680
rect 20732 3534 20760 3674
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 19996 2746 20116 2774
rect 20088 2689 20116 2746
rect 20074 2680 20130 2689
rect 20074 2615 20130 2624
rect 20272 800 20300 2790
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 20548 1329 20576 2382
rect 20534 1320 20590 1329
rect 20534 1255 20590 1264
rect 20548 1057 20576 1255
rect 20534 1048 20590 1057
rect 20534 983 20590 992
rect 20640 800 20668 2858
rect 20732 2774 20760 3470
rect 20824 2990 20852 5646
rect 20916 3602 20944 18634
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21008 17338 21036 18226
rect 21086 18184 21142 18193
rect 21086 18119 21088 18128
rect 21140 18119 21142 18128
rect 21088 18090 21140 18096
rect 21192 18086 21220 19314
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21284 17882 21312 19790
rect 21376 18222 21404 20334
rect 21560 20330 21588 22200
rect 21548 20324 21600 20330
rect 21548 20266 21600 20272
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21468 19417 21496 19654
rect 21454 19408 21510 19417
rect 21454 19343 21510 19352
rect 21456 19168 21508 19174
rect 21456 19110 21508 19116
rect 21468 19009 21496 19110
rect 21454 19000 21510 19009
rect 21454 18935 21510 18944
rect 21454 18728 21510 18737
rect 21454 18663 21510 18672
rect 21468 18630 21496 18663
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21652 18426 21680 22222
rect 21836 22114 21864 22222
rect 21914 22200 21970 23000
rect 22282 22200 22338 23000
rect 21928 22114 21956 22200
rect 21836 22086 21956 22114
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 22296 19514 22324 22200
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 21364 18216 21416 18222
rect 21364 18158 21416 18164
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 21468 17785 21496 18022
rect 22100 17808 22152 17814
rect 21454 17776 21510 17785
rect 22100 17750 22152 17756
rect 21454 17711 21510 17720
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 21284 16794 21312 17614
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21468 17241 21496 17478
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21454 17232 21510 17241
rect 21454 17167 21510 17176
rect 21456 16992 21508 16998
rect 21454 16960 21456 16969
rect 21508 16960 21510 16969
rect 21454 16895 21510 16904
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 21086 16552 21142 16561
rect 21008 16250 21036 16526
rect 21086 16487 21142 16496
rect 21100 16454 21128 16487
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 21468 16153 21496 16390
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21454 16144 21510 16153
rect 21272 16108 21324 16114
rect 21454 16079 21510 16088
rect 21272 16050 21324 16056
rect 21284 15706 21312 16050
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21468 15745 21496 15846
rect 21454 15736 21510 15745
rect 21272 15700 21324 15706
rect 21454 15671 21510 15680
rect 21272 15642 21324 15648
rect 21454 15464 21510 15473
rect 21454 15399 21510 15408
rect 21468 15366 21496 15399
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21008 14618 21036 14962
rect 21086 14920 21142 14929
rect 21086 14855 21088 14864
rect 21140 14855 21142 14864
rect 21088 14826 21140 14832
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 21008 14074 21036 14350
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 21008 12986 21036 13874
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21100 12889 21128 13126
rect 21086 12880 21142 12889
rect 20996 12844 21048 12850
rect 21086 12815 21142 12824
rect 20996 12786 21048 12792
rect 21008 10130 21036 12786
rect 21088 12164 21140 12170
rect 21088 12106 21140 12112
rect 21100 11257 21128 12106
rect 21192 11336 21220 15302
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21272 13796 21324 13802
rect 21272 13738 21324 13744
rect 21284 13326 21312 13738
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21284 11830 21312 12786
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21376 11558 21404 14894
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 14521 21496 14758
rect 21454 14512 21510 14521
rect 21454 14447 21510 14456
rect 21456 14272 21508 14278
rect 21456 14214 21508 14220
rect 21468 13977 21496 14214
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21454 13968 21510 13977
rect 21454 13903 21510 13912
rect 21456 13728 21508 13734
rect 21454 13696 21456 13705
rect 21508 13696 21510 13705
rect 21454 13631 21510 13640
rect 21638 13424 21694 13433
rect 21638 13359 21694 13368
rect 21454 13288 21510 13297
rect 21454 13223 21510 13232
rect 21468 13190 21496 13223
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21468 12481 21496 12582
rect 21454 12472 21510 12481
rect 21454 12407 21510 12416
rect 21454 12200 21510 12209
rect 21454 12135 21510 12144
rect 21468 12102 21496 12135
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21560 11694 21588 12650
rect 21652 12434 21680 13359
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21652 12406 22048 12434
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 22020 12186 22048 12406
rect 22112 12306 22140 17750
rect 22836 17060 22888 17066
rect 22836 17002 22888 17008
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 22204 12322 22232 15030
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 22296 12442 22324 14826
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22560 12368 22612 12374
rect 22100 12300 22152 12306
rect 22204 12294 22324 12322
rect 22560 12310 22612 12316
rect 22100 12242 22152 12248
rect 21548 11688 21600 11694
rect 21546 11656 21548 11665
rect 21600 11656 21602 11665
rect 21546 11591 21602 11600
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21192 11308 21588 11336
rect 21086 11248 21142 11257
rect 21086 11183 21142 11192
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21178 10840 21234 10849
rect 21178 10775 21234 10784
rect 21192 10742 21220 10775
rect 21180 10736 21232 10742
rect 21086 10704 21142 10713
rect 21180 10678 21232 10684
rect 21086 10639 21088 10648
rect 21140 10639 21142 10648
rect 21088 10610 21140 10616
rect 21178 10432 21234 10441
rect 21178 10367 21234 10376
rect 20996 10124 21048 10130
rect 20996 10066 21048 10072
rect 21192 9738 21220 10367
rect 21284 10198 21312 11154
rect 21454 10704 21510 10713
rect 21454 10639 21456 10648
rect 21508 10639 21510 10648
rect 21456 10610 21508 10616
rect 21272 10192 21324 10198
rect 21324 10152 21404 10180
rect 21272 10134 21324 10140
rect 21270 9752 21326 9761
rect 21192 9710 21270 9738
rect 21270 9687 21326 9696
rect 21284 9654 21312 9687
rect 20996 9648 21048 9654
rect 20996 9590 21048 9596
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21008 7478 21036 9590
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 21100 8945 21128 9386
rect 21086 8936 21142 8945
rect 21086 8871 21142 8880
rect 21270 8936 21326 8945
rect 21270 8871 21326 8880
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21100 8090 21128 8774
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 20994 7304 21050 7313
rect 20994 7239 21050 7248
rect 21008 6866 21036 7239
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 21100 5914 21128 7142
rect 21192 6458 21220 8774
rect 21284 8566 21312 8871
rect 21272 8560 21324 8566
rect 21272 8502 21324 8508
rect 21376 8430 21404 10152
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21284 7002 21312 7686
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 21008 4214 21036 5646
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 21100 5137 21128 5510
rect 21086 5128 21142 5137
rect 21086 5063 21142 5072
rect 21086 4720 21142 4729
rect 21086 4655 21142 4664
rect 21100 4214 21128 4655
rect 21284 4486 21312 6938
rect 21376 6769 21404 8230
rect 21468 8090 21496 10610
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21362 6760 21418 6769
rect 21362 6695 21418 6704
rect 21468 6644 21496 7890
rect 21376 6616 21496 6644
rect 21376 4622 21404 6616
rect 21454 5536 21510 5545
rect 21454 5471 21510 5480
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 21468 4214 21496 5471
rect 21560 5234 21588 11308
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21560 5137 21588 5170
rect 21546 5128 21602 5137
rect 21546 5063 21602 5072
rect 21652 4826 21680 12174
rect 22020 12158 22232 12186
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 22006 9208 22062 9217
rect 22006 9143 22062 9152
rect 22020 8838 22048 9143
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21730 8528 21786 8537
rect 21730 8463 21786 8472
rect 21744 7954 21772 8463
rect 21732 7948 21784 7954
rect 21732 7890 21784 7896
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21914 7440 21970 7449
rect 21914 7375 21970 7384
rect 21928 6644 21956 7375
rect 22112 6798 22140 11494
rect 22100 6792 22152 6798
rect 22006 6760 22062 6769
rect 22062 6740 22100 6746
rect 22062 6734 22152 6740
rect 22062 6718 22140 6734
rect 22006 6695 22062 6704
rect 21928 6616 22140 6644
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 22112 5166 22140 6616
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 21640 4820 21692 4826
rect 21640 4762 21692 4768
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 20996 4208 21048 4214
rect 20996 4150 21048 4156
rect 21088 4208 21140 4214
rect 21088 4150 21140 4156
rect 21456 4208 21508 4214
rect 22008 4208 22060 4214
rect 21456 4150 21508 4156
rect 22006 4176 22008 4185
rect 22060 4176 22062 4185
rect 22006 4111 22062 4120
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 21364 3936 21416 3942
rect 22020 3913 22048 4014
rect 22204 4010 22232 12158
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 21364 3878 21416 3884
rect 22006 3904 22062 3913
rect 20996 3664 21048 3670
rect 21376 3641 21404 3878
rect 22296 3890 22324 12294
rect 22376 12300 22428 12306
rect 22376 12242 22428 12248
rect 22062 3862 22324 3890
rect 22006 3839 22062 3848
rect 22006 3768 22062 3777
rect 22388 3754 22416 12242
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22480 6730 22508 7890
rect 22468 6724 22520 6730
rect 22468 6666 22520 6672
rect 22572 4690 22600 12310
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22572 4214 22600 4626
rect 22560 4208 22612 4214
rect 22560 4150 22612 4156
rect 22062 3726 22416 3754
rect 22664 3738 22692 15098
rect 22848 11898 22876 17002
rect 22928 14340 22980 14346
rect 22928 14282 22980 14288
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22836 11620 22888 11626
rect 22836 11562 22888 11568
rect 22652 3732 22704 3738
rect 22006 3703 22062 3712
rect 22652 3674 22704 3680
rect 20996 3606 21048 3612
rect 21362 3632 21418 3641
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20732 2746 20852 2774
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 20732 2417 20760 2450
rect 20718 2408 20774 2417
rect 20718 2343 20774 2352
rect 20824 1465 20852 2746
rect 20916 2514 20944 3402
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 20810 1456 20866 1465
rect 20810 1391 20866 1400
rect 21008 800 21036 3606
rect 21362 3567 21418 3576
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 21100 3194 21128 3470
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 21376 800 21404 3334
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 22756 3058 22784 11562
rect 22848 7954 22876 11562
rect 22836 7948 22888 7954
rect 22836 7890 22888 7896
rect 22836 7812 22888 7818
rect 22836 7754 22888 7760
rect 21640 3052 21692 3058
rect 21640 2994 21692 3000
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 17420 734 17632 762
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21652 649 21680 2994
rect 22848 2514 22876 7754
rect 22940 5642 22968 14282
rect 22928 5636 22980 5642
rect 22928 5578 22980 5584
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 21638 640 21694 649
rect 21638 575 21694 584
<< via2 >>
rect 18 22480 74 22536
rect 1582 22208 1638 22264
rect 938 14320 994 14376
rect 1490 20204 1492 20224
rect 1492 20204 1544 20224
rect 1544 20204 1546 20224
rect 1490 20168 1546 20204
rect 1122 16224 1178 16280
rect 938 7964 940 7984
rect 940 7964 992 7984
rect 992 7964 994 7984
rect 938 7928 994 7964
rect 938 6740 940 6760
rect 940 6740 992 6760
rect 992 6740 994 6760
rect 938 6704 994 6740
rect 1950 21392 2006 21448
rect 1858 20596 1914 20632
rect 1858 20576 1860 20596
rect 1860 20576 1912 20596
rect 1912 20576 1914 20596
rect 1490 19352 1546 19408
rect 1490 18944 1546 19000
rect 1858 19760 1914 19816
rect 1490 18128 1546 18184
rect 1490 17720 1546 17776
rect 1490 17312 1546 17368
rect 1490 16940 1492 16960
rect 1492 16940 1544 16960
rect 1544 16940 1546 16960
rect 1490 16904 1546 16940
rect 1490 16088 1546 16144
rect 1490 15680 1546 15736
rect 1950 19372 2006 19408
rect 1950 19352 1952 19372
rect 1952 19352 2004 19372
rect 2004 19352 2006 19372
rect 1950 18572 1952 18592
rect 1952 18572 2004 18592
rect 2004 18572 2006 18592
rect 1950 18536 2006 18572
rect 1858 16496 1914 16552
rect 2226 20984 2282 21040
rect 2410 20460 2466 20496
rect 2410 20440 2412 20460
rect 2412 20440 2464 20460
rect 2464 20440 2466 20460
rect 2410 19896 2466 19952
rect 2594 18808 2650 18864
rect 1490 15308 1492 15328
rect 1492 15308 1544 15328
rect 1544 15308 1546 15328
rect 1490 15272 1546 15308
rect 1858 14884 1914 14920
rect 1858 14864 1860 14884
rect 1860 14864 1912 14884
rect 1912 14864 1914 14884
rect 1490 14456 1546 14512
rect 1490 14048 1546 14104
rect 2042 14184 2098 14240
rect 1950 13912 2006 13968
rect 2226 17076 2228 17096
rect 2228 17076 2280 17096
rect 2280 17076 2282 17096
rect 2226 17040 2282 17076
rect 2594 17584 2650 17640
rect 2594 17312 2650 17368
rect 2502 16360 2558 16416
rect 2962 19624 3018 19680
rect 2962 19488 3018 19544
rect 3238 21256 3294 21312
rect 3330 20984 3386 21040
rect 3514 20304 3570 20360
rect 3238 19216 3294 19272
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 4158 21800 4214 21856
rect 3974 20168 4030 20224
rect 3606 19216 3662 19272
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3882 18808 3938 18864
rect 3422 18264 3478 18320
rect 4066 18672 4122 18728
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 2594 15952 2650 16008
rect 2318 15544 2374 15600
rect 3606 17584 3662 17640
rect 2594 15136 2650 15192
rect 3054 15308 3056 15328
rect 3056 15308 3108 15328
rect 3108 15308 3110 15328
rect 3054 15272 3110 15308
rect 3238 15000 3294 15056
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 1490 13676 1492 13696
rect 1492 13676 1544 13696
rect 1544 13676 1546 13696
rect 1490 13640 1546 13676
rect 1490 13232 1546 13288
rect 1858 12824 1914 12880
rect 1490 12436 1546 12472
rect 1490 12416 1492 12436
rect 1492 12416 1544 12436
rect 1544 12416 1546 12436
rect 1306 12280 1362 12336
rect 1214 9424 1270 9480
rect 1214 8336 1270 8392
rect 1030 6160 1086 6216
rect 1122 5888 1178 5944
rect 1214 5208 1270 5264
rect 1858 12044 1860 12064
rect 1860 12044 1912 12064
rect 1912 12044 1914 12064
rect 1858 12008 1914 12044
rect 1674 11328 1730 11384
rect 1490 11192 1546 11248
rect 2410 13096 2466 13152
rect 2318 12144 2374 12200
rect 2226 11636 2228 11656
rect 2228 11636 2280 11656
rect 2280 11636 2282 11656
rect 2226 11600 2282 11636
rect 2042 11328 2098 11384
rect 1858 10784 1914 10840
rect 1582 9968 1638 10024
rect 1490 9560 1546 9616
rect 2042 10648 2098 10704
rect 1950 10376 2006 10432
rect 1398 9152 1454 9208
rect 1398 8200 1454 8256
rect 1582 8628 1638 8664
rect 1582 8608 1584 8628
rect 1584 8608 1636 8628
rect 1636 8608 1638 8628
rect 1582 7792 1638 7848
rect 1674 7268 1730 7304
rect 1674 7248 1676 7268
rect 1676 7248 1728 7268
rect 1728 7248 1730 7268
rect 1398 7112 1454 7168
rect 1582 6840 1638 6896
rect 1490 5752 1546 5808
rect 1306 4800 1362 4856
rect 1490 3712 1546 3768
rect 1398 3168 1454 3224
rect 2042 6840 2098 6896
rect 2042 6432 2098 6488
rect 1950 5344 2006 5400
rect 1950 4936 2006 4992
rect 2502 8608 2558 8664
rect 2594 7656 2650 7712
rect 2870 8880 2926 8936
rect 3054 8744 3110 8800
rect 2870 8492 2926 8528
rect 2870 8472 2872 8492
rect 2872 8472 2924 8492
rect 2924 8472 2926 8492
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 4802 21120 4858 21176
rect 4250 17720 4306 17776
rect 4066 15408 4122 15464
rect 4158 15308 4160 15328
rect 4160 15308 4212 15328
rect 4212 15308 4214 15328
rect 4158 15272 4214 15308
rect 4066 13932 4122 13968
rect 4526 18400 4582 18456
rect 4526 17856 4582 17912
rect 4894 20848 4950 20904
rect 5078 19080 5134 19136
rect 4526 17584 4582 17640
rect 4526 15816 4582 15872
rect 4710 17720 4766 17776
rect 5078 17584 5134 17640
rect 5446 20168 5502 20224
rect 5354 19760 5410 19816
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 5998 19508 6054 19544
rect 5998 19488 6000 19508
rect 6000 19488 6052 19508
rect 6052 19488 6054 19508
rect 5906 19216 5962 19272
rect 5354 17720 5410 17776
rect 5170 17176 5226 17232
rect 5354 16632 5410 16688
rect 5722 17312 5778 17368
rect 5722 16904 5778 16960
rect 4526 15136 4582 15192
rect 4066 13912 4068 13932
rect 4068 13912 4120 13932
rect 4120 13912 4122 13932
rect 4158 13812 4160 13832
rect 4160 13812 4212 13832
rect 4212 13812 4214 13832
rect 4158 13776 4214 13812
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 4066 13096 4122 13152
rect 4618 13776 4674 13832
rect 4342 13096 4398 13152
rect 3698 12008 3754 12064
rect 4158 12824 4214 12880
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 4618 12688 4674 12744
rect 5078 16360 5134 16416
rect 5354 15428 5410 15464
rect 5354 15408 5356 15428
rect 5356 15408 5408 15428
rect 5408 15408 5410 15428
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 7010 20304 7066 20360
rect 6458 17720 6514 17776
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 5998 16224 6054 16280
rect 5998 15952 6054 16008
rect 5906 15544 5962 15600
rect 6642 15544 6698 15600
rect 5906 15136 5962 15192
rect 4710 12552 4766 12608
rect 4986 12588 4988 12608
rect 4988 12588 5040 12608
rect 5040 12588 5042 12608
rect 4986 12552 5042 12588
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3422 10104 3478 10160
rect 3606 10124 3662 10160
rect 3606 10104 3608 10124
rect 3608 10104 3660 10124
rect 3660 10104 3662 10124
rect 3422 9968 3478 10024
rect 3238 9424 3294 9480
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 4342 9560 4398 9616
rect 2870 7520 2926 7576
rect 3146 7520 3202 7576
rect 2686 6568 2742 6624
rect 3330 6840 3386 6896
rect 2226 5108 2228 5128
rect 2228 5108 2280 5128
rect 2280 5108 2282 5128
rect 2226 5072 2282 5108
rect 2226 4120 2282 4176
rect 2410 5072 2466 5128
rect 2410 4528 2466 4584
rect 2502 4392 2558 4448
rect 2594 3440 2650 3496
rect 2502 3168 2558 3224
rect 2226 2488 2282 2544
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3974 8200 4030 8256
rect 3698 7384 3754 7440
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3514 6840 3570 6896
rect 3514 6296 3570 6352
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3790 5652 3792 5672
rect 3792 5652 3844 5672
rect 3844 5652 3846 5672
rect 3790 5616 3846 5652
rect 3514 5480 3570 5536
rect 3422 5244 3424 5264
rect 3424 5244 3476 5264
rect 3476 5244 3478 5264
rect 3422 5208 3478 5244
rect 3974 7112 4030 7168
rect 4342 6976 4398 7032
rect 4250 6840 4306 6896
rect 4250 5752 4306 5808
rect 3790 5072 3846 5128
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3422 4256 3478 4312
rect 3330 3848 3386 3904
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 2870 2624 2926 2680
rect 2778 1128 2834 1184
rect 3146 3304 3202 3360
rect 3146 2508 3202 2544
rect 3146 2488 3148 2508
rect 3148 2488 3200 2508
rect 3200 2488 3202 2508
rect 3790 3032 3846 3088
rect 3330 2896 3386 2952
rect 3514 2896 3570 2952
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 3422 2352 3478 2408
rect 3698 2216 3754 2272
rect 3790 1808 3846 1864
rect 3974 1808 4030 1864
rect 4342 4800 4398 4856
rect 4250 4664 4306 4720
rect 4802 10240 4858 10296
rect 4894 8744 4950 8800
rect 4802 7656 4858 7712
rect 4710 6604 4712 6624
rect 4712 6604 4764 6624
rect 4764 6604 4766 6624
rect 4710 6568 4766 6604
rect 5722 15000 5778 15056
rect 5446 13132 5448 13152
rect 5448 13132 5500 13152
rect 5500 13132 5502 13152
rect 5446 13096 5502 13132
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 5262 12008 5318 12064
rect 5170 11056 5226 11112
rect 5078 9968 5134 10024
rect 6550 13640 6606 13696
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 5262 8916 5264 8936
rect 5264 8916 5316 8936
rect 5316 8916 5318 8936
rect 5262 8880 5318 8916
rect 5262 8744 5318 8800
rect 5538 9868 5540 9888
rect 5540 9868 5592 9888
rect 5592 9868 5594 9888
rect 5538 9832 5594 9868
rect 5538 9016 5594 9072
rect 5538 8472 5594 8528
rect 5078 7792 5134 7848
rect 4986 6704 5042 6760
rect 4986 6568 5042 6624
rect 4894 5888 4950 5944
rect 5262 6296 5318 6352
rect 5170 5752 5226 5808
rect 4802 4664 4858 4720
rect 4802 4428 4804 4448
rect 4804 4428 4856 4448
rect 4856 4428 4858 4448
rect 4802 4392 4858 4428
rect 4894 4256 4950 4312
rect 4526 2896 4582 2952
rect 4710 2624 4766 2680
rect 5262 4936 5318 4992
rect 5262 4664 5318 4720
rect 4986 2896 5042 2952
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 5906 11328 5962 11384
rect 6090 11328 6146 11384
rect 5906 11056 5962 11112
rect 6366 11736 6422 11792
rect 6642 13096 6698 13152
rect 7102 19488 7158 19544
rect 7010 19216 7066 19272
rect 7378 19080 7434 19136
rect 6918 14456 6974 14512
rect 7286 14456 7342 14512
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 5998 10648 6054 10704
rect 6182 10648 6238 10704
rect 5906 9460 5908 9480
rect 5908 9460 5960 9480
rect 5960 9460 5962 9480
rect 5906 9424 5962 9460
rect 5814 7792 5870 7848
rect 6274 10240 6330 10296
rect 6458 10376 6514 10432
rect 6458 10240 6514 10296
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6090 9016 6146 9072
rect 7010 12688 7066 12744
rect 7102 12300 7158 12336
rect 7102 12280 7104 12300
rect 7104 12280 7156 12300
rect 7156 12280 7158 12300
rect 7010 11872 7066 11928
rect 7378 14048 7434 14104
rect 7102 11600 7158 11656
rect 7378 11328 7434 11384
rect 7838 20168 7894 20224
rect 7930 19080 7986 19136
rect 7654 18128 7710 18184
rect 7654 17212 7656 17232
rect 7656 17212 7708 17232
rect 7708 17212 7710 17232
rect 7654 17176 7710 17212
rect 7562 16768 7618 16824
rect 7838 17448 7894 17504
rect 7746 16632 7802 16688
rect 7562 16496 7618 16552
rect 7838 15680 7894 15736
rect 8298 19488 8354 19544
rect 8206 17584 8262 17640
rect 8022 15972 8078 16008
rect 8022 15952 8024 15972
rect 8024 15952 8076 15972
rect 8076 15952 8078 15972
rect 8298 15272 8354 15328
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8758 17484 8760 17504
rect 8760 17484 8812 17504
rect 8812 17484 8814 17504
rect 8758 17448 8814 17484
rect 8666 17196 8722 17232
rect 8666 17176 8668 17196
rect 8668 17176 8720 17196
rect 8720 17176 8722 17196
rect 8574 16904 8630 16960
rect 8574 15816 8630 15872
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 9678 19488 9734 19544
rect 10046 19080 10102 19136
rect 9494 18808 9550 18864
rect 9218 17856 9274 17912
rect 9218 17584 9274 17640
rect 9770 17992 9826 18048
rect 11058 20304 11114 20360
rect 10506 18944 10562 19000
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 9126 15272 9182 15328
rect 8666 15136 8722 15192
rect 8206 14592 8262 14648
rect 8298 13776 8354 13832
rect 8022 12960 8078 13016
rect 8022 12688 8078 12744
rect 7746 12300 7802 12336
rect 7746 12280 7748 12300
rect 7748 12280 7800 12300
rect 7800 12280 7802 12300
rect 7654 11600 7710 11656
rect 7102 10648 7158 10704
rect 7010 10376 7066 10432
rect 6918 10240 6974 10296
rect 6826 9696 6882 9752
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6550 8608 6606 8664
rect 6090 8084 6146 8120
rect 6090 8064 6092 8084
rect 6092 8064 6144 8084
rect 6144 8064 6146 8084
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 7194 10376 7250 10432
rect 7378 10240 7434 10296
rect 7102 8472 7158 8528
rect 8022 11872 8078 11928
rect 7838 10240 7894 10296
rect 7470 8472 7526 8528
rect 5722 6568 5778 6624
rect 5722 5480 5778 5536
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6182 6024 6238 6080
rect 5814 5364 5870 5400
rect 5814 5344 5816 5364
rect 5816 5344 5868 5364
rect 5868 5344 5870 5364
rect 5538 3168 5594 3224
rect 5722 4528 5778 4584
rect 6366 6296 6422 6352
rect 6550 6296 6606 6352
rect 6366 5616 6422 5672
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6090 4664 6146 4720
rect 6458 5108 6460 5128
rect 6460 5108 6512 5128
rect 6512 5108 6514 5128
rect 6458 5072 6514 5108
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6090 3440 6146 3496
rect 6366 4020 6368 4040
rect 6368 4020 6420 4040
rect 6420 4020 6422 4040
rect 6366 3984 6422 4020
rect 6274 3712 6330 3768
rect 6458 3576 6514 3632
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 6826 6296 6882 6352
rect 6918 4528 6974 4584
rect 6918 3576 6974 3632
rect 7378 7656 7434 7712
rect 7378 7112 7434 7168
rect 8298 13096 8354 13152
rect 8206 12552 8262 12608
rect 9126 14728 9182 14784
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 9494 15000 9550 15056
rect 9402 14592 9458 14648
rect 8942 14476 8998 14512
rect 8942 14456 8944 14476
rect 8944 14456 8996 14476
rect 8996 14456 8998 14476
rect 9310 14456 9366 14512
rect 9586 14456 9642 14512
rect 9034 14184 9090 14240
rect 9770 14048 9826 14104
rect 8942 13796 8998 13832
rect 8942 13776 8944 13796
rect 8944 13776 8996 13796
rect 8996 13776 8998 13796
rect 8574 13524 8630 13560
rect 8574 13504 8576 13524
rect 8576 13504 8628 13524
rect 8628 13504 8630 13524
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8574 12416 8630 12472
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8574 11872 8630 11928
rect 8574 11328 8630 11384
rect 9034 11892 9090 11928
rect 9034 11872 9036 11892
rect 9036 11872 9088 11892
rect 9088 11872 9090 11892
rect 9218 12552 9274 12608
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8574 11192 8630 11248
rect 8758 11192 8814 11248
rect 9310 11192 9366 11248
rect 8942 10784 8998 10840
rect 7838 8744 7894 8800
rect 7838 8064 7894 8120
rect 7746 7656 7802 7712
rect 7746 6840 7802 6896
rect 6642 1672 6698 1728
rect 7286 4800 7342 4856
rect 7286 4256 7342 4312
rect 7654 6452 7710 6488
rect 7654 6432 7656 6452
rect 7656 6432 7708 6452
rect 7708 6432 7710 6452
rect 7378 3304 7434 3360
rect 7562 6024 7618 6080
rect 7654 5480 7710 5536
rect 7562 5364 7618 5400
rect 7562 5344 7564 5364
rect 7564 5344 7616 5364
rect 7616 5344 7618 5364
rect 8574 10648 8630 10704
rect 8298 9152 8354 9208
rect 8298 8880 8354 8936
rect 8298 8608 8354 8664
rect 8114 8472 8170 8528
rect 9678 13912 9734 13968
rect 10138 17484 10140 17504
rect 10140 17484 10192 17504
rect 10192 17484 10194 17504
rect 10138 17448 10194 17484
rect 10046 13640 10102 13696
rect 9494 12436 9550 12472
rect 9494 12416 9496 12436
rect 9496 12416 9548 12436
rect 9548 12416 9550 12436
rect 9218 10376 9274 10432
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 9126 10240 9182 10296
rect 9862 12316 9864 12336
rect 9864 12316 9916 12336
rect 9916 12316 9918 12336
rect 9862 12280 9918 12316
rect 9770 10532 9826 10568
rect 9770 10512 9772 10532
rect 9772 10512 9824 10532
rect 9824 10512 9826 10532
rect 9218 9968 9274 10024
rect 9034 9832 9090 9888
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 9126 8744 9182 8800
rect 8574 8200 8630 8256
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8574 8064 8630 8120
rect 8114 6976 8170 7032
rect 8022 6840 8078 6896
rect 7930 6296 7986 6352
rect 8482 6296 8538 6352
rect 7746 3032 7802 3088
rect 7378 2508 7434 2544
rect 7378 2488 7380 2508
rect 7380 2488 7432 2508
rect 7432 2488 7434 2508
rect 7378 1964 7434 2000
rect 7378 1944 7380 1964
rect 7380 1944 7432 1964
rect 7432 1944 7434 1964
rect 3882 40 3938 96
rect 7562 2488 7618 2544
rect 8114 5072 8170 5128
rect 8482 4936 8538 4992
rect 9770 10104 9826 10160
rect 9586 9172 9642 9208
rect 9586 9152 9588 9172
rect 9588 9152 9640 9172
rect 9640 9152 9642 9172
rect 9402 8628 9458 8664
rect 9402 8608 9404 8628
rect 9404 8608 9456 8628
rect 9456 8608 9458 8628
rect 9310 7928 9366 7984
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 9310 6976 9366 7032
rect 9862 9288 9918 9344
rect 9862 8336 9918 8392
rect 10046 11056 10102 11112
rect 10046 10512 10102 10568
rect 10874 17484 10876 17504
rect 10876 17484 10928 17504
rect 10928 17484 10930 17504
rect 10874 17448 10930 17484
rect 10414 15136 10470 15192
rect 10322 14900 10324 14920
rect 10324 14900 10376 14920
rect 10376 14900 10378 14920
rect 10322 14864 10378 14900
rect 10322 13912 10378 13968
rect 10506 13776 10562 13832
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 12990 21392 13046 21448
rect 11610 19796 11612 19816
rect 11612 19796 11664 19816
rect 11664 19796 11666 19816
rect 11610 19760 11666 19796
rect 11794 19660 11796 19680
rect 11796 19660 11848 19680
rect 11848 19660 11850 19680
rect 11794 19624 11850 19660
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11150 17992 11206 18048
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 10966 14764 10968 14784
rect 10968 14764 11020 14784
rect 11020 14764 11022 14784
rect 10966 14728 11022 14764
rect 10322 13232 10378 13288
rect 10230 12280 10286 12336
rect 10230 11056 10286 11112
rect 10782 14320 10838 14376
rect 11058 14320 11114 14376
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 10782 13776 10838 13832
rect 10782 13640 10838 13696
rect 10598 13232 10654 13288
rect 10690 13096 10746 13152
rect 10598 12436 10654 12472
rect 10598 12416 10600 12436
rect 10600 12416 10652 12436
rect 10652 12416 10654 12436
rect 11058 13232 11114 13288
rect 10782 12416 10838 12472
rect 10874 12144 10930 12200
rect 10046 9832 10102 9888
rect 10138 9696 10194 9752
rect 10138 9016 10194 9072
rect 9310 6604 9312 6624
rect 9312 6604 9364 6624
rect 9364 6604 9366 6624
rect 9310 6568 9366 6604
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 9126 5752 9182 5808
rect 8758 5480 8814 5536
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 9310 5888 9366 5944
rect 9770 6432 9826 6488
rect 8114 2896 8170 2952
rect 8206 2644 8262 2680
rect 8206 2624 8208 2644
rect 8208 2624 8260 2644
rect 8260 2624 8262 2644
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 8574 3032 8630 3088
rect 9310 4256 9366 4312
rect 9678 5344 9734 5400
rect 9678 4936 9734 4992
rect 10046 7112 10102 7168
rect 10230 7112 10286 7168
rect 10138 3984 10194 4040
rect 10138 3440 10194 3496
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 10138 3188 10194 3224
rect 10138 3168 10140 3188
rect 10140 3168 10192 3188
rect 10192 3168 10194 3188
rect 10138 2488 10194 2544
rect 10966 11872 11022 11928
rect 12806 19624 12862 19680
rect 12806 19080 12862 19136
rect 12990 17856 13046 17912
rect 12070 16632 12126 16688
rect 12162 16088 12218 16144
rect 12346 16088 12402 16144
rect 11702 15544 11758 15600
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11518 13640 11574 13696
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11886 14184 11942 14240
rect 11794 14068 11850 14104
rect 11794 14048 11796 14068
rect 11796 14048 11848 14068
rect 11848 14048 11850 14068
rect 11794 13812 11796 13832
rect 11796 13812 11848 13832
rect 11848 13812 11850 13832
rect 11794 13776 11850 13812
rect 11794 12824 11850 12880
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 10782 10920 10838 10976
rect 10874 10784 10930 10840
rect 10690 9968 10746 10024
rect 11058 10648 11114 10704
rect 11610 11500 11612 11520
rect 11612 11500 11664 11520
rect 11664 11500 11666 11520
rect 11610 11464 11666 11500
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 10874 8608 10930 8664
rect 11518 9988 11574 10024
rect 11518 9968 11520 9988
rect 11520 9968 11572 9988
rect 11572 9968 11574 9988
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 12254 13812 12256 13832
rect 12256 13812 12308 13832
rect 12308 13812 12310 13832
rect 12254 13776 12310 13812
rect 11978 13368 12034 13424
rect 12254 13404 12256 13424
rect 12256 13404 12308 13424
rect 12308 13404 12310 13424
rect 12254 13368 12310 13404
rect 11978 12824 12034 12880
rect 11978 12436 12034 12472
rect 11978 12416 11980 12436
rect 11980 12416 12032 12436
rect 12032 12416 12034 12436
rect 11978 12144 12034 12200
rect 12162 13132 12164 13152
rect 12164 13132 12216 13152
rect 12216 13132 12218 13152
rect 12162 13096 12218 13132
rect 13082 16224 13138 16280
rect 12530 15000 12586 15056
rect 12438 13640 12494 13696
rect 12530 12824 12586 12880
rect 12254 11736 12310 11792
rect 11794 9288 11850 9344
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11334 8492 11390 8528
rect 11334 8472 11336 8492
rect 11336 8472 11388 8492
rect 11388 8472 11390 8492
rect 10506 7384 10562 7440
rect 10506 4800 10562 4856
rect 10690 5616 10746 5672
rect 11242 7928 11298 7984
rect 11702 7792 11758 7848
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11058 7520 11114 7576
rect 11794 7540 11850 7576
rect 11794 7520 11796 7540
rect 11796 7520 11848 7540
rect 11848 7520 11850 7540
rect 11702 7384 11758 7440
rect 11702 6976 11758 7032
rect 12806 14592 12862 14648
rect 12530 11736 12586 11792
rect 12530 10920 12586 10976
rect 12070 8608 12126 8664
rect 10966 6296 11022 6352
rect 11058 5516 11060 5536
rect 11060 5516 11112 5536
rect 11112 5516 11114 5536
rect 11058 5480 11114 5516
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11518 6024 11574 6080
rect 11334 5908 11390 5944
rect 11334 5888 11336 5908
rect 11336 5888 11388 5908
rect 11388 5888 11390 5908
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11334 5072 11390 5128
rect 10874 3848 10930 3904
rect 11794 4800 11850 4856
rect 11978 5888 12034 5944
rect 11978 5344 12034 5400
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11886 4256 11942 4312
rect 10690 2388 10692 2408
rect 10692 2388 10744 2408
rect 10744 2388 10746 2408
rect 10690 2352 10746 2388
rect 10598 1808 10654 1864
rect 11150 3168 11206 3224
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 11886 3984 11942 4040
rect 13450 18944 13506 19000
rect 13266 18128 13322 18184
rect 12806 11192 12862 11248
rect 12898 9832 12954 9888
rect 12622 9560 12678 9616
rect 12622 7792 12678 7848
rect 13450 17604 13506 17640
rect 13450 17584 13452 17604
rect 13452 17584 13504 17604
rect 13504 17584 13506 17604
rect 13726 19760 13782 19816
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16854 20440 16910 20496
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 14186 15308 14188 15328
rect 14188 15308 14240 15328
rect 14240 15308 14242 15328
rect 14186 15272 14242 15308
rect 14002 15000 14058 15056
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13818 14184 13874 14240
rect 14370 14184 14426 14240
rect 13450 13776 13506 13832
rect 13358 12980 13414 13016
rect 13358 12960 13360 12980
rect 13360 12960 13412 12980
rect 13412 12960 13414 12980
rect 13634 12824 13690 12880
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 14554 13776 14610 13832
rect 14278 13368 14334 13424
rect 13818 12552 13874 12608
rect 13266 11872 13322 11928
rect 13450 12164 13506 12200
rect 13450 12144 13452 12164
rect 13452 12144 13504 12164
rect 13504 12144 13506 12164
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13358 11348 13414 11384
rect 13358 11328 13360 11348
rect 13360 11328 13412 11348
rect 13412 11328 13414 11348
rect 13266 11192 13322 11248
rect 13082 10920 13138 10976
rect 13266 10784 13322 10840
rect 13266 10376 13322 10432
rect 13726 12008 13782 12064
rect 13542 11736 13598 11792
rect 13818 11872 13874 11928
rect 13818 11600 13874 11656
rect 14554 12688 14610 12744
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13634 11076 13690 11112
rect 13634 11056 13636 11076
rect 13636 11056 13688 11076
rect 13688 11056 13690 11076
rect 13174 9424 13230 9480
rect 12990 8744 13046 8800
rect 13082 8356 13138 8392
rect 13082 8336 13084 8356
rect 13084 8336 13136 8356
rect 13136 8336 13138 8356
rect 13082 7928 13138 7984
rect 12898 7520 12954 7576
rect 12530 6976 12586 7032
rect 12438 5616 12494 5672
rect 12438 5072 12494 5128
rect 12346 4936 12402 4992
rect 12622 5616 12678 5672
rect 12898 5616 12954 5672
rect 12162 3440 12218 3496
rect 12070 2896 12126 2952
rect 12438 3168 12494 3224
rect 12990 5072 13046 5128
rect 14462 10784 14518 10840
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13818 9172 13874 9208
rect 13818 9152 13820 9172
rect 13820 9152 13872 9172
rect 13872 9152 13874 9172
rect 14462 10376 14518 10432
rect 13726 8916 13728 8936
rect 13728 8916 13780 8936
rect 13780 8916 13782 8936
rect 13358 7792 13414 7848
rect 13726 8880 13782 8916
rect 13634 8744 13690 8800
rect 13450 6976 13506 7032
rect 13266 6840 13322 6896
rect 13266 6704 13322 6760
rect 13358 5480 13414 5536
rect 12714 3576 12770 3632
rect 13174 3848 13230 3904
rect 13358 4936 13414 4992
rect 13358 4528 13414 4584
rect 13726 6976 13782 7032
rect 14002 8628 14058 8664
rect 14002 8608 14004 8628
rect 14004 8608 14056 8628
rect 14056 8608 14058 8628
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 14278 6160 14334 6216
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 14646 11872 14702 11928
rect 14554 7384 14610 7440
rect 14094 5344 14150 5400
rect 14554 5752 14610 5808
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 14370 4936 14426 4992
rect 14186 3168 14242 3224
rect 13910 2896 13966 2952
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 13726 2624 13782 2680
rect 14462 3848 14518 3904
rect 15290 19236 15346 19272
rect 15290 19216 15292 19236
rect 15292 19216 15344 19236
rect 15344 19216 15346 19236
rect 15474 18672 15530 18728
rect 15658 18264 15714 18320
rect 16118 18808 16174 18864
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 17498 19352 17554 19408
rect 18050 20304 18106 20360
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16302 17876 16358 17912
rect 16302 17856 16304 17876
rect 16304 17856 16356 17876
rect 16356 17856 16358 17876
rect 15750 16496 15806 16552
rect 15014 12144 15070 12200
rect 15014 10240 15070 10296
rect 15290 10104 15346 10160
rect 14738 3712 14794 3768
rect 14738 3440 14794 3496
rect 14370 2932 14372 2952
rect 14372 2932 14424 2952
rect 14424 2932 14426 2952
rect 14370 2896 14426 2932
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16302 16244 16358 16280
rect 16302 16224 16304 16244
rect 16304 16224 16356 16244
rect 16356 16224 16358 16244
rect 16210 14456 16266 14512
rect 16118 13912 16174 13968
rect 15474 9968 15530 10024
rect 15382 8064 15438 8120
rect 15382 7520 15438 7576
rect 15198 7384 15254 7440
rect 15198 6860 15254 6896
rect 15198 6840 15200 6860
rect 15200 6840 15252 6860
rect 15252 6840 15254 6860
rect 15198 5364 15254 5400
rect 15198 5344 15200 5364
rect 15200 5344 15252 5364
rect 15252 5344 15254 5364
rect 15198 5208 15254 5264
rect 15290 4936 15346 4992
rect 15198 4800 15254 4856
rect 15198 4256 15254 4312
rect 15014 992 15070 1048
rect 15566 6024 15622 6080
rect 15566 5888 15622 5944
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 17130 16496 17186 16552
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 17314 14864 17370 14920
rect 17682 17176 17738 17232
rect 16394 14320 16450 14376
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16210 10512 16266 10568
rect 16026 10104 16082 10160
rect 15842 8200 15898 8256
rect 15934 8064 15990 8120
rect 15566 4020 15568 4040
rect 15568 4020 15620 4040
rect 15620 4020 15622 4040
rect 15566 3984 15622 4020
rect 15566 2760 15622 2816
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16762 12588 16764 12608
rect 16764 12588 16816 12608
rect 16816 12588 16818 12608
rect 16762 12552 16818 12588
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16578 11600 16634 11656
rect 17222 12688 17278 12744
rect 17038 11736 17094 11792
rect 16394 11500 16396 11520
rect 16396 11500 16448 11520
rect 16448 11500 16450 11520
rect 16394 11464 16450 11500
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 17038 10648 17094 10704
rect 16854 10376 16910 10432
rect 16118 9696 16174 9752
rect 16210 9560 16266 9616
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16762 9152 16818 9208
rect 16670 9016 16726 9072
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16118 5772 16174 5808
rect 16118 5752 16120 5772
rect 16120 5752 16172 5772
rect 16172 5752 16174 5772
rect 17406 11600 17462 11656
rect 18234 19372 18290 19408
rect 18510 19896 18566 19952
rect 18234 19352 18236 19372
rect 18236 19352 18288 19372
rect 18288 19352 18290 19372
rect 18234 16668 18236 16688
rect 18236 16668 18288 16688
rect 18288 16668 18290 16688
rect 18234 16632 18290 16668
rect 17866 12280 17922 12336
rect 17866 10920 17922 10976
rect 18510 16124 18512 16144
rect 18512 16124 18564 16144
rect 18564 16124 18566 16144
rect 18510 16088 18566 16124
rect 18234 11736 18290 11792
rect 17958 10512 18014 10568
rect 17774 9424 17830 9480
rect 17406 7656 17462 7712
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16302 5752 16358 5808
rect 16578 6160 16634 6216
rect 16946 5888 17002 5944
rect 17406 7112 17462 7168
rect 17314 6568 17370 6624
rect 16302 5480 16358 5536
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16302 5208 16358 5264
rect 16946 5208 17002 5264
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16946 4140 17002 4176
rect 16946 4120 16948 4140
rect 16948 4120 17000 4140
rect 17000 4120 17002 4140
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 17314 5072 17370 5128
rect 17498 6296 17554 6352
rect 17406 3032 17462 3088
rect 18050 9152 18106 9208
rect 17866 9016 17922 9072
rect 17774 7928 17830 7984
rect 17774 7828 17776 7848
rect 17776 7828 17828 7848
rect 17828 7828 17830 7848
rect 17774 7792 17830 7828
rect 17682 6840 17738 6896
rect 17958 8608 18014 8664
rect 17958 7928 18014 7984
rect 17958 7656 18014 7712
rect 17682 6432 17738 6488
rect 18142 6432 18198 6488
rect 17590 4936 17646 4992
rect 17222 2896 17278 2952
rect 17406 2932 17408 2952
rect 17408 2932 17460 2952
rect 17460 2932 17462 2952
rect 17406 2896 17462 2932
rect 16118 2760 16174 2816
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 19062 21800 19118 21856
rect 18970 19352 19026 19408
rect 19522 21392 19578 21448
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19430 19352 19486 19408
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19430 18844 19432 18864
rect 19432 18844 19484 18864
rect 19484 18844 19486 18864
rect 19430 18808 19486 18844
rect 19338 18672 19394 18728
rect 19982 20440 20038 20496
rect 20350 20168 20406 20224
rect 20626 22072 20682 22128
rect 20534 20984 20590 21040
rect 20810 20304 20866 20360
rect 19982 19488 20038 19544
rect 19890 19352 19946 19408
rect 19798 18944 19854 19000
rect 19614 18672 19670 18728
rect 19430 18400 19486 18456
rect 19890 18400 19946 18456
rect 19614 18128 19670 18184
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 20442 19216 20498 19272
rect 20166 18808 20222 18864
rect 20350 18808 20406 18864
rect 20534 18944 20590 19000
rect 20350 18672 20406 18728
rect 20166 18028 20168 18048
rect 20168 18028 20220 18048
rect 20220 18028 20222 18048
rect 20166 17992 20222 18028
rect 20350 18128 20406 18184
rect 21086 19760 21142 19816
rect 20810 17720 20866 17776
rect 20350 16632 20406 16688
rect 19614 16496 19670 16552
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19522 14048 19578 14104
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 18970 12688 19026 12744
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 18694 11192 18750 11248
rect 18326 9152 18382 9208
rect 18326 6160 18382 6216
rect 18326 6060 18328 6080
rect 18328 6060 18380 6080
rect 18380 6060 18382 6080
rect 18326 6024 18382 6060
rect 18326 5888 18382 5944
rect 18510 6568 18566 6624
rect 18510 6296 18566 6352
rect 18694 9968 18750 10024
rect 18786 9832 18842 9888
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 18970 10668 19026 10704
rect 18970 10648 18972 10668
rect 18972 10648 19024 10668
rect 19024 10648 19026 10668
rect 18970 9560 19026 9616
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19430 9424 19486 9480
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19706 13268 19708 13288
rect 19708 13268 19760 13288
rect 19760 13268 19762 13288
rect 19706 13232 19762 13268
rect 20350 16496 20406 16552
rect 18786 8064 18842 8120
rect 18878 6840 18934 6896
rect 18786 6316 18842 6352
rect 18786 6296 18788 6316
rect 18788 6296 18840 6316
rect 18840 6296 18842 6316
rect 18694 6160 18750 6216
rect 18418 5480 18474 5536
rect 18050 3052 18106 3088
rect 18050 3032 18052 3052
rect 18052 3032 18104 3052
rect 18104 3032 18106 3052
rect 18510 4392 18566 4448
rect 19154 8608 19210 8664
rect 19338 8372 19340 8392
rect 19340 8372 19392 8392
rect 19392 8372 19394 8392
rect 19338 8336 19394 8372
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19614 7792 19670 7848
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19246 6568 19302 6624
rect 19154 6432 19210 6488
rect 19614 7112 19670 7168
rect 19890 7928 19946 7984
rect 18878 6024 18934 6080
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 18970 5752 19026 5808
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19430 3984 19486 4040
rect 18970 3848 19026 3904
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 18970 3440 19026 3496
rect 19798 5616 19854 5672
rect 19706 3032 19762 3088
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19706 2896 19762 2952
rect 19890 3732 19946 3768
rect 19890 3712 19892 3732
rect 19892 3712 19944 3732
rect 19944 3712 19946 3732
rect 19798 1808 19854 1864
rect 20350 13812 20352 13832
rect 20352 13812 20404 13832
rect 20404 13812 20406 13832
rect 20350 13776 20406 13812
rect 20810 13912 20866 13968
rect 20626 13504 20682 13560
rect 20810 12280 20866 12336
rect 20718 11600 20774 11656
rect 20718 10920 20774 10976
rect 20166 9560 20222 9616
rect 20626 10004 20628 10024
rect 20628 10004 20680 10024
rect 20680 10004 20682 10024
rect 20626 9968 20682 10004
rect 20258 9288 20314 9344
rect 20534 9832 20590 9888
rect 20718 9016 20774 9072
rect 20350 8336 20406 8392
rect 20258 8200 20314 8256
rect 20442 7828 20444 7848
rect 20444 7828 20496 7848
rect 20496 7828 20498 7848
rect 20442 7792 20498 7828
rect 20166 6976 20222 7032
rect 20442 4664 20498 4720
rect 20258 3984 20314 4040
rect 20350 3848 20406 3904
rect 20626 3712 20682 3768
rect 20074 2624 20130 2680
rect 20534 1264 20590 1320
rect 20534 992 20590 1048
rect 21086 18148 21142 18184
rect 21086 18128 21088 18148
rect 21088 18128 21140 18148
rect 21140 18128 21142 18148
rect 21454 19352 21510 19408
rect 21454 18944 21510 19000
rect 21454 18672 21510 18728
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21454 17720 21510 17776
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21454 17176 21510 17232
rect 21454 16940 21456 16960
rect 21456 16940 21508 16960
rect 21508 16940 21510 16960
rect 21454 16904 21510 16940
rect 21086 16496 21142 16552
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21454 16088 21510 16144
rect 21454 15680 21510 15736
rect 21454 15408 21510 15464
rect 21086 14884 21142 14920
rect 21086 14864 21088 14884
rect 21088 14864 21140 14884
rect 21140 14864 21142 14884
rect 21086 12824 21142 12880
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21454 14456 21510 14512
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21454 13912 21510 13968
rect 21454 13676 21456 13696
rect 21456 13676 21508 13696
rect 21508 13676 21510 13696
rect 21454 13640 21510 13676
rect 21638 13368 21694 13424
rect 21454 13232 21510 13288
rect 21454 12416 21510 12472
rect 21454 12144 21510 12200
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21546 11636 21548 11656
rect 21548 11636 21600 11656
rect 21600 11636 21602 11656
rect 21546 11600 21602 11636
rect 21086 11192 21142 11248
rect 21178 10784 21234 10840
rect 21086 10668 21142 10704
rect 21086 10648 21088 10668
rect 21088 10648 21140 10668
rect 21140 10648 21142 10668
rect 21178 10376 21234 10432
rect 21454 10668 21510 10704
rect 21454 10648 21456 10668
rect 21456 10648 21508 10668
rect 21508 10648 21510 10668
rect 21270 9696 21326 9752
rect 21086 8880 21142 8936
rect 21270 8880 21326 8936
rect 20994 7248 21050 7304
rect 21086 5072 21142 5128
rect 21086 4664 21142 4720
rect 21362 6704 21418 6760
rect 21454 5480 21510 5536
rect 21546 5072 21602 5128
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 22006 9152 22062 9208
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21730 8472 21786 8528
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21914 7384 21970 7440
rect 22006 6704 22062 6760
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 22006 4156 22008 4176
rect 22008 4156 22060 4176
rect 22060 4156 22062 4176
rect 22006 4120 22062 4156
rect 22006 3848 22062 3904
rect 22006 3712 22062 3768
rect 20718 2352 20774 2408
rect 20810 1400 20866 1456
rect 21362 3576 21418 3632
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
rect 21638 584 21694 640
<< metal3 >>
rect 13 22538 79 22541
rect 14590 22538 14596 22540
rect 13 22536 14596 22538
rect 13 22480 18 22536
rect 74 22480 14596 22536
rect 13 22478 14596 22480
rect 13 22475 79 22478
rect 14590 22476 14596 22478
rect 14660 22476 14666 22540
rect 0 22266 800 22296
rect 1577 22266 1643 22269
rect 22200 22266 23000 22296
rect 0 22264 1643 22266
rect 0 22208 1582 22264
rect 1638 22208 1643 22264
rect 0 22206 1643 22208
rect 0 22176 800 22206
rect 1577 22203 1643 22206
rect 20670 22206 23000 22266
rect 20670 22133 20730 22206
rect 22200 22176 23000 22206
rect 20621 22128 20730 22133
rect 20621 22072 20626 22128
rect 20682 22072 20730 22128
rect 20621 22070 20730 22072
rect 20621 22067 20687 22070
rect 0 21858 800 21888
rect 4153 21858 4219 21861
rect 0 21856 4219 21858
rect 0 21800 4158 21856
rect 4214 21800 4219 21856
rect 0 21798 4219 21800
rect 0 21768 800 21798
rect 4153 21795 4219 21798
rect 19057 21858 19123 21861
rect 22200 21858 23000 21888
rect 19057 21856 23000 21858
rect 19057 21800 19062 21856
rect 19118 21800 23000 21856
rect 19057 21798 23000 21800
rect 19057 21795 19123 21798
rect 22200 21768 23000 21798
rect 1158 21660 1164 21724
rect 1228 21722 1234 21724
rect 12934 21722 12940 21724
rect 1228 21662 12940 21722
rect 1228 21660 1234 21662
rect 12934 21660 12940 21662
rect 13004 21660 13010 21724
rect 1710 21524 1716 21588
rect 1780 21586 1786 21588
rect 1780 21526 2790 21586
rect 1780 21524 1786 21526
rect 0 21450 800 21480
rect 1945 21450 2011 21453
rect 0 21448 2011 21450
rect 0 21392 1950 21448
rect 2006 21392 2011 21448
rect 0 21390 2011 21392
rect 2730 21450 2790 21526
rect 12985 21450 13051 21453
rect 2730 21448 13051 21450
rect 2730 21392 12990 21448
rect 13046 21392 13051 21448
rect 2730 21390 13051 21392
rect 0 21360 800 21390
rect 1945 21387 2011 21390
rect 12985 21387 13051 21390
rect 19517 21450 19583 21453
rect 22200 21450 23000 21480
rect 19517 21448 23000 21450
rect 19517 21392 19522 21448
rect 19578 21392 23000 21448
rect 19517 21390 23000 21392
rect 19517 21387 19583 21390
rect 22200 21360 23000 21390
rect 3233 21314 3299 21317
rect 13302 21314 13308 21316
rect 3233 21312 13308 21314
rect 3233 21256 3238 21312
rect 3294 21256 13308 21312
rect 3233 21254 13308 21256
rect 3233 21251 3299 21254
rect 13302 21252 13308 21254
rect 13372 21252 13378 21316
rect 4797 21178 4863 21181
rect 14406 21178 14412 21180
rect 4797 21176 14412 21178
rect 4797 21120 4802 21176
rect 4858 21120 14412 21176
rect 4797 21118 14412 21120
rect 4797 21115 4863 21118
rect 14406 21116 14412 21118
rect 14476 21116 14482 21180
rect 0 21042 800 21072
rect 2221 21042 2287 21045
rect 0 21040 2287 21042
rect 0 20984 2226 21040
rect 2282 20984 2287 21040
rect 0 20982 2287 20984
rect 0 20952 800 20982
rect 2221 20979 2287 20982
rect 3325 21042 3391 21045
rect 7414 21042 7420 21044
rect 3325 21040 7420 21042
rect 3325 20984 3330 21040
rect 3386 20984 7420 21040
rect 3325 20982 7420 20984
rect 3325 20979 3391 20982
rect 7414 20980 7420 20982
rect 7484 20980 7490 21044
rect 20529 21042 20595 21045
rect 22200 21042 23000 21072
rect 20529 21040 23000 21042
rect 20529 20984 20534 21040
rect 20590 20984 23000 21040
rect 20529 20982 23000 20984
rect 20529 20979 20595 20982
rect 22200 20952 23000 20982
rect 4889 20906 4955 20909
rect 7230 20906 7236 20908
rect 4889 20904 7236 20906
rect 4889 20848 4894 20904
rect 4950 20848 7236 20904
rect 4889 20846 7236 20848
rect 4889 20843 4955 20846
rect 7230 20844 7236 20846
rect 7300 20844 7306 20908
rect 6144 20704 6460 20705
rect 0 20634 800 20664
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 1853 20634 1919 20637
rect 22200 20634 23000 20664
rect 0 20632 1919 20634
rect 0 20576 1858 20632
rect 1914 20576 1919 20632
rect 0 20574 1919 20576
rect 0 20544 800 20574
rect 1853 20571 1919 20574
rect 22142 20544 23000 20634
rect 2405 20498 2471 20501
rect 16849 20498 16915 20501
rect 2405 20496 16915 20498
rect 2405 20440 2410 20496
rect 2466 20440 16854 20496
rect 16910 20440 16915 20496
rect 2405 20438 16915 20440
rect 2405 20435 2471 20438
rect 16849 20435 16915 20438
rect 19977 20498 20043 20501
rect 22142 20498 22202 20544
rect 19977 20496 22202 20498
rect 19977 20440 19982 20496
rect 20038 20440 22202 20496
rect 19977 20438 22202 20440
rect 19977 20435 20043 20438
rect 3509 20362 3575 20365
rect 7005 20362 7071 20365
rect 11053 20364 11119 20365
rect 10174 20362 10180 20364
rect 3509 20360 7071 20362
rect 3509 20304 3514 20360
rect 3570 20304 7010 20360
rect 7066 20304 7071 20360
rect 3509 20302 7071 20304
rect 3509 20299 3575 20302
rect 7005 20299 7071 20302
rect 8526 20302 10180 20362
rect 0 20226 800 20256
rect 1485 20226 1551 20229
rect 0 20224 1551 20226
rect 0 20168 1490 20224
rect 1546 20168 1551 20224
rect 0 20166 1551 20168
rect 0 20136 800 20166
rect 1485 20163 1551 20166
rect 3969 20226 4035 20229
rect 5441 20226 5507 20229
rect 7833 20226 7899 20229
rect 3969 20224 5274 20226
rect 3969 20168 3974 20224
rect 4030 20168 5274 20224
rect 3969 20166 5274 20168
rect 3969 20163 4035 20166
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 5214 20090 5274 20166
rect 5441 20224 7899 20226
rect 5441 20168 5446 20224
rect 5502 20168 7838 20224
rect 7894 20168 7899 20224
rect 5441 20166 7899 20168
rect 5441 20163 5507 20166
rect 7833 20163 7899 20166
rect 8526 20090 8586 20302
rect 10174 20300 10180 20302
rect 10244 20300 10250 20364
rect 11053 20362 11100 20364
rect 11008 20360 11100 20362
rect 11008 20304 11058 20360
rect 11008 20302 11100 20304
rect 11053 20300 11100 20302
rect 11164 20300 11170 20364
rect 18045 20362 18111 20365
rect 20805 20362 20871 20365
rect 18045 20360 20871 20362
rect 18045 20304 18050 20360
rect 18106 20304 20810 20360
rect 20866 20304 20871 20360
rect 18045 20302 20871 20304
rect 11053 20299 11119 20300
rect 18045 20299 18111 20302
rect 20805 20299 20871 20302
rect 20345 20226 20411 20229
rect 22200 20226 23000 20256
rect 20345 20224 23000 20226
rect 20345 20168 20350 20224
rect 20406 20168 23000 20224
rect 20345 20166 23000 20168
rect 20345 20163 20411 20166
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 22200 20136 23000 20166
rect 19139 20095 19455 20096
rect 5214 20030 8586 20090
rect 2405 19954 2471 19957
rect 18505 19954 18571 19957
rect 2405 19952 18571 19954
rect 2405 19896 2410 19952
rect 2466 19896 18510 19952
rect 18566 19896 18571 19952
rect 2405 19894 18571 19896
rect 2405 19891 2471 19894
rect 18505 19891 18571 19894
rect 0 19818 800 19848
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19728 800 19758
rect 1853 19755 1919 19758
rect 5349 19818 5415 19821
rect 10542 19818 10548 19820
rect 5349 19816 10548 19818
rect 5349 19760 5354 19816
rect 5410 19760 10548 19816
rect 5349 19758 10548 19760
rect 5349 19755 5415 19758
rect 10542 19756 10548 19758
rect 10612 19756 10618 19820
rect 11605 19818 11671 19821
rect 13721 19818 13787 19821
rect 11605 19816 13787 19818
rect 11605 19760 11610 19816
rect 11666 19760 13726 19816
rect 13782 19760 13787 19816
rect 11605 19758 13787 19760
rect 11605 19755 11671 19758
rect 13721 19755 13787 19758
rect 21081 19818 21147 19821
rect 22200 19818 23000 19848
rect 21081 19816 23000 19818
rect 21081 19760 21086 19816
rect 21142 19760 23000 19816
rect 21081 19758 23000 19760
rect 21081 19755 21147 19758
rect 22200 19728 23000 19758
rect 2957 19682 3023 19685
rect 5942 19682 5948 19684
rect 2957 19680 5948 19682
rect 2957 19624 2962 19680
rect 3018 19624 5948 19680
rect 2957 19622 5948 19624
rect 2957 19619 3023 19622
rect 5942 19620 5948 19622
rect 6012 19620 6018 19684
rect 11789 19682 11855 19685
rect 12801 19682 12867 19685
rect 11789 19680 12867 19682
rect 11789 19624 11794 19680
rect 11850 19624 12806 19680
rect 12862 19624 12867 19680
rect 11789 19622 12867 19624
rect 11789 19619 11855 19622
rect 12801 19619 12867 19622
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 2957 19548 3023 19549
rect 2957 19546 3004 19548
rect 2876 19544 3004 19546
rect 3068 19546 3074 19548
rect 5993 19546 6059 19549
rect 3068 19544 6059 19546
rect 2876 19488 2962 19544
rect 3068 19488 5998 19544
rect 6054 19488 6059 19544
rect 2876 19486 3004 19488
rect 2957 19484 3004 19486
rect 3068 19486 6059 19488
rect 3068 19484 3074 19486
rect 2957 19483 3023 19484
rect 5993 19483 6059 19486
rect 7097 19546 7163 19549
rect 8293 19546 8359 19549
rect 7097 19544 8359 19546
rect 7097 19488 7102 19544
rect 7158 19488 8298 19544
rect 8354 19488 8359 19544
rect 7097 19486 8359 19488
rect 7097 19483 7163 19486
rect 8293 19483 8359 19486
rect 9673 19546 9739 19549
rect 9806 19546 9812 19548
rect 9673 19544 9812 19546
rect 9673 19488 9678 19544
rect 9734 19488 9812 19544
rect 9673 19486 9812 19488
rect 9673 19483 9739 19486
rect 9806 19484 9812 19486
rect 9876 19484 9882 19548
rect 19977 19546 20043 19549
rect 19977 19544 20362 19546
rect 19977 19488 19982 19544
rect 20038 19488 20362 19544
rect 19977 19486 20362 19488
rect 19977 19483 20043 19486
rect 0 19410 800 19440
rect 1485 19410 1551 19413
rect 0 19408 1551 19410
rect 0 19352 1490 19408
rect 1546 19352 1551 19408
rect 0 19350 1551 19352
rect 0 19320 800 19350
rect 1485 19347 1551 19350
rect 1945 19410 2011 19413
rect 17493 19410 17559 19413
rect 1945 19408 17559 19410
rect 1945 19352 1950 19408
rect 2006 19352 17498 19408
rect 17554 19352 17559 19408
rect 1945 19350 17559 19352
rect 1945 19347 2011 19350
rect 17493 19347 17559 19350
rect 18229 19410 18295 19413
rect 18965 19410 19031 19413
rect 19425 19410 19491 19413
rect 18229 19408 19491 19410
rect 18229 19352 18234 19408
rect 18290 19352 18970 19408
rect 19026 19352 19430 19408
rect 19486 19352 19491 19408
rect 18229 19350 19491 19352
rect 18229 19347 18295 19350
rect 18965 19347 19031 19350
rect 19425 19347 19491 19350
rect 19558 19348 19564 19412
rect 19628 19410 19634 19412
rect 19885 19410 19951 19413
rect 19628 19408 19951 19410
rect 19628 19352 19890 19408
rect 19946 19352 19951 19408
rect 19628 19350 19951 19352
rect 19628 19348 19634 19350
rect 19885 19347 19951 19350
rect 3233 19274 3299 19277
rect 3366 19274 3372 19276
rect 3233 19272 3372 19274
rect 3233 19216 3238 19272
rect 3294 19216 3372 19272
rect 3233 19214 3372 19216
rect 3233 19211 3299 19214
rect 3366 19212 3372 19214
rect 3436 19212 3442 19276
rect 3601 19274 3667 19277
rect 5901 19274 5967 19277
rect 3601 19272 5967 19274
rect 3601 19216 3606 19272
rect 3662 19216 5906 19272
rect 5962 19216 5967 19272
rect 3601 19214 5967 19216
rect 3601 19211 3667 19214
rect 5901 19211 5967 19214
rect 7005 19274 7071 19277
rect 15285 19274 15351 19277
rect 7005 19272 15351 19274
rect 7005 19216 7010 19272
rect 7066 19216 15290 19272
rect 15346 19216 15351 19272
rect 7005 19214 15351 19216
rect 20302 19274 20362 19486
rect 21449 19410 21515 19413
rect 22200 19410 23000 19440
rect 21449 19408 23000 19410
rect 21449 19352 21454 19408
rect 21510 19352 23000 19408
rect 21449 19350 23000 19352
rect 21449 19347 21515 19350
rect 22200 19320 23000 19350
rect 20437 19274 20503 19277
rect 20302 19272 20503 19274
rect 20302 19216 20442 19272
rect 20498 19216 20503 19272
rect 20302 19214 20503 19216
rect 7005 19211 7071 19214
rect 15285 19211 15351 19214
rect 20437 19211 20503 19214
rect 5073 19138 5139 19141
rect 7373 19138 7439 19141
rect 7925 19138 7991 19141
rect 5073 19136 7991 19138
rect 5073 19080 5078 19136
rect 5134 19080 7378 19136
rect 7434 19080 7930 19136
rect 7986 19080 7991 19136
rect 5073 19078 7991 19080
rect 5073 19075 5139 19078
rect 7373 19075 7439 19078
rect 7925 19075 7991 19078
rect 10041 19138 10107 19141
rect 12801 19138 12867 19141
rect 10041 19136 12867 19138
rect 10041 19080 10046 19136
rect 10102 19080 12806 19136
rect 12862 19080 12867 19136
rect 10041 19078 12867 19080
rect 10041 19075 10107 19078
rect 12801 19075 12867 19078
rect 3545 19072 3861 19073
rect 0 19002 800 19032
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 1485 19002 1551 19005
rect 0 19000 1551 19002
rect 0 18944 1490 19000
rect 1546 18944 1551 19000
rect 0 18942 1551 18944
rect 0 18912 800 18942
rect 1485 18939 1551 18942
rect 10501 19002 10567 19005
rect 13445 19002 13511 19005
rect 10501 19000 13511 19002
rect 10501 18944 10506 19000
rect 10562 18944 13450 19000
rect 13506 18944 13511 19000
rect 10501 18942 13511 18944
rect 10501 18939 10567 18942
rect 13445 18939 13511 18942
rect 19793 19002 19859 19005
rect 20529 19002 20595 19005
rect 19793 19000 20595 19002
rect 19793 18944 19798 19000
rect 19854 18944 20534 19000
rect 20590 18944 20595 19000
rect 19793 18942 20595 18944
rect 19793 18939 19859 18942
rect 20529 18939 20595 18942
rect 21449 19002 21515 19005
rect 22200 19002 23000 19032
rect 21449 19000 23000 19002
rect 21449 18944 21454 19000
rect 21510 18944 23000 19000
rect 21449 18942 23000 18944
rect 21449 18939 21515 18942
rect 22200 18912 23000 18942
rect 2589 18866 2655 18869
rect 3877 18868 3943 18869
rect 3877 18866 3924 18868
rect 2589 18864 2698 18866
rect 2589 18808 2594 18864
rect 2650 18808 2698 18864
rect 2589 18803 2698 18808
rect 3832 18864 3924 18866
rect 3832 18808 3882 18864
rect 3832 18806 3924 18808
rect 3877 18804 3924 18806
rect 3988 18804 3994 18868
rect 9489 18866 9555 18869
rect 16113 18866 16179 18869
rect 9489 18864 16179 18866
rect 9489 18808 9494 18864
rect 9550 18808 16118 18864
rect 16174 18808 16179 18864
rect 9489 18806 16179 18808
rect 3877 18803 3943 18804
rect 9489 18803 9555 18806
rect 16113 18803 16179 18806
rect 19425 18866 19491 18869
rect 20161 18866 20227 18869
rect 19425 18864 20227 18866
rect 19425 18808 19430 18864
rect 19486 18808 20166 18864
rect 20222 18808 20227 18864
rect 19425 18806 20227 18808
rect 19425 18803 19491 18806
rect 20161 18803 20227 18806
rect 20345 18866 20411 18869
rect 20345 18864 20546 18866
rect 20345 18808 20350 18864
rect 20406 18808 20546 18864
rect 20345 18806 20546 18808
rect 20345 18803 20411 18806
rect 2638 18730 2698 18803
rect 4061 18730 4127 18733
rect 15469 18730 15535 18733
rect 2638 18670 2790 18730
rect 0 18594 800 18624
rect 1945 18594 2011 18597
rect 0 18592 2011 18594
rect 0 18536 1950 18592
rect 2006 18536 2011 18592
rect 0 18534 2011 18536
rect 0 18504 800 18534
rect 1945 18531 2011 18534
rect 2730 18458 2790 18670
rect 4061 18728 15535 18730
rect 4061 18672 4066 18728
rect 4122 18672 15474 18728
rect 15530 18672 15535 18728
rect 4061 18670 15535 18672
rect 4061 18667 4127 18670
rect 15469 18667 15535 18670
rect 19333 18730 19399 18733
rect 19609 18730 19675 18733
rect 20345 18730 20411 18733
rect 19333 18728 19442 18730
rect 19333 18672 19338 18728
rect 19394 18672 19442 18728
rect 19333 18667 19442 18672
rect 19609 18728 20411 18730
rect 19609 18672 19614 18728
rect 19670 18672 20350 18728
rect 20406 18672 20411 18728
rect 19609 18670 20411 18672
rect 19609 18667 19675 18670
rect 20345 18667 20411 18670
rect 19382 18594 19442 18667
rect 20486 18594 20546 18806
rect 21449 18730 21515 18733
rect 21449 18728 22202 18730
rect 21449 18672 21454 18728
rect 21510 18672 22202 18728
rect 21449 18670 22202 18672
rect 21449 18667 21515 18670
rect 19382 18534 20546 18594
rect 22142 18624 22202 18670
rect 22142 18534 23000 18624
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 22200 18504 23000 18534
rect 21738 18463 22054 18464
rect 4521 18458 4587 18461
rect 19425 18458 19491 18461
rect 19885 18458 19951 18461
rect 2730 18456 6010 18458
rect 2730 18400 4526 18456
rect 4582 18400 6010 18456
rect 2730 18398 6010 18400
rect 4521 18395 4587 18398
rect 3417 18322 3483 18325
rect 5022 18322 5028 18324
rect 3417 18320 5028 18322
rect 3417 18264 3422 18320
rect 3478 18264 5028 18320
rect 3417 18262 5028 18264
rect 3417 18259 3483 18262
rect 5022 18260 5028 18262
rect 5092 18260 5098 18324
rect 5950 18322 6010 18398
rect 19425 18456 19951 18458
rect 19425 18400 19430 18456
rect 19486 18400 19890 18456
rect 19946 18400 19951 18456
rect 19425 18398 19951 18400
rect 19425 18395 19491 18398
rect 19885 18395 19951 18398
rect 15653 18322 15719 18325
rect 5950 18320 15719 18322
rect 5950 18264 15658 18320
rect 15714 18264 15719 18320
rect 5950 18262 15719 18264
rect 15653 18259 15719 18262
rect 0 18186 800 18216
rect 1485 18186 1551 18189
rect 0 18184 1551 18186
rect 0 18128 1490 18184
rect 1546 18128 1551 18184
rect 0 18126 1551 18128
rect 0 18096 800 18126
rect 1485 18123 1551 18126
rect 7649 18186 7715 18189
rect 13261 18186 13327 18189
rect 7649 18184 13327 18186
rect 7649 18128 7654 18184
rect 7710 18128 13266 18184
rect 13322 18128 13327 18184
rect 7649 18126 13327 18128
rect 7649 18123 7715 18126
rect 13261 18123 13327 18126
rect 19609 18186 19675 18189
rect 20345 18186 20411 18189
rect 19609 18184 20411 18186
rect 19609 18128 19614 18184
rect 19670 18128 20350 18184
rect 20406 18128 20411 18184
rect 19609 18126 20411 18128
rect 19609 18123 19675 18126
rect 20345 18123 20411 18126
rect 21081 18186 21147 18189
rect 22200 18186 23000 18216
rect 21081 18184 23000 18186
rect 21081 18128 21086 18184
rect 21142 18128 23000 18184
rect 21081 18126 23000 18128
rect 21081 18123 21147 18126
rect 22200 18096 23000 18126
rect 9254 17988 9260 18052
rect 9324 18050 9330 18052
rect 9765 18050 9831 18053
rect 9324 18048 9831 18050
rect 9324 17992 9770 18048
rect 9826 17992 9831 18048
rect 9324 17990 9831 17992
rect 9324 17988 9330 17990
rect 9765 17987 9831 17990
rect 11145 18050 11211 18053
rect 12014 18050 12020 18052
rect 11145 18048 12020 18050
rect 11145 17992 11150 18048
rect 11206 17992 12020 18048
rect 11145 17990 12020 17992
rect 11145 17987 11211 17990
rect 12014 17988 12020 17990
rect 12084 17988 12090 18052
rect 20161 18050 20227 18053
rect 20478 18050 20484 18052
rect 20161 18048 20484 18050
rect 20161 17992 20166 18048
rect 20222 17992 20484 18048
rect 20161 17990 20484 17992
rect 20161 17987 20227 17990
rect 20478 17988 20484 17990
rect 20548 17988 20554 18052
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 4521 17914 4587 17917
rect 5206 17914 5212 17916
rect 4521 17912 5212 17914
rect 4521 17856 4526 17912
rect 4582 17856 5212 17912
rect 4521 17854 5212 17856
rect 4521 17851 4587 17854
rect 5206 17852 5212 17854
rect 5276 17852 5282 17916
rect 9213 17914 9279 17917
rect 12985 17914 13051 17917
rect 9213 17912 13051 17914
rect 9213 17856 9218 17912
rect 9274 17856 12990 17912
rect 13046 17856 13051 17912
rect 9213 17854 13051 17856
rect 9213 17851 9279 17854
rect 12985 17851 13051 17854
rect 16297 17914 16363 17917
rect 17166 17914 17172 17916
rect 16297 17912 17172 17914
rect 16297 17856 16302 17912
rect 16358 17856 17172 17912
rect 16297 17854 17172 17856
rect 16297 17851 16363 17854
rect 17166 17852 17172 17854
rect 17236 17852 17242 17916
rect 0 17778 800 17808
rect 1485 17778 1551 17781
rect 0 17776 1551 17778
rect 0 17720 1490 17776
rect 1546 17720 1551 17776
rect 0 17718 1551 17720
rect 0 17688 800 17718
rect 1485 17715 1551 17718
rect 4245 17778 4311 17781
rect 4705 17778 4771 17781
rect 4245 17776 4771 17778
rect 4245 17720 4250 17776
rect 4306 17720 4710 17776
rect 4766 17720 4771 17776
rect 4245 17718 4771 17720
rect 4245 17715 4311 17718
rect 4705 17715 4771 17718
rect 5349 17778 5415 17781
rect 6453 17778 6519 17781
rect 20805 17778 20871 17781
rect 5349 17776 20871 17778
rect 5349 17720 5354 17776
rect 5410 17720 6458 17776
rect 6514 17720 20810 17776
rect 20866 17720 20871 17776
rect 5349 17718 20871 17720
rect 5349 17715 5415 17718
rect 6453 17715 6519 17718
rect 20805 17715 20871 17718
rect 21449 17778 21515 17781
rect 22200 17778 23000 17808
rect 21449 17776 23000 17778
rect 21449 17720 21454 17776
rect 21510 17720 23000 17776
rect 21449 17718 23000 17720
rect 21449 17715 21515 17718
rect 22200 17688 23000 17718
rect 2589 17642 2655 17645
rect 3601 17642 3667 17645
rect 2589 17640 3667 17642
rect 2589 17584 2594 17640
rect 2650 17584 3606 17640
rect 3662 17584 3667 17640
rect 2589 17582 3667 17584
rect 2589 17579 2655 17582
rect 3601 17579 3667 17582
rect 4521 17642 4587 17645
rect 5073 17642 5139 17645
rect 8201 17642 8267 17645
rect 9213 17642 9279 17645
rect 13445 17642 13511 17645
rect 4521 17640 9279 17642
rect 4521 17584 4526 17640
rect 4582 17584 5078 17640
rect 5134 17584 8206 17640
rect 8262 17584 9218 17640
rect 9274 17584 9279 17640
rect 4521 17582 9279 17584
rect 4521 17579 4587 17582
rect 5073 17579 5139 17582
rect 8201 17579 8267 17582
rect 9213 17579 9279 17582
rect 9446 17640 13511 17642
rect 9446 17584 13450 17640
rect 13506 17584 13511 17640
rect 9446 17582 13511 17584
rect 7833 17506 7899 17509
rect 8753 17506 8819 17509
rect 7833 17504 8819 17506
rect 7833 17448 7838 17504
rect 7894 17448 8758 17504
rect 8814 17448 8819 17504
rect 7833 17446 8819 17448
rect 7833 17443 7899 17446
rect 8753 17443 8819 17446
rect 6144 17440 6460 17441
rect 0 17370 800 17400
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 1485 17370 1551 17373
rect 0 17368 1551 17370
rect 0 17312 1490 17368
rect 1546 17312 1551 17368
rect 0 17310 1551 17312
rect 0 17280 800 17310
rect 1485 17307 1551 17310
rect 2589 17370 2655 17373
rect 5717 17370 5783 17373
rect 9446 17370 9506 17582
rect 13445 17579 13511 17582
rect 10133 17506 10199 17509
rect 10869 17506 10935 17509
rect 10133 17504 10935 17506
rect 10133 17448 10138 17504
rect 10194 17448 10874 17504
rect 10930 17448 10935 17504
rect 10133 17446 10935 17448
rect 10133 17443 10199 17446
rect 10869 17443 10935 17446
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 22200 17370 23000 17400
rect 2589 17368 5783 17370
rect 2589 17312 2594 17368
rect 2650 17312 5722 17368
rect 5778 17312 5783 17368
rect 2589 17310 5783 17312
rect 2589 17307 2655 17310
rect 5717 17307 5783 17310
rect 6686 17310 9506 17370
rect 5165 17234 5231 17237
rect 6686 17234 6746 17310
rect 22142 17280 23000 17370
rect 7649 17236 7715 17237
rect 5165 17232 6746 17234
rect 5165 17176 5170 17232
rect 5226 17176 6746 17232
rect 5165 17174 6746 17176
rect 5165 17171 5231 17174
rect 7598 17172 7604 17236
rect 7668 17234 7715 17236
rect 8661 17234 8727 17237
rect 17677 17234 17743 17237
rect 7668 17232 7760 17234
rect 7710 17176 7760 17232
rect 7668 17174 7760 17176
rect 8661 17232 17743 17234
rect 8661 17176 8666 17232
rect 8722 17176 17682 17232
rect 17738 17176 17743 17232
rect 8661 17174 17743 17176
rect 7668 17172 7715 17174
rect 7606 17171 7715 17172
rect 8661 17171 8727 17174
rect 17677 17171 17743 17174
rect 21449 17234 21515 17237
rect 22142 17234 22202 17280
rect 21449 17232 22202 17234
rect 21449 17176 21454 17232
rect 21510 17176 22202 17232
rect 21449 17174 22202 17176
rect 21449 17171 21515 17174
rect 2221 17098 2287 17101
rect 7606 17098 7666 17171
rect 2221 17096 7666 17098
rect 2221 17040 2226 17096
rect 2282 17040 7666 17096
rect 2221 17038 7666 17040
rect 2221 17035 2287 17038
rect 0 16962 800 16992
rect 1485 16962 1551 16965
rect 0 16960 1551 16962
rect 0 16904 1490 16960
rect 1546 16904 1551 16960
rect 0 16902 1551 16904
rect 0 16872 800 16902
rect 1485 16899 1551 16902
rect 5717 16962 5783 16965
rect 6678 16962 6684 16964
rect 5717 16960 6684 16962
rect 5717 16904 5722 16960
rect 5778 16904 6684 16960
rect 5717 16902 6684 16904
rect 5717 16899 5783 16902
rect 6678 16900 6684 16902
rect 6748 16962 6754 16964
rect 8569 16962 8635 16965
rect 6748 16960 8635 16962
rect 6748 16904 8574 16960
rect 8630 16904 8635 16960
rect 6748 16902 8635 16904
rect 6748 16900 6754 16902
rect 8569 16899 8635 16902
rect 21449 16962 21515 16965
rect 22200 16962 23000 16992
rect 21449 16960 23000 16962
rect 21449 16904 21454 16960
rect 21510 16904 23000 16960
rect 21449 16902 23000 16904
rect 21449 16899 21515 16902
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 22200 16872 23000 16902
rect 19139 16831 19455 16832
rect 7557 16826 7623 16829
rect 7557 16824 8586 16826
rect 7557 16768 7562 16824
rect 7618 16768 8586 16824
rect 7557 16766 8586 16768
rect 7557 16763 7666 16766
rect 1894 16628 1900 16692
rect 1964 16690 1970 16692
rect 5349 16690 5415 16693
rect 1964 16688 5415 16690
rect 1964 16632 5354 16688
rect 5410 16632 5415 16688
rect 1964 16630 5415 16632
rect 7606 16690 7666 16763
rect 7741 16690 7807 16693
rect 7606 16688 7807 16690
rect 7606 16632 7746 16688
rect 7802 16632 7807 16688
rect 7606 16630 7807 16632
rect 8526 16690 8586 16766
rect 12065 16690 12131 16693
rect 8526 16688 12131 16690
rect 8526 16632 12070 16688
rect 12126 16632 12131 16688
rect 8526 16630 12131 16632
rect 1964 16628 1970 16630
rect 5349 16627 5415 16630
rect 7741 16627 7807 16630
rect 12065 16627 12131 16630
rect 18229 16690 18295 16693
rect 20345 16692 20411 16693
rect 19742 16690 19748 16692
rect 18229 16688 19748 16690
rect 18229 16632 18234 16688
rect 18290 16632 19748 16688
rect 18229 16630 19748 16632
rect 18229 16627 18295 16630
rect 19742 16628 19748 16630
rect 19812 16628 19818 16692
rect 20294 16690 20300 16692
rect 20254 16630 20300 16690
rect 20364 16688 20411 16692
rect 20406 16632 20411 16688
rect 20294 16628 20300 16630
rect 20364 16628 20411 16632
rect 20345 16627 20411 16628
rect 0 16554 800 16584
rect 1853 16554 1919 16557
rect 7557 16554 7623 16557
rect 15745 16556 15811 16557
rect 15694 16554 15700 16556
rect 0 16552 1919 16554
rect 0 16496 1858 16552
rect 1914 16496 1919 16552
rect 0 16494 1919 16496
rect 0 16464 800 16494
rect 1853 16491 1919 16494
rect 2086 16494 7436 16554
rect 974 16356 980 16420
rect 1044 16418 1050 16420
rect 2086 16418 2146 16494
rect 1044 16358 2146 16418
rect 2497 16418 2563 16421
rect 5073 16418 5139 16421
rect 2497 16416 5139 16418
rect 2497 16360 2502 16416
rect 2558 16360 5078 16416
rect 5134 16360 5139 16416
rect 2497 16358 5139 16360
rect 1044 16356 1050 16358
rect 2497 16355 2563 16358
rect 5073 16355 5139 16358
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 1117 16282 1183 16285
rect 5993 16282 6059 16285
rect 1117 16280 6059 16282
rect 1117 16224 1122 16280
rect 1178 16224 5998 16280
rect 6054 16224 6059 16280
rect 1117 16222 6059 16224
rect 1117 16219 1183 16222
rect 5993 16219 6059 16222
rect 0 16146 800 16176
rect 1485 16146 1551 16149
rect 0 16144 1551 16146
rect 0 16088 1490 16144
rect 1546 16088 1551 16144
rect 0 16086 1551 16088
rect 7376 16146 7436 16494
rect 7557 16552 15700 16554
rect 15764 16554 15811 16556
rect 17125 16554 17191 16557
rect 19609 16554 19675 16557
rect 20345 16554 20411 16557
rect 15764 16552 15892 16554
rect 7557 16496 7562 16552
rect 7618 16496 15700 16552
rect 15806 16496 15892 16552
rect 7557 16494 15700 16496
rect 7557 16491 7623 16494
rect 15694 16492 15700 16494
rect 15764 16494 15892 16496
rect 17125 16552 20411 16554
rect 17125 16496 17130 16552
rect 17186 16496 19614 16552
rect 19670 16496 20350 16552
rect 20406 16496 20411 16552
rect 17125 16494 20411 16496
rect 15764 16492 15811 16494
rect 15745 16491 15811 16492
rect 17125 16491 17191 16494
rect 19609 16491 19675 16494
rect 20345 16491 20411 16494
rect 21081 16554 21147 16557
rect 22200 16554 23000 16584
rect 21081 16552 23000 16554
rect 21081 16496 21086 16552
rect 21142 16496 23000 16552
rect 21081 16494 23000 16496
rect 21081 16491 21147 16494
rect 22200 16464 23000 16494
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 13077 16282 13143 16285
rect 16297 16282 16363 16285
rect 13077 16280 16363 16282
rect 13077 16224 13082 16280
rect 13138 16224 16302 16280
rect 16358 16224 16363 16280
rect 13077 16222 16363 16224
rect 13077 16219 13143 16222
rect 16297 16219 16363 16222
rect 12157 16146 12223 16149
rect 7376 16144 12223 16146
rect 7376 16088 12162 16144
rect 12218 16088 12223 16144
rect 7376 16086 12223 16088
rect 0 16056 800 16086
rect 1485 16083 1551 16086
rect 12157 16083 12223 16086
rect 12341 16146 12407 16149
rect 18505 16146 18571 16149
rect 12341 16144 18571 16146
rect 12341 16088 12346 16144
rect 12402 16088 18510 16144
rect 18566 16088 18571 16144
rect 12341 16086 18571 16088
rect 12341 16083 12407 16086
rect 18505 16083 18571 16086
rect 21449 16146 21515 16149
rect 22200 16146 23000 16176
rect 21449 16144 23000 16146
rect 21449 16088 21454 16144
rect 21510 16088 23000 16144
rect 21449 16086 23000 16088
rect 21449 16083 21515 16086
rect 22200 16056 23000 16086
rect 2589 16010 2655 16013
rect 5993 16010 6059 16013
rect 2589 16008 6059 16010
rect 2589 15952 2594 16008
rect 2650 15952 5998 16008
rect 6054 15952 6059 16008
rect 2589 15950 6059 15952
rect 2589 15947 2655 15950
rect 5993 15947 6059 15950
rect 8017 16010 8083 16013
rect 17534 16010 17540 16012
rect 8017 16008 17540 16010
rect 8017 15952 8022 16008
rect 8078 15952 17540 16008
rect 8017 15950 17540 15952
rect 8017 15947 8083 15950
rect 17534 15948 17540 15950
rect 17604 15948 17610 16012
rect 4521 15874 4587 15877
rect 8569 15874 8635 15877
rect 4521 15872 8635 15874
rect 4521 15816 4526 15872
rect 4582 15816 8574 15872
rect 8630 15816 8635 15872
rect 4521 15814 8635 15816
rect 4521 15811 4587 15814
rect 8569 15811 8635 15814
rect 3545 15808 3861 15809
rect 0 15738 800 15768
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 1485 15738 1551 15741
rect 0 15736 1551 15738
rect 0 15680 1490 15736
rect 1546 15680 1551 15736
rect 0 15678 1551 15680
rect 0 15648 800 15678
rect 1485 15675 1551 15678
rect 4838 15676 4844 15740
rect 4908 15738 4914 15740
rect 7833 15738 7899 15741
rect 4908 15736 7899 15738
rect 4908 15680 7838 15736
rect 7894 15680 7899 15736
rect 4908 15678 7899 15680
rect 4908 15676 4914 15678
rect 7833 15675 7899 15678
rect 21449 15738 21515 15741
rect 22200 15738 23000 15768
rect 21449 15736 23000 15738
rect 21449 15680 21454 15736
rect 21510 15680 23000 15736
rect 21449 15678 23000 15680
rect 21449 15675 21515 15678
rect 22200 15648 23000 15678
rect 2313 15602 2379 15605
rect 5901 15602 5967 15605
rect 2313 15600 5967 15602
rect 2313 15544 2318 15600
rect 2374 15544 5906 15600
rect 5962 15544 5967 15600
rect 2313 15542 5967 15544
rect 2313 15539 2379 15542
rect 5901 15539 5967 15542
rect 6637 15602 6703 15605
rect 11697 15602 11763 15605
rect 6637 15600 11763 15602
rect 6637 15544 6642 15600
rect 6698 15544 11702 15600
rect 11758 15544 11763 15600
rect 6637 15542 11763 15544
rect 6637 15539 6703 15542
rect 11697 15539 11763 15542
rect 3918 15404 3924 15468
rect 3988 15466 3994 15468
rect 4061 15466 4127 15469
rect 3988 15464 4127 15466
rect 3988 15408 4066 15464
rect 4122 15408 4127 15464
rect 3988 15406 4127 15408
rect 3988 15404 3994 15406
rect 4061 15403 4127 15406
rect 5349 15466 5415 15469
rect 19558 15466 19564 15468
rect 5349 15464 19564 15466
rect 5349 15408 5354 15464
rect 5410 15408 19564 15464
rect 5349 15406 19564 15408
rect 5349 15403 5415 15406
rect 19558 15404 19564 15406
rect 19628 15404 19634 15468
rect 21449 15466 21515 15469
rect 21449 15464 22202 15466
rect 21449 15408 21454 15464
rect 21510 15408 22202 15464
rect 21449 15406 22202 15408
rect 21449 15403 21515 15406
rect 22142 15360 22202 15406
rect 0 15330 800 15360
rect 1485 15330 1551 15333
rect 3049 15332 3115 15333
rect 0 15328 1551 15330
rect 0 15272 1490 15328
rect 1546 15272 1551 15328
rect 0 15270 1551 15272
rect 0 15240 800 15270
rect 1485 15267 1551 15270
rect 2998 15268 3004 15332
rect 3068 15330 3115 15332
rect 4153 15330 4219 15333
rect 8293 15332 8359 15333
rect 4286 15330 4292 15332
rect 3068 15328 3160 15330
rect 3110 15272 3160 15328
rect 3068 15270 3160 15272
rect 4153 15328 4292 15330
rect 4153 15272 4158 15328
rect 4214 15272 4292 15328
rect 4153 15270 4292 15272
rect 3068 15268 3115 15270
rect 3049 15267 3115 15268
rect 4153 15267 4219 15270
rect 4286 15268 4292 15270
rect 4356 15268 4362 15332
rect 8293 15328 8340 15332
rect 8404 15330 8410 15332
rect 9121 15330 9187 15333
rect 8293 15272 8298 15328
rect 8293 15268 8340 15272
rect 8404 15270 8450 15330
rect 8526 15328 9187 15330
rect 8526 15272 9126 15328
rect 9182 15272 9187 15328
rect 8526 15270 9187 15272
rect 8404 15268 8410 15270
rect 8293 15267 8359 15268
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 2589 15194 2655 15197
rect 4521 15194 4587 15197
rect 5901 15196 5967 15197
rect 5901 15194 5948 15196
rect 2589 15192 4587 15194
rect 2589 15136 2594 15192
rect 2650 15136 4526 15192
rect 4582 15136 4587 15192
rect 2589 15134 4587 15136
rect 5856 15192 5948 15194
rect 5856 15136 5906 15192
rect 5856 15134 5948 15136
rect 2589 15131 2655 15134
rect 4521 15131 4587 15134
rect 5901 15132 5948 15134
rect 6012 15132 6018 15196
rect 7046 15132 7052 15196
rect 7116 15194 7122 15196
rect 8526 15194 8586 15270
rect 9121 15267 9187 15270
rect 11830 15268 11836 15332
rect 11900 15330 11906 15332
rect 14181 15330 14247 15333
rect 11900 15328 14247 15330
rect 11900 15272 14186 15328
rect 14242 15272 14247 15328
rect 11900 15270 14247 15272
rect 22142 15270 23000 15360
rect 11900 15268 11906 15270
rect 14181 15267 14247 15270
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 22200 15240 23000 15270
rect 21738 15199 22054 15200
rect 7116 15134 8586 15194
rect 8661 15194 8727 15197
rect 10409 15194 10475 15197
rect 8661 15192 10475 15194
rect 8661 15136 8666 15192
rect 8722 15136 10414 15192
rect 10470 15136 10475 15192
rect 8661 15134 10475 15136
rect 7116 15132 7122 15134
rect 5901 15131 5967 15132
rect 8661 15131 8727 15134
rect 10409 15131 10475 15134
rect 3233 15058 3299 15061
rect 5717 15058 5783 15061
rect 9489 15058 9555 15061
rect 3233 15056 9555 15058
rect 3233 15000 3238 15056
rect 3294 15000 5722 15056
rect 5778 15000 9494 15056
rect 9550 15000 9555 15056
rect 3233 14998 9555 15000
rect 3233 14995 3299 14998
rect 5717 14995 5783 14998
rect 9489 14995 9555 14998
rect 12525 15058 12591 15061
rect 13997 15058 14063 15061
rect 12525 15056 14063 15058
rect 12525 15000 12530 15056
rect 12586 15000 14002 15056
rect 14058 15000 14063 15056
rect 12525 14998 14063 15000
rect 12525 14995 12591 14998
rect 13997 14995 14063 14998
rect 0 14922 800 14952
rect 1853 14922 1919 14925
rect 0 14920 1919 14922
rect 0 14864 1858 14920
rect 1914 14864 1919 14920
rect 0 14862 1919 14864
rect 0 14832 800 14862
rect 1853 14859 1919 14862
rect 10317 14922 10383 14925
rect 17309 14922 17375 14925
rect 10317 14920 17375 14922
rect 10317 14864 10322 14920
rect 10378 14864 17314 14920
rect 17370 14864 17375 14920
rect 10317 14862 17375 14864
rect 10317 14859 10383 14862
rect 17309 14859 17375 14862
rect 21081 14922 21147 14925
rect 22200 14922 23000 14952
rect 21081 14920 23000 14922
rect 21081 14864 21086 14920
rect 21142 14864 23000 14920
rect 21081 14862 23000 14864
rect 21081 14859 21147 14862
rect 22200 14832 23000 14862
rect 9121 14786 9187 14789
rect 10961 14786 11027 14789
rect 9121 14784 11027 14786
rect 9121 14728 9126 14784
rect 9182 14728 10966 14784
rect 11022 14728 11027 14784
rect 9121 14726 11027 14728
rect 9121 14723 9187 14726
rect 10961 14723 11027 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 8201 14652 8267 14653
rect 8150 14650 8156 14652
rect 8110 14590 8156 14650
rect 8220 14648 8267 14652
rect 8262 14592 8267 14648
rect 8150 14588 8156 14590
rect 8220 14588 8267 14592
rect 8201 14587 8267 14588
rect 9397 14650 9463 14653
rect 12801 14650 12867 14653
rect 9397 14648 12867 14650
rect 9397 14592 9402 14648
rect 9458 14592 12806 14648
rect 12862 14592 12867 14648
rect 9397 14590 12867 14592
rect 9397 14587 9463 14590
rect 12801 14587 12867 14590
rect 0 14514 800 14544
rect 1485 14514 1551 14517
rect 0 14512 1551 14514
rect 0 14456 1490 14512
rect 1546 14456 1551 14512
rect 0 14454 1551 14456
rect 0 14424 800 14454
rect 1485 14451 1551 14454
rect 3366 14452 3372 14516
rect 3436 14514 3442 14516
rect 6913 14514 6979 14517
rect 3436 14512 6979 14514
rect 3436 14456 6918 14512
rect 6974 14456 6979 14512
rect 3436 14454 6979 14456
rect 3436 14452 3442 14454
rect 6913 14451 6979 14454
rect 7281 14514 7347 14517
rect 7598 14514 7604 14516
rect 7281 14512 7604 14514
rect 7281 14456 7286 14512
rect 7342 14456 7604 14512
rect 7281 14454 7604 14456
rect 7281 14451 7347 14454
rect 7598 14452 7604 14454
rect 7668 14452 7674 14516
rect 8937 14514 9003 14517
rect 9305 14514 9371 14517
rect 8937 14512 9371 14514
rect 8937 14456 8942 14512
rect 8998 14456 9310 14512
rect 9366 14456 9371 14512
rect 8937 14454 9371 14456
rect 8937 14451 9003 14454
rect 9305 14451 9371 14454
rect 9581 14514 9647 14517
rect 16205 14514 16271 14517
rect 9581 14512 16271 14514
rect 9581 14456 9586 14512
rect 9642 14456 16210 14512
rect 16266 14456 16271 14512
rect 9581 14454 16271 14456
rect 9581 14451 9647 14454
rect 16205 14451 16271 14454
rect 21449 14514 21515 14517
rect 22200 14514 23000 14544
rect 21449 14512 23000 14514
rect 21449 14456 21454 14512
rect 21510 14456 23000 14512
rect 21449 14454 23000 14456
rect 21449 14451 21515 14454
rect 22200 14424 23000 14454
rect 933 14378 999 14381
rect 10777 14378 10843 14381
rect 933 14376 10843 14378
rect 933 14320 938 14376
rect 994 14320 10782 14376
rect 10838 14320 10843 14376
rect 933 14318 10843 14320
rect 933 14315 999 14318
rect 10777 14315 10843 14318
rect 11053 14378 11119 14381
rect 16389 14378 16455 14381
rect 11053 14376 16455 14378
rect 11053 14320 11058 14376
rect 11114 14320 16394 14376
rect 16450 14320 16455 14376
rect 11053 14318 16455 14320
rect 11053 14315 11119 14318
rect 2037 14242 2103 14245
rect 2262 14242 2268 14244
rect 2037 14240 2268 14242
rect 2037 14184 2042 14240
rect 2098 14184 2268 14240
rect 2037 14182 2268 14184
rect 2037 14179 2103 14182
rect 2262 14180 2268 14182
rect 2332 14180 2338 14244
rect 9029 14242 9095 14245
rect 11056 14242 11116 14315
rect 11884 14245 11944 14318
rect 16389 14315 16455 14318
rect 9029 14240 11116 14242
rect 9029 14184 9034 14240
rect 9090 14184 11116 14240
rect 9029 14182 11116 14184
rect 11881 14240 11947 14245
rect 11881 14184 11886 14240
rect 11942 14184 11947 14240
rect 9029 14179 9095 14182
rect 11881 14179 11947 14184
rect 13813 14242 13879 14245
rect 14365 14244 14431 14245
rect 14365 14242 14412 14244
rect 13813 14240 14412 14242
rect 13813 14184 13818 14240
rect 13874 14184 14370 14240
rect 13813 14182 14412 14184
rect 13813 14179 13879 14182
rect 14365 14180 14412 14182
rect 14476 14180 14482 14244
rect 14365 14179 14431 14180
rect 6144 14176 6460 14177
rect 0 14106 800 14136
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 1485 14106 1551 14109
rect 0 14104 1551 14106
rect 0 14048 1490 14104
rect 1546 14048 1551 14104
rect 0 14046 1551 14048
rect 0 14016 800 14046
rect 1485 14043 1551 14046
rect 7373 14106 7439 14109
rect 9765 14106 9831 14109
rect 7373 14104 9831 14106
rect 7373 14048 7378 14104
rect 7434 14048 9770 14104
rect 9826 14048 9831 14104
rect 7373 14046 9831 14048
rect 7373 14043 7439 14046
rect 9765 14043 9831 14046
rect 11789 14106 11855 14109
rect 19517 14108 19583 14109
rect 14406 14106 14412 14108
rect 11789 14104 14412 14106
rect 11789 14048 11794 14104
rect 11850 14048 14412 14104
rect 11789 14046 14412 14048
rect 11789 14043 11855 14046
rect 14406 14044 14412 14046
rect 14476 14044 14482 14108
rect 19517 14104 19564 14108
rect 19628 14106 19634 14108
rect 22200 14106 23000 14136
rect 19517 14048 19522 14104
rect 19517 14044 19564 14048
rect 19628 14046 19674 14106
rect 19628 14044 19634 14046
rect 19517 14043 19583 14044
rect 22142 14016 23000 14106
rect 1945 13970 2011 13973
rect 4061 13970 4127 13973
rect 9673 13970 9739 13973
rect 1945 13968 9739 13970
rect 1945 13912 1950 13968
rect 2006 13912 4066 13968
rect 4122 13912 9678 13968
rect 9734 13912 9739 13968
rect 1945 13910 9739 13912
rect 1945 13907 2011 13910
rect 4061 13907 4127 13910
rect 9673 13907 9739 13910
rect 10317 13970 10383 13973
rect 16113 13970 16179 13973
rect 20805 13970 20871 13973
rect 10317 13968 16179 13970
rect 10317 13912 10322 13968
rect 10378 13912 16118 13968
rect 16174 13912 16179 13968
rect 10317 13910 16179 13912
rect 10317 13907 10383 13910
rect 16113 13907 16179 13910
rect 16254 13968 20871 13970
rect 16254 13912 20810 13968
rect 20866 13912 20871 13968
rect 16254 13910 20871 13912
rect 4153 13834 4219 13837
rect 4613 13834 4679 13837
rect 8293 13834 8359 13837
rect 4153 13832 8359 13834
rect 4153 13776 4158 13832
rect 4214 13776 4618 13832
rect 4674 13776 8298 13832
rect 8354 13776 8359 13832
rect 4153 13774 8359 13776
rect 4153 13771 4219 13774
rect 4613 13771 4679 13774
rect 8293 13771 8359 13774
rect 8937 13834 9003 13837
rect 9438 13834 9444 13836
rect 8937 13832 9444 13834
rect 8937 13776 8942 13832
rect 8998 13776 9444 13832
rect 8937 13774 9444 13776
rect 8937 13771 9003 13774
rect 9438 13772 9444 13774
rect 9508 13834 9514 13836
rect 10501 13834 10567 13837
rect 9508 13832 10567 13834
rect 9508 13776 10506 13832
rect 10562 13776 10567 13832
rect 9508 13774 10567 13776
rect 9508 13772 9514 13774
rect 10501 13771 10567 13774
rect 10777 13834 10843 13837
rect 10777 13832 10978 13834
rect 10777 13776 10782 13832
rect 10838 13776 10978 13832
rect 10777 13774 10978 13776
rect 10777 13771 10843 13774
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 5574 13636 5580 13700
rect 5644 13698 5650 13700
rect 6545 13698 6611 13701
rect 5644 13696 6611 13698
rect 5644 13640 6550 13696
rect 6606 13640 6611 13696
rect 5644 13638 6611 13640
rect 5644 13636 5650 13638
rect 6545 13635 6611 13638
rect 10041 13698 10107 13701
rect 10777 13698 10843 13701
rect 10041 13696 10843 13698
rect 10041 13640 10046 13696
rect 10102 13640 10782 13696
rect 10838 13640 10843 13696
rect 10041 13638 10843 13640
rect 10918 13698 10978 13774
rect 11094 13772 11100 13836
rect 11164 13834 11170 13836
rect 11789 13834 11855 13837
rect 12249 13836 12315 13837
rect 12198 13834 12204 13836
rect 11164 13832 11855 13834
rect 11164 13776 11794 13832
rect 11850 13776 11855 13832
rect 11164 13774 11855 13776
rect 12158 13774 12204 13834
rect 12268 13832 12315 13836
rect 12310 13776 12315 13832
rect 11164 13772 11170 13774
rect 11789 13771 11855 13774
rect 12198 13772 12204 13774
rect 12268 13772 12315 13776
rect 12249 13771 12315 13772
rect 13445 13836 13511 13837
rect 13445 13832 13492 13836
rect 13556 13834 13562 13836
rect 14549 13834 14615 13837
rect 14958 13834 14964 13836
rect 13445 13776 13450 13832
rect 13445 13772 13492 13776
rect 13556 13774 13602 13834
rect 14549 13832 14964 13834
rect 14549 13776 14554 13832
rect 14610 13776 14964 13832
rect 14549 13774 14964 13776
rect 13556 13772 13562 13774
rect 13445 13771 13511 13772
rect 14549 13771 14615 13774
rect 14958 13772 14964 13774
rect 15028 13834 15034 13836
rect 16254 13834 16314 13910
rect 20805 13907 20871 13910
rect 21449 13970 21515 13973
rect 22142 13970 22202 14016
rect 21449 13968 22202 13970
rect 21449 13912 21454 13968
rect 21510 13912 22202 13968
rect 21449 13910 22202 13912
rect 21449 13907 21515 13910
rect 15028 13774 16314 13834
rect 15028 13772 15034 13774
rect 19926 13772 19932 13836
rect 19996 13834 20002 13836
rect 20345 13834 20411 13837
rect 19996 13832 20411 13834
rect 19996 13776 20350 13832
rect 20406 13776 20411 13832
rect 19996 13774 20411 13776
rect 19996 13772 20002 13774
rect 20345 13771 20411 13774
rect 11513 13698 11579 13701
rect 12433 13698 12499 13701
rect 10918 13696 11579 13698
rect 10918 13640 11518 13696
rect 11574 13640 11579 13696
rect 10918 13638 11579 13640
rect 10041 13635 10107 13638
rect 10777 13635 10843 13638
rect 11513 13635 11579 13638
rect 12390 13696 12499 13698
rect 12390 13640 12438 13696
rect 12494 13640 12499 13696
rect 12390 13635 12499 13640
rect 21449 13698 21515 13701
rect 22200 13698 23000 13728
rect 21449 13696 23000 13698
rect 21449 13640 21454 13696
rect 21510 13640 23000 13696
rect 21449 13638 23000 13640
rect 21449 13635 21515 13638
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 1342 13500 1348 13564
rect 1412 13562 1418 13564
rect 1412 13502 2790 13562
rect 1412 13500 1418 13502
rect 2730 13426 2790 13502
rect 4102 13500 4108 13564
rect 4172 13562 4178 13564
rect 8569 13562 8635 13565
rect 12390 13562 12450 13635
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 22200 13608 23000 13638
rect 19139 13567 19455 13568
rect 4172 13560 8635 13562
rect 4172 13504 8574 13560
rect 8630 13504 8635 13560
rect 4172 13502 8635 13504
rect 4172 13500 4178 13502
rect 8569 13499 8635 13502
rect 9262 13502 12450 13562
rect 20621 13562 20687 13565
rect 21030 13562 21036 13564
rect 20621 13560 21036 13562
rect 20621 13504 20626 13560
rect 20682 13504 21036 13560
rect 20621 13502 21036 13504
rect 9262 13426 9322 13502
rect 20621 13499 20687 13502
rect 21030 13500 21036 13502
rect 21100 13500 21106 13564
rect 11973 13426 12039 13429
rect 2730 13366 9322 13426
rect 9446 13424 12039 13426
rect 9446 13368 11978 13424
rect 12034 13368 12039 13424
rect 9446 13366 12039 13368
rect 0 13290 800 13320
rect 1485 13290 1551 13293
rect 0 13288 1551 13290
rect 0 13232 1490 13288
rect 1546 13232 1551 13288
rect 0 13230 1551 13232
rect 0 13200 800 13230
rect 1485 13227 1551 13230
rect 2814 13228 2820 13292
rect 2884 13290 2890 13292
rect 9446 13290 9506 13366
rect 11973 13363 12039 13366
rect 12249 13426 12315 13429
rect 12566 13426 12572 13428
rect 12249 13424 12572 13426
rect 12249 13368 12254 13424
rect 12310 13368 12572 13424
rect 12249 13366 12572 13368
rect 12249 13363 12315 13366
rect 12566 13364 12572 13366
rect 12636 13364 12642 13428
rect 14273 13426 14339 13429
rect 21633 13426 21699 13429
rect 14273 13424 21699 13426
rect 14273 13368 14278 13424
rect 14334 13368 21638 13424
rect 21694 13368 21699 13424
rect 14273 13366 21699 13368
rect 14273 13363 14339 13366
rect 21633 13363 21699 13366
rect 2884 13230 9506 13290
rect 2884 13228 2890 13230
rect 10174 13228 10180 13292
rect 10244 13290 10250 13292
rect 10317 13290 10383 13293
rect 10593 13290 10659 13293
rect 10244 13288 10659 13290
rect 10244 13232 10322 13288
rect 10378 13232 10598 13288
rect 10654 13232 10659 13288
rect 10244 13230 10659 13232
rect 10244 13228 10250 13230
rect 10317 13227 10383 13230
rect 10593 13227 10659 13230
rect 11053 13290 11119 13293
rect 16062 13290 16068 13292
rect 11053 13288 16068 13290
rect 11053 13232 11058 13288
rect 11114 13232 16068 13288
rect 11053 13230 16068 13232
rect 11053 13227 11119 13230
rect 16062 13228 16068 13230
rect 16132 13228 16138 13292
rect 19558 13228 19564 13292
rect 19628 13290 19634 13292
rect 19701 13290 19767 13293
rect 19628 13288 19767 13290
rect 19628 13232 19706 13288
rect 19762 13232 19767 13288
rect 19628 13230 19767 13232
rect 19628 13228 19634 13230
rect 19701 13227 19767 13230
rect 21449 13290 21515 13293
rect 22200 13290 23000 13320
rect 21449 13288 23000 13290
rect 21449 13232 21454 13288
rect 21510 13232 23000 13288
rect 21449 13230 23000 13232
rect 21449 13227 21515 13230
rect 22200 13200 23000 13230
rect 2405 13154 2471 13157
rect 4061 13154 4127 13157
rect 2405 13152 4127 13154
rect 2405 13096 2410 13152
rect 2466 13096 4066 13152
rect 4122 13096 4127 13152
rect 2405 13094 4127 13096
rect 2405 13091 2471 13094
rect 4061 13091 4127 13094
rect 4337 13154 4403 13157
rect 5441 13154 5507 13157
rect 4337 13152 5507 13154
rect 4337 13096 4342 13152
rect 4398 13096 5446 13152
rect 5502 13096 5507 13152
rect 4337 13094 5507 13096
rect 4337 13091 4403 13094
rect 5441 13091 5507 13094
rect 6637 13154 6703 13157
rect 7782 13154 7788 13156
rect 6637 13152 7788 13154
rect 6637 13096 6642 13152
rect 6698 13096 7788 13152
rect 6637 13094 7788 13096
rect 6637 13091 6703 13094
rect 7782 13092 7788 13094
rect 7852 13092 7858 13156
rect 8293 13154 8359 13157
rect 10685 13154 10751 13157
rect 8293 13152 10751 13154
rect 8293 13096 8298 13152
rect 8354 13096 10690 13152
rect 10746 13096 10751 13152
rect 8293 13094 10751 13096
rect 8293 13091 8359 13094
rect 10685 13091 10751 13094
rect 12157 13154 12223 13157
rect 12157 13152 14658 13154
rect 12157 13096 12162 13152
rect 12218 13096 14658 13152
rect 12157 13094 14658 13096
rect 12157 13091 12223 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 3182 12956 3188 13020
rect 3252 13018 3258 13020
rect 4102 13018 4108 13020
rect 3252 12958 4108 13018
rect 3252 12956 3258 12958
rect 4102 12956 4108 12958
rect 4172 12956 4178 13020
rect 6862 12956 6868 13020
rect 6932 13018 6938 13020
rect 8017 13018 8083 13021
rect 10358 13018 10364 13020
rect 6932 13016 10364 13018
rect 6932 12960 8022 13016
rect 8078 12960 10364 13016
rect 6932 12958 10364 12960
rect 6932 12956 6938 12958
rect 8017 12955 8083 12958
rect 10358 12956 10364 12958
rect 10428 12956 10434 13020
rect 12934 12956 12940 13020
rect 13004 13018 13010 13020
rect 13353 13018 13419 13021
rect 13004 13016 13419 13018
rect 13004 12960 13358 13016
rect 13414 12960 13419 13016
rect 13004 12958 13419 12960
rect 13004 12956 13010 12958
rect 13353 12955 13419 12958
rect 0 12882 800 12912
rect 1853 12882 1919 12885
rect 0 12880 1919 12882
rect 0 12824 1858 12880
rect 1914 12824 1919 12880
rect 0 12822 1919 12824
rect 0 12792 800 12822
rect 1853 12819 1919 12822
rect 4153 12882 4219 12885
rect 11789 12882 11855 12885
rect 4153 12880 11855 12882
rect 4153 12824 4158 12880
rect 4214 12824 11794 12880
rect 11850 12824 11855 12880
rect 4153 12822 11855 12824
rect 4153 12819 4219 12822
rect 11789 12819 11855 12822
rect 11973 12882 12039 12885
rect 12525 12882 12591 12885
rect 11973 12880 12591 12882
rect 11973 12824 11978 12880
rect 12034 12824 12530 12880
rect 12586 12824 12591 12880
rect 11973 12822 12591 12824
rect 11973 12819 12039 12822
rect 12525 12819 12591 12822
rect 13629 12884 13695 12885
rect 13629 12880 13676 12884
rect 13740 12882 13746 12884
rect 14598 12882 14658 13094
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 16982 12882 16988 12884
rect 13629 12824 13634 12880
rect 13629 12820 13676 12824
rect 13740 12822 13786 12882
rect 14598 12822 16988 12882
rect 13740 12820 13746 12822
rect 16982 12820 16988 12822
rect 17052 12820 17058 12884
rect 21081 12882 21147 12885
rect 22200 12882 23000 12912
rect 21081 12880 23000 12882
rect 21081 12824 21086 12880
rect 21142 12824 23000 12880
rect 21081 12822 23000 12824
rect 13629 12819 13695 12820
rect 21081 12819 21147 12822
rect 22200 12792 23000 12822
rect 974 12684 980 12748
rect 1044 12746 1050 12748
rect 4613 12746 4679 12749
rect 7005 12746 7071 12749
rect 1044 12686 3986 12746
rect 1044 12684 1050 12686
rect 3545 12544 3861 12545
rect 0 12474 800 12504
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 1485 12474 1551 12477
rect 0 12472 1551 12474
rect 0 12416 1490 12472
rect 1546 12416 1551 12472
rect 0 12414 1551 12416
rect 3926 12474 3986 12686
rect 4613 12744 7071 12746
rect 4613 12688 4618 12744
rect 4674 12688 7010 12744
rect 7066 12688 7071 12744
rect 4613 12686 7071 12688
rect 4613 12683 4679 12686
rect 7005 12683 7071 12686
rect 7598 12684 7604 12748
rect 7668 12746 7674 12748
rect 8017 12746 8083 12749
rect 14549 12746 14615 12749
rect 7668 12744 14615 12746
rect 7668 12688 8022 12744
rect 8078 12688 14554 12744
rect 14610 12688 14615 12744
rect 7668 12686 14615 12688
rect 7668 12684 7674 12686
rect 8017 12683 8083 12686
rect 14549 12683 14615 12686
rect 17217 12746 17283 12749
rect 18965 12746 19031 12749
rect 17217 12744 19031 12746
rect 17217 12688 17222 12744
rect 17278 12688 18970 12744
rect 19026 12688 19031 12744
rect 17217 12686 19031 12688
rect 17217 12683 17283 12686
rect 18965 12683 19031 12686
rect 4705 12610 4771 12613
rect 4981 12610 5047 12613
rect 8201 12610 8267 12613
rect 4705 12608 8267 12610
rect 4705 12552 4710 12608
rect 4766 12552 4986 12608
rect 5042 12552 8206 12608
rect 8262 12552 8267 12608
rect 4705 12550 8267 12552
rect 4705 12547 4771 12550
rect 4981 12547 5047 12550
rect 8201 12547 8267 12550
rect 9213 12610 9279 12613
rect 13813 12610 13879 12613
rect 9213 12608 13879 12610
rect 9213 12552 9218 12608
rect 9274 12552 13818 12608
rect 13874 12552 13879 12608
rect 9213 12550 13879 12552
rect 9213 12547 9279 12550
rect 13813 12547 13879 12550
rect 16757 12610 16823 12613
rect 17718 12610 17724 12612
rect 16757 12608 17724 12610
rect 16757 12552 16762 12608
rect 16818 12552 17724 12608
rect 16757 12550 17724 12552
rect 16757 12547 16823 12550
rect 17718 12548 17724 12550
rect 17788 12548 17794 12612
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 8569 12474 8635 12477
rect 3926 12472 8635 12474
rect 3926 12416 8574 12472
rect 8630 12416 8635 12472
rect 3926 12414 8635 12416
rect 0 12384 800 12414
rect 1485 12411 1551 12414
rect 8569 12411 8635 12414
rect 9489 12474 9555 12477
rect 10593 12476 10659 12477
rect 9622 12474 9628 12476
rect 9489 12472 9628 12474
rect 9489 12416 9494 12472
rect 9550 12416 9628 12472
rect 9489 12414 9628 12416
rect 9489 12411 9555 12414
rect 9622 12412 9628 12414
rect 9692 12412 9698 12476
rect 10542 12412 10548 12476
rect 10612 12474 10659 12476
rect 10777 12474 10843 12477
rect 11973 12476 12039 12477
rect 11973 12474 12020 12476
rect 10612 12472 10704 12474
rect 10654 12416 10704 12472
rect 10612 12414 10704 12416
rect 10777 12472 11116 12474
rect 10777 12416 10782 12472
rect 10838 12416 11116 12472
rect 10777 12414 11116 12416
rect 11928 12472 12020 12474
rect 11928 12416 11978 12472
rect 11928 12414 12020 12416
rect 10612 12412 10659 12414
rect 10593 12411 10659 12412
rect 10777 12411 10843 12414
rect 1301 12338 1367 12341
rect 7097 12338 7163 12341
rect 7230 12338 7236 12340
rect 1301 12336 6792 12338
rect 1301 12280 1306 12336
rect 1362 12280 6792 12336
rect 1301 12278 6792 12280
rect 1301 12275 1367 12278
rect 2313 12202 2379 12205
rect 6732 12202 6792 12278
rect 7097 12336 7236 12338
rect 7097 12280 7102 12336
rect 7158 12280 7236 12336
rect 7097 12278 7236 12280
rect 7097 12275 7163 12278
rect 7230 12276 7236 12278
rect 7300 12276 7306 12340
rect 7414 12276 7420 12340
rect 7484 12338 7490 12340
rect 7741 12338 7807 12341
rect 7484 12336 7807 12338
rect 7484 12280 7746 12336
rect 7802 12280 7807 12336
rect 7484 12278 7807 12280
rect 7484 12276 7490 12278
rect 7741 12275 7807 12278
rect 7966 12276 7972 12340
rect 8036 12338 8042 12340
rect 9857 12338 9923 12341
rect 8036 12336 9923 12338
rect 8036 12280 9862 12336
rect 9918 12280 9923 12336
rect 8036 12278 9923 12280
rect 8036 12276 8042 12278
rect 9857 12275 9923 12278
rect 9990 12276 9996 12340
rect 10060 12338 10066 12340
rect 10225 12338 10291 12341
rect 10060 12336 10291 12338
rect 10060 12280 10230 12336
rect 10286 12280 10291 12336
rect 10060 12278 10291 12280
rect 11056 12338 11116 12414
rect 11973 12412 12020 12414
rect 12084 12412 12090 12476
rect 21449 12474 21515 12477
rect 22200 12474 23000 12504
rect 21449 12472 23000 12474
rect 21449 12416 21454 12472
rect 21510 12416 23000 12472
rect 21449 12414 23000 12416
rect 11973 12411 12039 12412
rect 21449 12411 21515 12414
rect 22200 12384 23000 12414
rect 11056 12278 12450 12338
rect 10060 12276 10066 12278
rect 10225 12275 10291 12278
rect 10869 12202 10935 12205
rect 11973 12202 12039 12205
rect 2313 12200 6608 12202
rect 2313 12144 2318 12200
rect 2374 12144 6608 12200
rect 2313 12142 6608 12144
rect 6732 12200 10935 12202
rect 6732 12144 10874 12200
rect 10930 12144 10935 12200
rect 6732 12142 10935 12144
rect 2313 12139 2379 12142
rect 0 12066 800 12096
rect 1853 12066 1919 12069
rect 0 12064 1919 12066
rect 0 12008 1858 12064
rect 1914 12008 1919 12064
rect 0 12006 1919 12008
rect 0 11976 800 12006
rect 1853 12003 1919 12006
rect 3693 12066 3759 12069
rect 5257 12066 5323 12069
rect 3693 12064 5323 12066
rect 3693 12008 3698 12064
rect 3754 12008 5262 12064
rect 5318 12008 5323 12064
rect 3693 12006 5323 12008
rect 6548 12066 6608 12142
rect 10869 12139 10935 12142
rect 11102 12200 12039 12202
rect 11102 12144 11978 12200
rect 12034 12144 12039 12200
rect 11102 12142 12039 12144
rect 12390 12202 12450 12278
rect 12934 12276 12940 12340
rect 13004 12338 13010 12340
rect 13004 12278 15762 12338
rect 13004 12276 13010 12278
rect 13445 12202 13511 12205
rect 15009 12202 15075 12205
rect 12390 12200 13511 12202
rect 12390 12144 13450 12200
rect 13506 12144 13511 12200
rect 12390 12142 13511 12144
rect 11102 12066 11162 12142
rect 11973 12139 12039 12142
rect 13445 12139 13511 12142
rect 13724 12200 15075 12202
rect 13724 12144 15014 12200
rect 15070 12144 15075 12200
rect 13724 12142 15075 12144
rect 15702 12202 15762 12278
rect 15878 12276 15884 12340
rect 15948 12338 15954 12340
rect 17861 12338 17927 12341
rect 20805 12338 20871 12341
rect 15948 12336 20871 12338
rect 15948 12280 17866 12336
rect 17922 12280 20810 12336
rect 20866 12280 20871 12336
rect 15948 12278 20871 12280
rect 15948 12276 15954 12278
rect 17861 12275 17927 12278
rect 20805 12275 20871 12278
rect 21449 12202 21515 12205
rect 15702 12142 18154 12202
rect 13724 12069 13784 12142
rect 15009 12139 15075 12142
rect 13721 12066 13787 12069
rect 6548 12006 11162 12066
rect 12390 12064 13787 12066
rect 12390 12008 13726 12064
rect 13782 12008 13787 12064
rect 12390 12006 13787 12008
rect 3693 12003 3759 12006
rect 5257 12003 5323 12006
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 7005 11932 7071 11933
rect 7005 11930 7052 11932
rect 6960 11928 7052 11930
rect 6960 11872 7010 11928
rect 6960 11870 7052 11872
rect 7005 11868 7052 11870
rect 7116 11868 7122 11932
rect 7230 11868 7236 11932
rect 7300 11930 7306 11932
rect 8017 11930 8083 11933
rect 8569 11932 8635 11933
rect 8518 11930 8524 11932
rect 7300 11928 8083 11930
rect 7300 11872 8022 11928
rect 8078 11872 8083 11928
rect 7300 11870 8083 11872
rect 8478 11870 8524 11930
rect 8588 11928 8635 11932
rect 8630 11872 8635 11928
rect 7300 11868 7306 11870
rect 7005 11867 7071 11868
rect 8017 11867 8083 11870
rect 8518 11868 8524 11870
rect 8588 11868 8635 11872
rect 8569 11867 8635 11868
rect 9029 11930 9095 11933
rect 9254 11930 9260 11932
rect 9029 11928 9260 11930
rect 9029 11872 9034 11928
rect 9090 11872 9260 11928
rect 9029 11870 9260 11872
rect 9029 11867 9095 11870
rect 9254 11868 9260 11870
rect 9324 11868 9330 11932
rect 9400 11870 9874 11930
rect 6361 11794 6427 11797
rect 9400 11794 9460 11870
rect 6361 11792 9460 11794
rect 6361 11736 6366 11792
rect 6422 11736 9460 11792
rect 6361 11734 9460 11736
rect 9814 11794 9874 11870
rect 10542 11868 10548 11932
rect 10612 11930 10618 11932
rect 10961 11930 11027 11933
rect 12390 11930 12450 12006
rect 13721 12003 13787 12006
rect 14406 12004 14412 12068
rect 14476 12066 14482 12068
rect 14774 12066 14780 12068
rect 14476 12006 14780 12066
rect 14476 12004 14482 12006
rect 14774 12004 14780 12006
rect 14844 12004 14850 12068
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 10612 11928 11027 11930
rect 10612 11872 10966 11928
rect 11022 11872 11027 11928
rect 10612 11870 11027 11872
rect 10612 11868 10618 11870
rect 10961 11867 11027 11870
rect 11838 11870 12450 11930
rect 13261 11930 13327 11933
rect 13813 11930 13879 11933
rect 14406 11930 14412 11932
rect 13261 11928 13554 11930
rect 13261 11872 13266 11928
rect 13322 11872 13554 11928
rect 13261 11870 13554 11872
rect 11838 11794 11898 11870
rect 13261 11867 13327 11870
rect 13494 11797 13554 11870
rect 13813 11928 14412 11930
rect 13813 11872 13818 11928
rect 13874 11872 14412 11928
rect 13813 11870 14412 11872
rect 13813 11867 13879 11870
rect 14406 11868 14412 11870
rect 14476 11868 14482 11932
rect 14641 11930 14707 11933
rect 15326 11930 15332 11932
rect 14641 11928 15332 11930
rect 14641 11872 14646 11928
rect 14702 11872 15332 11928
rect 14641 11870 15332 11872
rect 14641 11867 14707 11870
rect 15326 11868 15332 11870
rect 15396 11868 15402 11932
rect 9814 11734 11898 11794
rect 6361 11731 6427 11734
rect 12014 11732 12020 11796
rect 12084 11794 12090 11796
rect 12249 11794 12315 11797
rect 12084 11792 12315 11794
rect 12084 11736 12254 11792
rect 12310 11736 12315 11792
rect 12084 11734 12315 11736
rect 12084 11732 12090 11734
rect 12249 11731 12315 11734
rect 12382 11732 12388 11796
rect 12452 11794 12458 11796
rect 12525 11794 12591 11797
rect 12452 11792 12591 11794
rect 12452 11736 12530 11792
rect 12586 11736 12591 11792
rect 12452 11734 12591 11736
rect 13494 11792 13603 11797
rect 17033 11794 17099 11797
rect 13494 11736 13542 11792
rect 13598 11736 13603 11792
rect 13494 11734 13603 11736
rect 12452 11732 12458 11734
rect 12525 11731 12591 11734
rect 13537 11731 13603 11734
rect 13678 11792 17099 11794
rect 13678 11736 17038 11792
rect 17094 11736 17099 11792
rect 13678 11734 17099 11736
rect 18094 11794 18154 12142
rect 21449 12200 22202 12202
rect 21449 12144 21454 12200
rect 21510 12144 22202 12200
rect 21449 12142 22202 12144
rect 21449 12139 21515 12142
rect 22142 12096 22202 12142
rect 22142 12006 23000 12096
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 22200 11976 23000 12006
rect 21738 11935 22054 11936
rect 18229 11794 18295 11797
rect 18094 11792 18295 11794
rect 18094 11736 18234 11792
rect 18290 11736 18295 11792
rect 18094 11734 18295 11736
rect 0 11658 800 11688
rect 2221 11658 2287 11661
rect 5574 11658 5580 11660
rect 0 11656 2287 11658
rect 0 11600 2226 11656
rect 2282 11600 2287 11656
rect 0 11598 2287 11600
rect 0 11568 800 11598
rect 2221 11595 2287 11598
rect 2408 11598 5580 11658
rect 1669 11388 1735 11389
rect 1669 11386 1716 11388
rect 1624 11384 1716 11386
rect 1624 11328 1674 11384
rect 1624 11326 1716 11328
rect 1669 11324 1716 11326
rect 1780 11324 1786 11388
rect 2037 11386 2103 11389
rect 2408 11386 2468 11598
rect 5574 11596 5580 11598
rect 5644 11596 5650 11660
rect 7097 11658 7163 11661
rect 7649 11658 7715 11661
rect 13678 11658 13738 11734
rect 17033 11731 17099 11734
rect 18229 11731 18295 11734
rect 7097 11656 13738 11658
rect 7097 11600 7102 11656
rect 7158 11600 7654 11656
rect 7710 11600 13738 11656
rect 7097 11598 13738 11600
rect 13813 11658 13879 11661
rect 14590 11658 14596 11660
rect 13813 11656 14596 11658
rect 13813 11600 13818 11656
rect 13874 11600 14596 11656
rect 13813 11598 14596 11600
rect 7097 11595 7163 11598
rect 7649 11595 7715 11598
rect 13813 11595 13879 11598
rect 14590 11596 14596 11598
rect 14660 11596 14666 11660
rect 16573 11658 16639 11661
rect 17166 11658 17172 11660
rect 16573 11656 17172 11658
rect 16573 11600 16578 11656
rect 16634 11600 17172 11656
rect 16573 11598 17172 11600
rect 16573 11595 16639 11598
rect 17166 11596 17172 11598
rect 17236 11596 17242 11660
rect 17401 11658 17467 11661
rect 17358 11656 17467 11658
rect 17358 11600 17406 11656
rect 17462 11600 17467 11656
rect 17358 11595 17467 11600
rect 18638 11596 18644 11660
rect 18708 11658 18714 11660
rect 20713 11658 20779 11661
rect 18708 11656 20779 11658
rect 18708 11600 20718 11656
rect 20774 11600 20779 11656
rect 18708 11598 20779 11600
rect 18708 11596 18714 11598
rect 20713 11595 20779 11598
rect 21541 11658 21607 11661
rect 22200 11658 23000 11688
rect 21541 11656 23000 11658
rect 21541 11600 21546 11656
rect 21602 11600 23000 11656
rect 21541 11598 23000 11600
rect 21541 11595 21607 11598
rect 4470 11460 4476 11524
rect 4540 11522 4546 11524
rect 7966 11522 7972 11524
rect 4540 11462 7972 11522
rect 4540 11460 4546 11462
rect 7966 11460 7972 11462
rect 8036 11460 8042 11524
rect 11605 11522 11671 11525
rect 12014 11522 12020 11524
rect 11605 11520 12020 11522
rect 11605 11464 11610 11520
rect 11666 11464 12020 11520
rect 11605 11462 12020 11464
rect 11605 11459 11671 11462
rect 12014 11460 12020 11462
rect 12084 11460 12090 11524
rect 15326 11460 15332 11524
rect 15396 11522 15402 11524
rect 16389 11522 16455 11525
rect 15396 11520 16455 11522
rect 15396 11464 16394 11520
rect 16450 11464 16455 11520
rect 15396 11462 16455 11464
rect 15396 11460 15402 11462
rect 16389 11459 16455 11462
rect 17166 11460 17172 11524
rect 17236 11522 17242 11524
rect 17358 11522 17418 11595
rect 22200 11568 23000 11598
rect 17236 11462 17418 11522
rect 17236 11460 17242 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 19139 11391 19455 11392
rect 5901 11386 5967 11389
rect 2037 11384 2468 11386
rect 2037 11328 2042 11384
rect 2098 11328 2468 11384
rect 2037 11326 2468 11328
rect 3926 11384 5967 11386
rect 3926 11328 5906 11384
rect 5962 11328 5967 11384
rect 3926 11326 5967 11328
rect 1669 11323 1735 11324
rect 2037 11323 2103 11326
rect 0 11250 800 11280
rect 1485 11250 1551 11253
rect 3926 11252 3986 11326
rect 5901 11323 5967 11326
rect 6085 11386 6151 11389
rect 6678 11386 6684 11388
rect 6085 11384 6684 11386
rect 6085 11328 6090 11384
rect 6146 11328 6684 11384
rect 6085 11326 6684 11328
rect 6085 11323 6151 11326
rect 6678 11324 6684 11326
rect 6748 11324 6754 11388
rect 7373 11386 7439 11389
rect 7966 11386 7972 11388
rect 7373 11384 7972 11386
rect 7373 11328 7378 11384
rect 7434 11328 7972 11384
rect 7373 11326 7972 11328
rect 7373 11323 7439 11326
rect 7966 11324 7972 11326
rect 8036 11386 8042 11388
rect 8569 11386 8635 11389
rect 13353 11388 13419 11389
rect 8036 11384 8635 11386
rect 8036 11328 8574 11384
rect 8630 11328 8635 11384
rect 8036 11326 8635 11328
rect 8036 11324 8042 11326
rect 8569 11323 8635 11326
rect 9622 11324 9628 11388
rect 9692 11386 9698 11388
rect 12934 11386 12940 11388
rect 9692 11326 12940 11386
rect 9692 11324 9698 11326
rect 12934 11324 12940 11326
rect 13004 11324 13010 11388
rect 13302 11324 13308 11388
rect 13372 11386 13419 11388
rect 13372 11384 13784 11386
rect 13414 11328 13784 11384
rect 13372 11326 13784 11328
rect 13372 11324 13419 11326
rect 13353 11323 13419 11324
rect 0 11248 1551 11250
rect 0 11192 1490 11248
rect 1546 11192 1551 11248
rect 0 11190 1551 11192
rect 0 11160 800 11190
rect 1485 11187 1551 11190
rect 3918 11188 3924 11252
rect 3988 11188 3994 11252
rect 4102 11188 4108 11252
rect 4172 11250 4178 11252
rect 8334 11250 8340 11252
rect 4172 11190 8340 11250
rect 4172 11188 4178 11190
rect 8334 11188 8340 11190
rect 8404 11250 8410 11252
rect 8569 11250 8635 11253
rect 8404 11248 8635 11250
rect 8404 11192 8574 11248
rect 8630 11192 8635 11248
rect 8404 11190 8635 11192
rect 8404 11188 8410 11190
rect 8569 11187 8635 11190
rect 8753 11250 8819 11253
rect 9305 11250 9371 11253
rect 8753 11248 9371 11250
rect 8753 11192 8758 11248
rect 8814 11192 9310 11248
rect 9366 11192 9371 11248
rect 8753 11190 9371 11192
rect 8753 11187 8819 11190
rect 9305 11187 9371 11190
rect 10726 11188 10732 11252
rect 10796 11250 10802 11252
rect 12382 11250 12388 11252
rect 10796 11190 12388 11250
rect 10796 11188 10802 11190
rect 12382 11188 12388 11190
rect 12452 11188 12458 11252
rect 12801 11250 12867 11253
rect 13261 11250 13327 11253
rect 12801 11248 13327 11250
rect 12801 11192 12806 11248
rect 12862 11192 13266 11248
rect 13322 11192 13327 11248
rect 12801 11190 13327 11192
rect 13724 11250 13784 11326
rect 15142 11250 15148 11252
rect 13724 11190 15148 11250
rect 12801 11187 12867 11190
rect 13261 11187 13327 11190
rect 15142 11188 15148 11190
rect 15212 11188 15218 11252
rect 18689 11250 18755 11253
rect 19742 11250 19748 11252
rect 18689 11248 19748 11250
rect 18689 11192 18694 11248
rect 18750 11192 19748 11248
rect 18689 11190 19748 11192
rect 18689 11187 18755 11190
rect 19742 11188 19748 11190
rect 19812 11188 19818 11252
rect 21081 11250 21147 11253
rect 22200 11250 23000 11280
rect 21081 11248 23000 11250
rect 21081 11192 21086 11248
rect 21142 11192 23000 11248
rect 21081 11190 23000 11192
rect 21081 11187 21147 11190
rect 22200 11160 23000 11190
rect 5165 11114 5231 11117
rect 5390 11114 5396 11116
rect 5165 11112 5396 11114
rect 5165 11056 5170 11112
rect 5226 11056 5396 11112
rect 5165 11054 5396 11056
rect 5165 11051 5231 11054
rect 5390 11052 5396 11054
rect 5460 11052 5466 11116
rect 5901 11114 5967 11117
rect 10041 11114 10107 11117
rect 5901 11112 10107 11114
rect 5901 11056 5906 11112
rect 5962 11056 10046 11112
rect 10102 11056 10107 11112
rect 5901 11054 10107 11056
rect 5901 11051 5967 11054
rect 10041 11051 10107 11054
rect 10225 11114 10291 11117
rect 12750 11114 12756 11116
rect 10225 11112 12756 11114
rect 10225 11056 10230 11112
rect 10286 11056 12756 11112
rect 10225 11054 12756 11056
rect 10225 11051 10291 11054
rect 12750 11052 12756 11054
rect 12820 11052 12826 11116
rect 13629 11114 13695 11117
rect 19926 11114 19932 11116
rect 13629 11112 19932 11114
rect 13629 11056 13634 11112
rect 13690 11056 19932 11112
rect 13629 11054 19932 11056
rect 13629 11051 13695 11054
rect 19926 11052 19932 11054
rect 19996 11052 20002 11116
rect 6870 10918 7160 10978
rect 6144 10912 6460 10913
rect 0 10842 800 10872
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 1853 10842 1919 10845
rect 6870 10842 6930 10918
rect 0 10840 1919 10842
rect 0 10784 1858 10840
rect 1914 10784 1919 10840
rect 0 10782 1919 10784
rect 0 10752 800 10782
rect 1853 10779 1919 10782
rect 6548 10782 6930 10842
rect 7100 10842 7160 10918
rect 8334 10916 8340 10980
rect 8404 10978 8410 10980
rect 10777 10978 10843 10981
rect 8404 10976 10843 10978
rect 8404 10920 10782 10976
rect 10838 10920 10843 10976
rect 8404 10918 10843 10920
rect 8404 10916 8410 10918
rect 10777 10915 10843 10918
rect 12525 10978 12591 10981
rect 13077 10978 13143 10981
rect 12525 10976 13143 10978
rect 12525 10920 12530 10976
rect 12586 10920 13082 10976
rect 13138 10920 13143 10976
rect 12525 10918 13143 10920
rect 12525 10915 12591 10918
rect 13077 10915 13143 10918
rect 17861 10978 17927 10981
rect 20713 10978 20779 10981
rect 17861 10976 20779 10978
rect 17861 10920 17866 10976
rect 17922 10920 20718 10976
rect 20774 10920 20779 10976
rect 17861 10918 20779 10920
rect 17861 10915 17927 10918
rect 20713 10915 20779 10918
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 8937 10842 9003 10845
rect 10869 10842 10935 10845
rect 7100 10782 8816 10842
rect 2037 10706 2103 10709
rect 5993 10708 6059 10709
rect 2037 10704 5136 10706
rect 2037 10648 2042 10704
rect 2098 10648 5136 10704
rect 2037 10646 5136 10648
rect 2037 10643 2103 10646
rect 5076 10570 5136 10646
rect 5942 10644 5948 10708
rect 6012 10706 6059 10708
rect 6177 10706 6243 10709
rect 6548 10706 6608 10782
rect 6012 10704 6104 10706
rect 6054 10648 6104 10704
rect 6012 10646 6104 10648
rect 6177 10704 6608 10706
rect 6177 10648 6182 10704
rect 6238 10648 6608 10704
rect 6177 10646 6608 10648
rect 7097 10706 7163 10709
rect 7414 10706 7420 10708
rect 7097 10704 7420 10706
rect 7097 10648 7102 10704
rect 7158 10648 7420 10704
rect 7097 10646 7420 10648
rect 6012 10644 6059 10646
rect 5993 10643 6059 10644
rect 6177 10643 6243 10646
rect 7097 10643 7163 10646
rect 7414 10644 7420 10646
rect 7484 10644 7490 10708
rect 7782 10644 7788 10708
rect 7852 10706 7858 10708
rect 8569 10706 8635 10709
rect 7852 10704 8635 10706
rect 7852 10648 8574 10704
rect 8630 10648 8635 10704
rect 7852 10646 8635 10648
rect 8756 10706 8816 10782
rect 8937 10840 10935 10842
rect 8937 10784 8942 10840
rect 8998 10784 10874 10840
rect 10930 10784 10935 10840
rect 8937 10782 10935 10784
rect 8937 10779 9003 10782
rect 10869 10779 10935 10782
rect 13261 10842 13327 10845
rect 14457 10842 14523 10845
rect 14590 10842 14596 10844
rect 13261 10840 14596 10842
rect 13261 10784 13266 10840
rect 13322 10784 14462 10840
rect 14518 10784 14596 10840
rect 13261 10782 14596 10784
rect 13261 10779 13327 10782
rect 14457 10779 14523 10782
rect 14590 10780 14596 10782
rect 14660 10780 14666 10844
rect 21030 10780 21036 10844
rect 21100 10842 21106 10844
rect 21173 10842 21239 10845
rect 22200 10842 23000 10872
rect 21100 10840 21239 10842
rect 21100 10784 21178 10840
rect 21234 10784 21239 10840
rect 21100 10782 21239 10784
rect 21100 10780 21106 10782
rect 21173 10779 21239 10782
rect 22142 10752 23000 10842
rect 11053 10706 11119 10709
rect 17033 10706 17099 10709
rect 8756 10704 11119 10706
rect 8756 10648 11058 10704
rect 11114 10648 11119 10704
rect 8756 10646 11119 10648
rect 7852 10644 7858 10646
rect 8569 10643 8635 10646
rect 11053 10643 11119 10646
rect 12390 10704 17099 10706
rect 12390 10648 17038 10704
rect 17094 10648 17099 10704
rect 12390 10646 17099 10648
rect 9765 10570 9831 10573
rect 5076 10568 9831 10570
rect 5076 10512 9770 10568
rect 9826 10512 9831 10568
rect 5076 10510 9831 10512
rect 9765 10507 9831 10510
rect 10041 10570 10107 10573
rect 12390 10570 12450 10646
rect 17033 10643 17099 10646
rect 18965 10706 19031 10709
rect 21081 10706 21147 10709
rect 18965 10704 21147 10706
rect 18965 10648 18970 10704
rect 19026 10648 21086 10704
rect 21142 10648 21147 10704
rect 18965 10646 21147 10648
rect 18965 10643 19031 10646
rect 21081 10643 21147 10646
rect 21449 10706 21515 10709
rect 22142 10706 22202 10752
rect 21449 10704 22202 10706
rect 21449 10648 21454 10704
rect 21510 10648 22202 10704
rect 21449 10646 22202 10648
rect 21449 10643 21515 10646
rect 16205 10570 16271 10573
rect 10041 10568 12450 10570
rect 10041 10512 10046 10568
rect 10102 10512 12450 10568
rect 10041 10510 12450 10512
rect 13724 10568 16271 10570
rect 13724 10512 16210 10568
rect 16266 10512 16271 10568
rect 13724 10510 16271 10512
rect 10041 10507 10107 10510
rect 0 10434 800 10464
rect 1945 10434 2011 10437
rect 0 10432 2011 10434
rect 0 10376 1950 10432
rect 2006 10376 2011 10432
rect 0 10374 2011 10376
rect 0 10344 800 10374
rect 1945 10371 2011 10374
rect 5574 10372 5580 10436
rect 5644 10434 5650 10436
rect 6453 10434 6519 10437
rect 7005 10436 7071 10437
rect 7005 10434 7052 10436
rect 5644 10432 6519 10434
rect 5644 10376 6458 10432
rect 6514 10376 6519 10432
rect 5644 10374 6519 10376
rect 6960 10432 7052 10434
rect 6960 10376 7010 10432
rect 6960 10374 7052 10376
rect 5644 10372 5650 10374
rect 6453 10371 6519 10374
rect 7005 10372 7052 10374
rect 7116 10372 7122 10436
rect 7189 10434 7255 10437
rect 9213 10434 9279 10437
rect 13261 10434 13327 10437
rect 7189 10432 8448 10434
rect 7189 10376 7194 10432
rect 7250 10376 8448 10432
rect 7189 10374 8448 10376
rect 7005 10371 7071 10372
rect 7189 10371 7255 10374
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 4797 10298 4863 10301
rect 6269 10298 6335 10301
rect 4797 10296 6335 10298
rect 4797 10240 4802 10296
rect 4858 10240 6274 10296
rect 6330 10240 6335 10296
rect 4797 10238 6335 10240
rect 4797 10235 4863 10238
rect 6269 10235 6335 10238
rect 6453 10298 6519 10301
rect 6913 10298 6979 10301
rect 6453 10296 6979 10298
rect 6453 10240 6458 10296
rect 6514 10240 6918 10296
rect 6974 10240 6979 10296
rect 6453 10238 6979 10240
rect 6453 10235 6519 10238
rect 6913 10235 6979 10238
rect 7373 10298 7439 10301
rect 7833 10300 7899 10301
rect 7782 10298 7788 10300
rect 7373 10296 7788 10298
rect 7852 10298 7899 10300
rect 7852 10296 7980 10298
rect 7373 10240 7378 10296
rect 7434 10240 7788 10296
rect 7894 10240 7980 10296
rect 7373 10238 7788 10240
rect 7373 10235 7439 10238
rect 7782 10236 7788 10238
rect 7852 10238 7980 10240
rect 7852 10236 7899 10238
rect 7833 10235 7899 10236
rect 3417 10162 3483 10165
rect 3236 10160 3483 10162
rect 3236 10104 3422 10160
rect 3478 10104 3483 10160
rect 3236 10102 3483 10104
rect 0 10026 800 10056
rect 1577 10026 1643 10029
rect 3236 10026 3296 10102
rect 3417 10099 3483 10102
rect 3601 10162 3667 10165
rect 4838 10162 4844 10164
rect 3601 10160 4844 10162
rect 3601 10104 3606 10160
rect 3662 10104 4844 10160
rect 3601 10102 4844 10104
rect 3601 10099 3667 10102
rect 4838 10100 4844 10102
rect 4908 10162 4914 10164
rect 7230 10162 7236 10164
rect 4908 10102 7236 10162
rect 4908 10100 4914 10102
rect 7230 10100 7236 10102
rect 7300 10100 7306 10164
rect 8388 10162 8448 10374
rect 9213 10432 13327 10434
rect 9213 10376 9218 10432
rect 9274 10376 13266 10432
rect 13322 10376 13327 10432
rect 9213 10374 13327 10376
rect 9213 10371 9279 10374
rect 13261 10371 13327 10374
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 9121 10298 9187 10301
rect 9121 10296 10288 10298
rect 9121 10240 9126 10296
rect 9182 10240 10288 10296
rect 9121 10238 10288 10240
rect 9121 10235 9187 10238
rect 9765 10162 9831 10165
rect 8388 10160 9831 10162
rect 8388 10104 9770 10160
rect 9826 10104 9831 10160
rect 8388 10102 9831 10104
rect 10228 10162 10288 10238
rect 10358 10236 10364 10300
rect 10428 10298 10434 10300
rect 13724 10298 13784 10510
rect 16205 10507 16271 10510
rect 17534 10508 17540 10572
rect 17604 10570 17610 10572
rect 17953 10570 18019 10573
rect 17604 10568 18019 10570
rect 17604 10512 17958 10568
rect 18014 10512 18019 10568
rect 17604 10510 18019 10512
rect 17604 10508 17610 10510
rect 17953 10507 18019 10510
rect 14457 10434 14523 10437
rect 16849 10434 16915 10437
rect 17534 10434 17540 10436
rect 14457 10432 17540 10434
rect 14457 10376 14462 10432
rect 14518 10376 16854 10432
rect 16910 10376 17540 10432
rect 14457 10374 17540 10376
rect 14457 10371 14523 10374
rect 16849 10371 16915 10374
rect 17534 10372 17540 10374
rect 17604 10372 17610 10436
rect 21173 10434 21239 10437
rect 22200 10434 23000 10464
rect 21173 10432 23000 10434
rect 21173 10376 21178 10432
rect 21234 10376 23000 10432
rect 21173 10374 23000 10376
rect 21173 10371 21239 10374
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 22200 10344 23000 10374
rect 19139 10303 19455 10304
rect 10428 10238 13784 10298
rect 15009 10298 15075 10301
rect 18822 10298 18828 10300
rect 15009 10296 18828 10298
rect 15009 10240 15014 10296
rect 15070 10240 18828 10296
rect 15009 10238 18828 10240
rect 10428 10236 10434 10238
rect 15009 10235 15075 10238
rect 18822 10236 18828 10238
rect 18892 10236 18898 10300
rect 15285 10162 15351 10165
rect 10228 10160 15351 10162
rect 10228 10104 15290 10160
rect 15346 10104 15351 10160
rect 10228 10102 15351 10104
rect 9765 10099 9831 10102
rect 15285 10099 15351 10102
rect 16021 10162 16087 10165
rect 20110 10162 20116 10164
rect 16021 10160 20116 10162
rect 16021 10104 16026 10160
rect 16082 10104 20116 10160
rect 16021 10102 20116 10104
rect 16021 10099 16087 10102
rect 20110 10100 20116 10102
rect 20180 10100 20186 10164
rect 0 10024 3296 10026
rect 0 9968 1582 10024
rect 1638 9968 3296 10024
rect 0 9966 3296 9968
rect 3417 10026 3483 10029
rect 5073 10026 5139 10029
rect 9213 10026 9279 10029
rect 10685 10026 10751 10029
rect 3417 10024 9279 10026
rect 3417 9968 3422 10024
rect 3478 9968 5078 10024
rect 5134 9968 9218 10024
rect 9274 9968 9279 10024
rect 3417 9966 9279 9968
rect 0 9936 800 9966
rect 1577 9963 1643 9966
rect 3417 9963 3483 9966
rect 5073 9963 5139 9966
rect 9213 9963 9279 9966
rect 9492 10024 10751 10026
rect 9492 9968 10690 10024
rect 10746 9968 10751 10024
rect 9492 9966 10751 9968
rect 5533 9892 5599 9893
rect 5533 9890 5580 9892
rect 5488 9888 5580 9890
rect 5488 9832 5538 9888
rect 5488 9830 5580 9832
rect 5533 9828 5580 9830
rect 5644 9828 5650 9892
rect 7046 9828 7052 9892
rect 7116 9890 7122 9892
rect 9029 9890 9095 9893
rect 7116 9888 9095 9890
rect 7116 9832 9034 9888
rect 9090 9832 9095 9888
rect 7116 9830 9095 9832
rect 7116 9828 7122 9830
rect 5533 9827 5599 9828
rect 9029 9827 9095 9830
rect 9254 9828 9260 9892
rect 9324 9890 9330 9892
rect 9492 9890 9552 9966
rect 10685 9963 10751 9966
rect 11094 9964 11100 10028
rect 11164 10026 11170 10028
rect 11513 10026 11579 10029
rect 11164 10024 11579 10026
rect 11164 9968 11518 10024
rect 11574 9968 11579 10024
rect 11164 9966 11579 9968
rect 11164 9964 11170 9966
rect 11513 9963 11579 9966
rect 15469 10026 15535 10029
rect 18689 10026 18755 10029
rect 15469 10024 18755 10026
rect 15469 9968 15474 10024
rect 15530 9968 18694 10024
rect 18750 9968 18755 10024
rect 15469 9966 18755 9968
rect 15469 9963 15535 9966
rect 18689 9963 18755 9966
rect 20621 10026 20687 10029
rect 22200 10026 23000 10056
rect 20621 10024 23000 10026
rect 20621 9968 20626 10024
rect 20682 9968 23000 10024
rect 20621 9966 23000 9968
rect 20621 9963 20687 9966
rect 22200 9936 23000 9966
rect 10041 9890 10107 9893
rect 9324 9830 9552 9890
rect 9630 9888 10107 9890
rect 9630 9832 10046 9888
rect 10102 9832 10107 9888
rect 9630 9830 10107 9832
rect 9324 9828 9330 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 6821 9754 6887 9757
rect 9630 9754 9690 9830
rect 10041 9827 10107 9830
rect 12566 9828 12572 9892
rect 12636 9890 12642 9892
rect 12893 9890 12959 9893
rect 12636 9888 12959 9890
rect 12636 9832 12898 9888
rect 12954 9832 12959 9888
rect 12636 9830 12959 9832
rect 12636 9828 12642 9830
rect 12893 9827 12959 9830
rect 18781 9890 18847 9893
rect 20529 9890 20595 9893
rect 18781 9888 20595 9890
rect 18781 9832 18786 9888
rect 18842 9832 20534 9888
rect 20590 9832 20595 9888
rect 18781 9830 20595 9832
rect 18781 9827 18847 9830
rect 20529 9827 20595 9830
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 6821 9752 9690 9754
rect 6821 9696 6826 9752
rect 6882 9696 9690 9752
rect 6821 9694 9690 9696
rect 10133 9756 10199 9757
rect 10133 9752 10180 9756
rect 10244 9754 10250 9756
rect 10133 9696 10138 9752
rect 6821 9691 6887 9694
rect 10133 9692 10180 9696
rect 10244 9694 10290 9754
rect 10244 9692 10250 9694
rect 12566 9692 12572 9756
rect 12636 9754 12642 9756
rect 16113 9754 16179 9757
rect 21265 9754 21331 9757
rect 12636 9752 16179 9754
rect 12636 9696 16118 9752
rect 16174 9696 16179 9752
rect 12636 9694 16179 9696
rect 12636 9692 12642 9694
rect 10133 9691 10199 9692
rect 16113 9691 16179 9694
rect 17910 9752 21331 9754
rect 17910 9696 21270 9752
rect 21326 9696 21331 9752
rect 17910 9694 21331 9696
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 2998 9556 3004 9620
rect 3068 9618 3074 9620
rect 4337 9618 4403 9621
rect 3068 9616 4403 9618
rect 3068 9560 4342 9616
rect 4398 9560 4403 9616
rect 3068 9558 4403 9560
rect 3068 9556 3074 9558
rect 4337 9555 4403 9558
rect 5206 9556 5212 9620
rect 5276 9618 5282 9620
rect 12617 9618 12683 9621
rect 5276 9584 7896 9618
rect 8112 9616 12683 9618
rect 8112 9584 12622 9616
rect 5276 9560 12622 9584
rect 12678 9560 12683 9616
rect 5276 9558 12683 9560
rect 5276 9556 5282 9558
rect 7836 9524 8172 9558
rect 12617 9555 12683 9558
rect 16205 9618 16271 9621
rect 17910 9618 17970 9694
rect 21265 9691 21331 9694
rect 16205 9616 17970 9618
rect 16205 9560 16210 9616
rect 16266 9560 17970 9616
rect 16205 9558 17970 9560
rect 18965 9618 19031 9621
rect 20161 9618 20227 9621
rect 22200 9618 23000 9648
rect 18965 9616 23000 9618
rect 18965 9560 18970 9616
rect 19026 9560 20166 9616
rect 20222 9560 23000 9616
rect 18965 9558 23000 9560
rect 16205 9555 16271 9558
rect 18965 9555 19031 9558
rect 20161 9555 20227 9558
rect 22200 9528 23000 9558
rect 1209 9482 1275 9485
rect 3233 9482 3299 9485
rect 1209 9480 3299 9482
rect 1209 9424 1214 9480
rect 1270 9424 3238 9480
rect 3294 9424 3299 9480
rect 1209 9422 3299 9424
rect 1209 9419 1275 9422
rect 3233 9419 3299 9422
rect 5901 9482 5967 9485
rect 6862 9482 6868 9484
rect 5901 9480 6868 9482
rect 5901 9424 5906 9480
rect 5962 9424 6868 9480
rect 5901 9422 6868 9424
rect 5901 9419 5967 9422
rect 6862 9420 6868 9422
rect 6932 9420 6938 9484
rect 13169 9482 13235 9485
rect 17769 9482 17835 9485
rect 8250 9480 13235 9482
rect 8250 9424 13174 9480
rect 13230 9424 13235 9480
rect 8250 9422 13235 9424
rect 4654 9284 4660 9348
rect 4724 9346 4730 9348
rect 8250 9346 8310 9422
rect 13169 9419 13235 9422
rect 13310 9480 17835 9482
rect 13310 9424 17774 9480
rect 17830 9424 17835 9480
rect 13310 9422 17835 9424
rect 4724 9286 8310 9346
rect 9857 9346 9923 9349
rect 9990 9346 9996 9348
rect 9857 9344 9996 9346
rect 9857 9288 9862 9344
rect 9918 9288 9996 9344
rect 9857 9286 9996 9288
rect 4724 9284 4730 9286
rect 9857 9283 9923 9286
rect 9990 9284 9996 9286
rect 10060 9284 10066 9348
rect 11789 9346 11855 9349
rect 13310 9346 13370 9422
rect 17769 9419 17835 9422
rect 19425 9482 19491 9485
rect 19425 9480 20316 9482
rect 19425 9424 19430 9480
rect 19486 9424 20316 9480
rect 19425 9422 20316 9424
rect 19425 9419 19491 9422
rect 20256 9349 20316 9422
rect 11789 9344 13370 9346
rect 11789 9288 11794 9344
rect 11850 9288 13370 9344
rect 11789 9286 13370 9288
rect 11789 9283 11855 9286
rect 14774 9284 14780 9348
rect 14844 9346 14850 9348
rect 17350 9346 17356 9348
rect 14844 9286 17356 9346
rect 14844 9284 14850 9286
rect 17350 9284 17356 9286
rect 17420 9284 17426 9348
rect 20253 9344 20319 9349
rect 20253 9288 20258 9344
rect 20314 9288 20319 9344
rect 20253 9283 20319 9288
rect 3545 9280 3861 9281
rect 0 9210 800 9240
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 1393 9210 1459 9213
rect 8293 9210 8359 9213
rect 0 9208 3296 9210
rect 0 9152 1398 9208
rect 1454 9152 3296 9208
rect 0 9150 3296 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 3236 9074 3296 9150
rect 3926 9208 8359 9210
rect 3926 9152 8298 9208
rect 8354 9152 8359 9208
rect 3926 9150 8359 9152
rect 3926 9074 3986 9150
rect 8293 9147 8359 9150
rect 9438 9148 9444 9212
rect 9508 9210 9514 9212
rect 9581 9210 9647 9213
rect 13813 9210 13879 9213
rect 9508 9208 9647 9210
rect 9508 9152 9586 9208
rect 9642 9152 9647 9208
rect 9508 9150 9647 9152
rect 9508 9148 9514 9150
rect 9581 9147 9647 9150
rect 9814 9208 13879 9210
rect 9814 9152 13818 9208
rect 13874 9152 13879 9208
rect 9814 9150 13879 9152
rect 3236 9014 3986 9074
rect 5206 9012 5212 9076
rect 5276 9074 5282 9076
rect 5533 9074 5599 9077
rect 5276 9072 5599 9074
rect 5276 9016 5538 9072
rect 5594 9016 5599 9072
rect 5276 9014 5599 9016
rect 5276 9012 5282 9014
rect 5533 9011 5599 9014
rect 6085 9074 6151 9077
rect 9814 9076 9874 9150
rect 13813 9147 13879 9150
rect 16757 9210 16823 9213
rect 18045 9210 18111 9213
rect 18321 9210 18387 9213
rect 16757 9208 18387 9210
rect 16757 9152 16762 9208
rect 16818 9152 18050 9208
rect 18106 9152 18326 9208
rect 18382 9152 18387 9208
rect 16757 9150 18387 9152
rect 16757 9147 16823 9150
rect 18045 9147 18111 9150
rect 18321 9147 18387 9150
rect 22001 9210 22067 9213
rect 22200 9210 23000 9240
rect 22001 9208 23000 9210
rect 22001 9152 22006 9208
rect 22062 9152 23000 9208
rect 22001 9150 23000 9152
rect 22001 9147 22067 9150
rect 22200 9120 23000 9150
rect 9806 9074 9812 9076
rect 6085 9072 9812 9074
rect 6085 9016 6090 9072
rect 6146 9016 9812 9072
rect 6085 9014 9812 9016
rect 6085 9011 6151 9014
rect 9806 9012 9812 9014
rect 9876 9012 9882 9076
rect 10133 9074 10199 9077
rect 16665 9074 16731 9077
rect 10133 9072 16731 9074
rect 10133 9016 10138 9072
rect 10194 9016 16670 9072
rect 16726 9016 16731 9072
rect 10133 9014 16731 9016
rect 10133 9011 10199 9014
rect 16665 9011 16731 9014
rect 16982 9012 16988 9076
rect 17052 9074 17058 9076
rect 17861 9074 17927 9077
rect 20713 9074 20779 9077
rect 17052 9072 20779 9074
rect 17052 9016 17866 9072
rect 17922 9016 20718 9072
rect 20774 9016 20779 9072
rect 17052 9014 20779 9016
rect 17052 9012 17058 9014
rect 17861 9011 17927 9014
rect 20713 9011 20779 9014
rect 2865 8938 2931 8941
rect 5022 8938 5028 8940
rect 2865 8936 5028 8938
rect 2865 8880 2870 8936
rect 2926 8880 5028 8936
rect 2865 8878 5028 8880
rect 2865 8875 2931 8878
rect 5022 8876 5028 8878
rect 5092 8938 5098 8940
rect 5257 8938 5323 8941
rect 8293 8938 8359 8941
rect 13721 8938 13787 8941
rect 21081 8938 21147 8941
rect 5092 8936 8359 8938
rect 5092 8880 5262 8936
rect 5318 8880 8298 8936
rect 8354 8880 8359 8936
rect 5092 8878 8359 8880
rect 5092 8876 5098 8878
rect 5257 8875 5323 8878
rect 8293 8875 8359 8878
rect 9262 8936 13787 8938
rect 9262 8880 13726 8936
rect 13782 8880 13787 8936
rect 9262 8878 13787 8880
rect 0 8802 800 8832
rect 3049 8802 3115 8805
rect 0 8800 3115 8802
rect 0 8744 3054 8800
rect 3110 8744 3115 8800
rect 0 8742 3115 8744
rect 0 8712 800 8742
rect 3049 8739 3115 8742
rect 4889 8800 4955 8805
rect 4889 8744 4894 8800
rect 4950 8744 4955 8800
rect 4889 8739 4955 8744
rect 5257 8802 5323 8805
rect 5942 8802 5948 8804
rect 5257 8800 5948 8802
rect 5257 8744 5262 8800
rect 5318 8744 5948 8800
rect 5257 8742 5948 8744
rect 5257 8739 5323 8742
rect 5942 8740 5948 8742
rect 6012 8740 6018 8804
rect 6678 8740 6684 8804
rect 6748 8802 6754 8804
rect 7833 8802 7899 8805
rect 9121 8802 9187 8805
rect 6748 8800 7899 8802
rect 6748 8744 7838 8800
rect 7894 8744 7899 8800
rect 6748 8742 7899 8744
rect 6748 8740 6754 8742
rect 7833 8739 7899 8742
rect 7974 8800 9187 8802
rect 7974 8744 9126 8800
rect 9182 8744 9187 8800
rect 7974 8742 9187 8744
rect 1577 8666 1643 8669
rect 2497 8668 2563 8669
rect 1894 8666 1900 8668
rect 1577 8664 1900 8666
rect 1577 8608 1582 8664
rect 1638 8608 1900 8664
rect 1577 8606 1900 8608
rect 1577 8603 1643 8606
rect 1894 8604 1900 8606
rect 1964 8604 1970 8668
rect 2446 8604 2452 8668
rect 2516 8666 2563 8668
rect 4892 8666 4952 8739
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 6545 8666 6611 8669
rect 7974 8666 8034 8742
rect 9121 8739 9187 8742
rect 8150 8666 8156 8668
rect 2516 8664 2608 8666
rect 2558 8608 2608 8664
rect 2516 8606 2608 8608
rect 4892 8606 6010 8666
rect 2516 8604 2563 8606
rect 2497 8603 2563 8604
rect 1710 8468 1716 8532
rect 1780 8530 1786 8532
rect 2865 8530 2931 8533
rect 5533 8530 5599 8533
rect 1780 8470 2790 8530
rect 1780 8468 1786 8470
rect 0 8394 800 8424
rect 1209 8394 1275 8397
rect 0 8392 1275 8394
rect 0 8336 1214 8392
rect 1270 8336 1275 8392
rect 0 8334 1275 8336
rect 2730 8394 2790 8470
rect 2865 8528 5599 8530
rect 2865 8472 2870 8528
rect 2926 8472 5538 8528
rect 5594 8472 5599 8528
rect 2865 8470 5599 8472
rect 5950 8530 6010 8606
rect 6545 8664 8034 8666
rect 6545 8608 6550 8664
rect 6606 8608 8034 8664
rect 6545 8606 8034 8608
rect 6545 8603 6611 8606
rect 8112 8604 8156 8666
rect 8220 8604 8226 8668
rect 8293 8666 8359 8669
rect 9262 8666 9322 8878
rect 13721 8875 13787 8878
rect 13862 8936 21147 8938
rect 13862 8880 21086 8936
rect 21142 8880 21147 8936
rect 13862 8878 21147 8880
rect 12985 8802 13051 8805
rect 13629 8802 13695 8805
rect 13862 8802 13922 8878
rect 21081 8875 21147 8878
rect 21265 8938 21331 8941
rect 21265 8936 22202 8938
rect 21265 8880 21270 8936
rect 21326 8880 22202 8936
rect 21265 8878 22202 8880
rect 21265 8875 21331 8878
rect 12985 8800 13922 8802
rect 12985 8744 12990 8800
rect 13046 8744 13634 8800
rect 13690 8744 13922 8800
rect 12985 8742 13922 8744
rect 22142 8832 22202 8878
rect 22142 8742 23000 8832
rect 12985 8739 13051 8742
rect 13629 8739 13695 8742
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 22200 8712 23000 8742
rect 21738 8671 22054 8672
rect 8293 8664 9322 8666
rect 8293 8608 8298 8664
rect 8354 8608 9322 8664
rect 8293 8606 9322 8608
rect 9397 8666 9463 8669
rect 10869 8666 10935 8669
rect 9397 8664 10935 8666
rect 9397 8608 9402 8664
rect 9458 8608 10874 8664
rect 10930 8608 10935 8664
rect 9397 8606 10935 8608
rect 8112 8533 8172 8604
rect 8293 8603 8359 8606
rect 9397 8603 9463 8606
rect 10869 8603 10935 8606
rect 12065 8666 12131 8669
rect 13997 8666 14063 8669
rect 12065 8664 14063 8666
rect 12065 8608 12070 8664
rect 12126 8608 14002 8664
rect 14058 8608 14063 8664
rect 12065 8606 14063 8608
rect 12065 8603 12131 8606
rect 13997 8603 14063 8606
rect 17953 8666 18019 8669
rect 19149 8666 19215 8669
rect 17953 8664 19215 8666
rect 17953 8608 17958 8664
rect 18014 8608 19154 8664
rect 19210 8608 19215 8664
rect 17953 8606 19215 8608
rect 17953 8603 18019 8606
rect 19149 8603 19215 8606
rect 7097 8530 7163 8533
rect 7465 8532 7531 8533
rect 5950 8528 7163 8530
rect 5950 8472 7102 8528
rect 7158 8472 7163 8528
rect 5950 8470 7163 8472
rect 2865 8467 2931 8470
rect 5533 8467 5599 8470
rect 7097 8467 7163 8470
rect 7414 8468 7420 8532
rect 7484 8530 7531 8532
rect 7484 8528 7576 8530
rect 7526 8472 7576 8528
rect 7484 8470 7576 8472
rect 8109 8528 8175 8533
rect 8109 8472 8114 8528
rect 8170 8472 8175 8528
rect 7484 8468 7531 8470
rect 7465 8467 7531 8468
rect 8109 8467 8175 8472
rect 11329 8530 11395 8533
rect 21725 8530 21791 8533
rect 11329 8528 21791 8530
rect 11329 8472 11334 8528
rect 11390 8472 21730 8528
rect 21786 8472 21791 8528
rect 11329 8470 21791 8472
rect 11329 8467 11395 8470
rect 21725 8467 21791 8470
rect 8250 8394 8770 8428
rect 9857 8394 9923 8397
rect 2730 8392 9923 8394
rect 2730 8368 9862 8392
rect 2730 8334 8310 8368
rect 8710 8336 9862 8368
rect 9918 8336 9923 8392
rect 8710 8334 9923 8336
rect 0 8304 800 8334
rect 1209 8331 1275 8334
rect 9857 8331 9923 8334
rect 13077 8394 13143 8397
rect 17902 8394 17908 8396
rect 13077 8392 17908 8394
rect 13077 8336 13082 8392
rect 13138 8336 17908 8392
rect 13077 8334 17908 8336
rect 13077 8331 13143 8334
rect 17902 8332 17908 8334
rect 17972 8332 17978 8396
rect 19333 8394 19399 8397
rect 19014 8392 19399 8394
rect 19014 8336 19338 8392
rect 19394 8336 19399 8392
rect 19014 8334 19399 8336
rect 1393 8258 1459 8261
rect 3969 8258 4035 8261
rect 8569 8258 8635 8261
rect 1393 8256 2790 8258
rect 1393 8200 1398 8256
rect 1454 8200 2790 8256
rect 1393 8198 2790 8200
rect 1393 8195 1459 8198
rect 0 7986 800 8016
rect 933 7986 999 7989
rect 0 7984 999 7986
rect 0 7928 938 7984
rect 994 7928 999 7984
rect 0 7926 999 7928
rect 2730 7986 2790 8198
rect 3969 8256 8635 8258
rect 3969 8200 3974 8256
rect 4030 8200 8574 8256
rect 8630 8200 8635 8256
rect 3969 8198 8635 8200
rect 3969 8195 4035 8198
rect 8569 8195 8635 8198
rect 15837 8258 15903 8261
rect 19014 8258 19074 8334
rect 19333 8331 19399 8334
rect 20345 8394 20411 8397
rect 22200 8394 23000 8424
rect 20345 8392 23000 8394
rect 20345 8336 20350 8392
rect 20406 8336 23000 8392
rect 20345 8334 23000 8336
rect 20345 8331 20411 8334
rect 22200 8304 23000 8334
rect 15837 8256 19074 8258
rect 15837 8200 15842 8256
rect 15898 8200 19074 8256
rect 15837 8198 19074 8200
rect 15837 8195 15903 8198
rect 19926 8196 19932 8260
rect 19996 8258 20002 8260
rect 20253 8258 20319 8261
rect 19996 8256 20319 8258
rect 19996 8200 20258 8256
rect 20314 8200 20319 8256
rect 19996 8198 20319 8200
rect 19996 8196 20002 8198
rect 20253 8195 20319 8198
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 5390 8060 5396 8124
rect 5460 8122 5466 8124
rect 6085 8122 6151 8125
rect 5460 8120 6151 8122
rect 5460 8064 6090 8120
rect 6146 8064 6151 8120
rect 5460 8062 6151 8064
rect 5460 8060 5466 8062
rect 6085 8059 6151 8062
rect 7833 8122 7899 8125
rect 8569 8122 8635 8125
rect 7833 8120 8635 8122
rect 7833 8064 7838 8120
rect 7894 8064 8574 8120
rect 8630 8064 8635 8120
rect 7833 8062 8635 8064
rect 7833 8059 7899 8062
rect 8569 8059 8635 8062
rect 15377 8122 15443 8125
rect 15929 8122 15995 8125
rect 18781 8122 18847 8125
rect 15377 8120 18847 8122
rect 15377 8064 15382 8120
rect 15438 8064 15934 8120
rect 15990 8064 18786 8120
rect 18842 8064 18847 8120
rect 15377 8062 18847 8064
rect 15377 8059 15443 8062
rect 15929 8059 15995 8062
rect 18781 8059 18847 8062
rect 9305 7986 9371 7989
rect 2730 7984 9371 7986
rect 2730 7928 9310 7984
rect 9366 7928 9371 7984
rect 2730 7926 9371 7928
rect 0 7896 800 7926
rect 933 7923 999 7926
rect 9305 7923 9371 7926
rect 10358 7924 10364 7988
rect 10428 7986 10434 7988
rect 11237 7986 11303 7989
rect 10428 7984 11303 7986
rect 10428 7928 11242 7984
rect 11298 7928 11303 7984
rect 10428 7926 11303 7928
rect 10428 7924 10434 7926
rect 11237 7923 11303 7926
rect 13077 7986 13143 7989
rect 15326 7986 15332 7988
rect 13077 7984 15332 7986
rect 13077 7928 13082 7984
rect 13138 7928 15332 7984
rect 13077 7926 15332 7928
rect 13077 7923 13143 7926
rect 15326 7924 15332 7926
rect 15396 7924 15402 7988
rect 17769 7986 17835 7989
rect 16990 7984 17835 7986
rect 16990 7928 17774 7984
rect 17830 7928 17835 7984
rect 16990 7926 17835 7928
rect 1577 7850 1643 7853
rect 4102 7850 4108 7852
rect 1577 7848 4108 7850
rect 1577 7792 1582 7848
rect 1638 7792 4108 7848
rect 1577 7790 4108 7792
rect 1577 7787 1643 7790
rect 4102 7788 4108 7790
rect 4172 7788 4178 7852
rect 5073 7850 5139 7853
rect 5206 7850 5212 7852
rect 5073 7848 5212 7850
rect 5073 7792 5078 7848
rect 5134 7792 5212 7848
rect 5073 7790 5212 7792
rect 5073 7787 5139 7790
rect 5206 7788 5212 7790
rect 5276 7788 5282 7852
rect 5809 7850 5875 7853
rect 5942 7850 5948 7852
rect 5809 7848 5948 7850
rect 5809 7792 5814 7848
rect 5870 7792 5948 7848
rect 5809 7790 5948 7792
rect 5809 7787 5875 7790
rect 5942 7788 5948 7790
rect 6012 7850 6018 7852
rect 11697 7850 11763 7853
rect 6012 7848 11763 7850
rect 6012 7792 11702 7848
rect 11758 7792 11763 7848
rect 6012 7790 11763 7792
rect 6012 7788 6018 7790
rect 11697 7787 11763 7790
rect 12617 7850 12683 7853
rect 13353 7850 13419 7853
rect 16990 7850 17050 7926
rect 17769 7923 17835 7926
rect 17953 7986 18019 7989
rect 19885 7986 19951 7989
rect 22200 7986 23000 8016
rect 17953 7984 23000 7986
rect 17953 7928 17958 7984
rect 18014 7928 19890 7984
rect 19946 7928 23000 7984
rect 17953 7926 23000 7928
rect 17953 7923 18019 7926
rect 19885 7923 19951 7926
rect 22200 7896 23000 7926
rect 12617 7848 17050 7850
rect 12617 7792 12622 7848
rect 12678 7792 13358 7848
rect 13414 7792 17050 7848
rect 12617 7790 17050 7792
rect 12617 7787 12683 7790
rect 13353 7787 13419 7790
rect 2589 7714 2655 7717
rect 4286 7714 4292 7716
rect 2589 7712 4292 7714
rect 2589 7656 2594 7712
rect 2650 7656 4292 7712
rect 2589 7654 4292 7656
rect 2589 7651 2655 7654
rect 4286 7652 4292 7654
rect 4356 7652 4362 7716
rect 4797 7714 4863 7717
rect 5022 7714 5028 7716
rect 4797 7712 5028 7714
rect 4797 7656 4802 7712
rect 4858 7656 5028 7712
rect 4797 7654 5028 7656
rect 4797 7651 4863 7654
rect 5022 7652 5028 7654
rect 5092 7652 5098 7716
rect 7230 7652 7236 7716
rect 7300 7714 7306 7716
rect 7373 7714 7439 7717
rect 7300 7712 7439 7714
rect 7300 7656 7378 7712
rect 7434 7656 7439 7712
rect 7300 7654 7439 7656
rect 7300 7652 7306 7654
rect 7373 7651 7439 7654
rect 7741 7714 7807 7717
rect 10542 7714 10548 7716
rect 7741 7712 10548 7714
rect 7741 7656 7746 7712
rect 7802 7656 10548 7712
rect 7741 7654 10548 7656
rect 7741 7651 7807 7654
rect 10542 7652 10548 7654
rect 10612 7652 10618 7716
rect 6144 7648 6460 7649
rect 0 7578 800 7608
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 2865 7578 2931 7581
rect 0 7576 2931 7578
rect 0 7520 2870 7576
rect 2926 7520 2931 7576
rect 0 7518 2931 7520
rect 0 7488 800 7518
rect 2865 7515 2931 7518
rect 3141 7578 3207 7581
rect 5574 7578 5580 7580
rect 3141 7576 5580 7578
rect 3141 7520 3146 7576
rect 3202 7520 5580 7576
rect 3141 7518 5580 7520
rect 3141 7515 3207 7518
rect 5574 7516 5580 7518
rect 5644 7516 5650 7580
rect 7376 7578 7436 7651
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 11053 7578 11119 7581
rect 7376 7576 11119 7578
rect 7376 7520 11058 7576
rect 11114 7520 11119 7576
rect 7376 7518 11119 7520
rect 11053 7515 11119 7518
rect 11789 7578 11855 7581
rect 12893 7578 12959 7581
rect 15377 7578 15443 7581
rect 11789 7576 12959 7578
rect 11789 7520 11794 7576
rect 11850 7520 12898 7576
rect 12954 7520 12959 7576
rect 11789 7518 12959 7520
rect 11789 7515 11855 7518
rect 12893 7515 12959 7518
rect 13310 7576 15443 7578
rect 13310 7520 15382 7576
rect 15438 7520 15443 7576
rect 13310 7518 15443 7520
rect 16990 7578 17050 7790
rect 17769 7850 17835 7853
rect 19609 7850 19675 7853
rect 17769 7848 19675 7850
rect 17769 7792 17774 7848
rect 17830 7792 19614 7848
rect 19670 7792 19675 7848
rect 17769 7790 19675 7792
rect 17769 7787 17835 7790
rect 19609 7787 19675 7790
rect 20437 7850 20503 7853
rect 20437 7848 22018 7850
rect 20437 7792 20442 7848
rect 20498 7816 22018 7848
rect 20498 7792 22202 7816
rect 20437 7790 22202 7792
rect 20437 7787 20503 7790
rect 21958 7756 22202 7790
rect 17401 7714 17467 7717
rect 17953 7714 18019 7717
rect 17401 7712 18019 7714
rect 17401 7656 17406 7712
rect 17462 7656 17958 7712
rect 18014 7656 18019 7712
rect 17401 7654 18019 7656
rect 17401 7651 17467 7654
rect 17953 7651 18019 7654
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 22142 7608 22202 7756
rect 16990 7518 17786 7578
rect 22142 7518 23000 7608
rect 3693 7442 3759 7445
rect 10501 7442 10567 7445
rect 3693 7440 10567 7442
rect 3693 7384 3698 7440
rect 3754 7384 10506 7440
rect 10562 7384 10567 7440
rect 3693 7382 10567 7384
rect 3693 7379 3759 7382
rect 10501 7379 10567 7382
rect 11697 7442 11763 7445
rect 13310 7442 13370 7518
rect 15377 7515 15443 7518
rect 14549 7442 14615 7445
rect 11697 7440 13370 7442
rect 11697 7384 11702 7440
rect 11758 7384 13370 7440
rect 11697 7382 13370 7384
rect 13494 7440 14615 7442
rect 13494 7384 14554 7440
rect 14610 7384 14615 7440
rect 13494 7382 14615 7384
rect 11697 7379 11763 7382
rect 1669 7306 1735 7309
rect 13494 7306 13554 7382
rect 14549 7379 14615 7382
rect 15193 7442 15259 7445
rect 17534 7442 17540 7444
rect 15193 7440 17540 7442
rect 15193 7384 15198 7440
rect 15254 7384 17540 7440
rect 15193 7382 17540 7384
rect 15193 7379 15259 7382
rect 17534 7380 17540 7382
rect 17604 7380 17610 7444
rect 17726 7442 17786 7518
rect 22200 7488 23000 7518
rect 21909 7442 21975 7445
rect 17726 7440 21975 7442
rect 17726 7384 21914 7440
rect 21970 7384 21975 7440
rect 17726 7382 21975 7384
rect 21909 7379 21975 7382
rect 20989 7306 21055 7309
rect 1669 7304 13554 7306
rect 1669 7248 1674 7304
rect 1730 7248 13554 7304
rect 1669 7246 13554 7248
rect 13724 7304 21055 7306
rect 13724 7248 20994 7304
rect 21050 7248 21055 7304
rect 13724 7246 21055 7248
rect 1669 7243 1735 7246
rect 0 7170 800 7200
rect 1393 7170 1459 7173
rect 0 7168 1459 7170
rect 0 7112 1398 7168
rect 1454 7112 1459 7168
rect 0 7110 1459 7112
rect 0 7080 800 7110
rect 1393 7107 1459 7110
rect 3969 7170 4035 7173
rect 7373 7172 7439 7173
rect 10041 7172 10107 7173
rect 6678 7170 6684 7172
rect 3969 7168 6684 7170
rect 3969 7112 3974 7168
rect 4030 7112 6684 7168
rect 3969 7110 6684 7112
rect 3969 7107 4035 7110
rect 6678 7108 6684 7110
rect 6748 7108 6754 7172
rect 7373 7170 7420 7172
rect 7328 7168 7420 7170
rect 7328 7112 7378 7168
rect 7328 7110 7420 7112
rect 7373 7108 7420 7110
rect 7484 7108 7490 7172
rect 9990 7170 9996 7172
rect 9950 7110 9996 7170
rect 10060 7168 10107 7172
rect 10102 7112 10107 7168
rect 9990 7108 9996 7110
rect 10060 7108 10107 7112
rect 7373 7107 7439 7108
rect 10041 7107 10107 7108
rect 10225 7170 10291 7173
rect 13724 7170 13784 7246
rect 20989 7243 21055 7246
rect 10225 7168 13784 7170
rect 10225 7112 10230 7168
rect 10286 7112 13784 7168
rect 10225 7110 13784 7112
rect 10225 7107 10291 7110
rect 17166 7108 17172 7172
rect 17236 7170 17242 7172
rect 17401 7170 17467 7173
rect 17236 7168 17467 7170
rect 17236 7112 17406 7168
rect 17462 7112 17467 7168
rect 17236 7110 17467 7112
rect 17236 7108 17242 7110
rect 17401 7107 17467 7110
rect 19609 7170 19675 7173
rect 22200 7170 23000 7200
rect 19609 7168 23000 7170
rect 19609 7112 19614 7168
rect 19670 7112 23000 7168
rect 19609 7110 23000 7112
rect 19609 7107 19675 7110
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 22200 7080 23000 7110
rect 19139 7039 19455 7040
rect 4337 7034 4403 7037
rect 4838 7034 4844 7036
rect 4337 7032 4844 7034
rect 4337 6976 4342 7032
rect 4398 6976 4844 7032
rect 4337 6974 4844 6976
rect 4337 6971 4403 6974
rect 4838 6972 4844 6974
rect 4908 6972 4914 7036
rect 8109 7034 8175 7037
rect 8518 7034 8524 7036
rect 8109 7032 8524 7034
rect 8109 6976 8114 7032
rect 8170 6976 8524 7032
rect 8109 6974 8524 6976
rect 8109 6971 8175 6974
rect 8518 6972 8524 6974
rect 8588 6972 8594 7036
rect 9305 7034 9371 7037
rect 9438 7034 9444 7036
rect 9305 7032 9444 7034
rect 9305 6976 9310 7032
rect 9366 6976 9444 7032
rect 9305 6974 9444 6976
rect 9305 6971 9371 6974
rect 9438 6972 9444 6974
rect 9508 7034 9514 7036
rect 11697 7034 11763 7037
rect 9508 7032 11763 7034
rect 9508 6976 11702 7032
rect 11758 6976 11763 7032
rect 9508 6974 11763 6976
rect 9508 6972 9514 6974
rect 11697 6971 11763 6974
rect 12525 7034 12591 7037
rect 13445 7034 13511 7037
rect 12525 7032 13511 7034
rect 12525 6976 12530 7032
rect 12586 6976 13450 7032
rect 13506 6976 13511 7032
rect 12525 6974 13511 6976
rect 12525 6971 12591 6974
rect 13445 6971 13511 6974
rect 13721 7032 13787 7037
rect 20161 7034 20227 7037
rect 13721 6976 13726 7032
rect 13782 6976 13787 7032
rect 13721 6971 13787 6976
rect 14414 6974 19074 7034
rect 1577 6898 1643 6901
rect 1710 6898 1716 6900
rect 1577 6896 1716 6898
rect 1577 6840 1582 6896
rect 1638 6840 1716 6896
rect 1577 6838 1716 6840
rect 1577 6835 1643 6838
rect 1710 6836 1716 6838
rect 1780 6836 1786 6900
rect 2037 6898 2103 6901
rect 3325 6898 3391 6901
rect 2037 6896 3391 6898
rect 2037 6840 2042 6896
rect 2098 6840 3330 6896
rect 3386 6840 3391 6896
rect 2037 6838 3391 6840
rect 2037 6835 2103 6838
rect 3325 6835 3391 6838
rect 3509 6898 3575 6901
rect 3918 6898 3924 6900
rect 3509 6896 3924 6898
rect 3509 6840 3514 6896
rect 3570 6840 3924 6896
rect 3509 6838 3924 6840
rect 3509 6835 3575 6838
rect 3918 6836 3924 6838
rect 3988 6836 3994 6900
rect 4245 6898 4311 6901
rect 7741 6898 7807 6901
rect 4245 6896 7807 6898
rect 4245 6840 4250 6896
rect 4306 6840 7746 6896
rect 7802 6840 7807 6896
rect 4245 6838 7807 6840
rect 4245 6835 4311 6838
rect 7741 6835 7807 6838
rect 8017 6898 8083 6901
rect 13261 6898 13327 6901
rect 8017 6896 13327 6898
rect 8017 6840 8022 6896
rect 8078 6840 13266 6896
rect 13322 6840 13327 6896
rect 8017 6838 13327 6840
rect 13724 6898 13784 6971
rect 14414 6898 14474 6974
rect 13724 6838 14474 6898
rect 15193 6898 15259 6901
rect 15878 6898 15884 6900
rect 15193 6896 15884 6898
rect 15193 6840 15198 6896
rect 15254 6840 15884 6896
rect 15193 6838 15884 6840
rect 8017 6835 8083 6838
rect 13261 6835 13327 6838
rect 15193 6835 15259 6838
rect 15878 6836 15884 6838
rect 15948 6836 15954 6900
rect 17677 6898 17743 6901
rect 18638 6898 18644 6900
rect 17677 6896 18644 6898
rect 17677 6840 17682 6896
rect 17738 6840 18644 6896
rect 17677 6838 18644 6840
rect 17677 6835 17743 6838
rect 18638 6836 18644 6838
rect 18708 6898 18714 6900
rect 18873 6898 18939 6901
rect 18708 6896 18939 6898
rect 18708 6840 18878 6896
rect 18934 6840 18939 6896
rect 18708 6838 18939 6840
rect 19014 6898 19074 6974
rect 19566 7032 20227 7034
rect 19566 6976 20166 7032
rect 20222 6976 20227 7032
rect 19566 6974 20227 6976
rect 19566 6898 19626 6974
rect 20161 6971 20227 6974
rect 19014 6838 19626 6898
rect 18708 6836 18714 6838
rect 18873 6835 18939 6838
rect 0 6762 800 6792
rect 933 6762 999 6765
rect 4981 6762 5047 6765
rect 13261 6762 13327 6765
rect 21357 6762 21423 6765
rect 0 6760 999 6762
rect 0 6704 938 6760
rect 994 6704 999 6760
rect 0 6702 999 6704
rect 0 6672 800 6702
rect 933 6699 999 6702
rect 2730 6760 8402 6762
rect 2730 6704 4986 6760
rect 5042 6704 8402 6760
rect 2730 6702 8402 6704
rect 2730 6629 2790 6702
rect 4981 6699 5047 6702
rect 2681 6628 2790 6629
rect 4705 6628 4771 6629
rect 2630 6626 2636 6628
rect 2554 6566 2636 6626
rect 2700 6624 2790 6628
rect 2742 6568 2790 6624
rect 2630 6564 2636 6566
rect 2700 6566 2790 6568
rect 2700 6564 2747 6566
rect 4654 6564 4660 6628
rect 4724 6626 4771 6628
rect 4981 6626 5047 6629
rect 5717 6626 5783 6629
rect 4724 6624 4816 6626
rect 4766 6568 4816 6624
rect 4724 6566 4816 6568
rect 4981 6624 5783 6626
rect 4981 6568 4986 6624
rect 5042 6568 5722 6624
rect 5778 6568 5783 6624
rect 4981 6566 5783 6568
rect 8342 6626 8402 6702
rect 11148 6760 21423 6762
rect 11148 6704 13266 6760
rect 13322 6704 21362 6760
rect 21418 6704 21423 6760
rect 11148 6702 21423 6704
rect 9305 6626 9371 6629
rect 8342 6624 9371 6626
rect 8342 6568 9310 6624
rect 9366 6568 9371 6624
rect 8342 6566 9371 6568
rect 4724 6564 4771 6566
rect 2681 6563 2747 6564
rect 4705 6563 4771 6564
rect 4981 6563 5047 6566
rect 5717 6563 5783 6566
rect 9305 6563 9371 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 2037 6490 2103 6493
rect 2262 6490 2268 6492
rect 2037 6488 2268 6490
rect 2037 6432 2042 6488
rect 2098 6432 2268 6488
rect 2037 6430 2268 6432
rect 2037 6427 2103 6430
rect 2262 6428 2268 6430
rect 2332 6490 2338 6492
rect 7649 6490 7715 6493
rect 9765 6490 9831 6493
rect 11148 6490 11208 6702
rect 13261 6699 13327 6702
rect 21357 6699 21423 6702
rect 22001 6762 22067 6765
rect 22200 6762 23000 6792
rect 22001 6760 23000 6762
rect 22001 6704 22006 6760
rect 22062 6704 23000 6760
rect 22001 6702 23000 6704
rect 22001 6699 22067 6702
rect 22200 6672 23000 6702
rect 17309 6626 17375 6629
rect 18505 6626 18571 6629
rect 19241 6626 19307 6629
rect 17309 6624 19307 6626
rect 17309 6568 17314 6624
rect 17370 6568 18510 6624
rect 18566 6568 19246 6624
rect 19302 6568 19307 6624
rect 17309 6566 19307 6568
rect 17309 6563 17375 6566
rect 18505 6563 18571 6566
rect 19241 6563 19307 6566
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 17677 6490 17743 6493
rect 2332 6430 6010 6490
rect 2332 6428 2338 6430
rect 0 6354 800 6384
rect 3509 6354 3575 6357
rect 0 6352 3575 6354
rect 0 6296 3514 6352
rect 3570 6296 3575 6352
rect 0 6294 3575 6296
rect 0 6264 800 6294
rect 3509 6291 3575 6294
rect 4102 6292 4108 6356
rect 4172 6354 4178 6356
rect 5257 6354 5323 6357
rect 4172 6352 5323 6354
rect 4172 6296 5262 6352
rect 5318 6296 5323 6352
rect 4172 6294 5323 6296
rect 5950 6354 6010 6430
rect 7649 6488 9831 6490
rect 7649 6432 7654 6488
rect 7710 6432 9770 6488
rect 9826 6432 9831 6488
rect 7649 6430 9831 6432
rect 7649 6427 7715 6430
rect 9765 6427 9831 6430
rect 10550 6430 11208 6490
rect 16944 6488 17743 6490
rect 16944 6432 17682 6488
rect 17738 6432 17743 6488
rect 16944 6430 17743 6432
rect 6361 6354 6427 6357
rect 5950 6352 6427 6354
rect 5950 6296 6366 6352
rect 6422 6296 6427 6352
rect 5950 6294 6427 6296
rect 4172 6292 4178 6294
rect 5257 6291 5323 6294
rect 6361 6291 6427 6294
rect 6545 6354 6611 6357
rect 6821 6354 6887 6357
rect 6545 6352 6887 6354
rect 6545 6296 6550 6352
rect 6606 6296 6826 6352
rect 6882 6296 6887 6352
rect 6545 6294 6887 6296
rect 6545 6291 6611 6294
rect 6821 6291 6887 6294
rect 7925 6354 7991 6357
rect 8477 6354 8543 6357
rect 10550 6354 10610 6430
rect 10961 6354 11027 6357
rect 16944 6354 17004 6430
rect 17677 6427 17743 6430
rect 18137 6490 18203 6493
rect 19149 6490 19215 6493
rect 18137 6488 19215 6490
rect 18137 6432 18142 6488
rect 18198 6432 19154 6488
rect 19210 6432 19215 6488
rect 18137 6430 19215 6432
rect 18137 6427 18203 6430
rect 19149 6427 19215 6430
rect 7925 6352 10610 6354
rect 7925 6296 7930 6352
rect 7986 6296 8482 6352
rect 8538 6296 10610 6352
rect 7925 6294 10610 6296
rect 10918 6352 17004 6354
rect 10918 6296 10966 6352
rect 11022 6296 17004 6352
rect 10918 6294 17004 6296
rect 17493 6352 17559 6357
rect 18505 6354 18571 6357
rect 17493 6296 17498 6352
rect 17554 6296 17559 6352
rect 7925 6291 7991 6294
rect 8477 6291 8543 6294
rect 10918 6291 11027 6294
rect 17493 6291 17559 6296
rect 17726 6352 18571 6354
rect 17726 6296 18510 6352
rect 18566 6296 18571 6352
rect 17726 6294 18571 6296
rect 1025 6218 1091 6221
rect 10918 6218 10978 6291
rect 1025 6216 10978 6218
rect 1025 6160 1030 6216
rect 1086 6160 10978 6216
rect 1025 6158 10978 6160
rect 14273 6218 14339 6221
rect 14958 6218 14964 6220
rect 14273 6216 14964 6218
rect 14273 6160 14278 6216
rect 14334 6160 14964 6216
rect 14273 6158 14964 6160
rect 1025 6155 1091 6158
rect 14273 6155 14339 6158
rect 14958 6156 14964 6158
rect 15028 6156 15034 6220
rect 16573 6218 16639 6221
rect 17496 6218 17556 6291
rect 16573 6216 17556 6218
rect 16573 6160 16578 6216
rect 16634 6160 17556 6216
rect 16573 6158 17556 6160
rect 16573 6155 16639 6158
rect 4470 6020 4476 6084
rect 4540 6082 4546 6084
rect 6177 6082 6243 6085
rect 7046 6082 7052 6084
rect 4540 6080 7052 6082
rect 4540 6024 6182 6080
rect 6238 6024 7052 6080
rect 4540 6022 7052 6024
rect 4540 6020 4546 6022
rect 6177 6019 6243 6022
rect 7046 6020 7052 6022
rect 7116 6020 7122 6084
rect 7230 6020 7236 6084
rect 7300 6082 7306 6084
rect 7557 6082 7623 6085
rect 7300 6080 7623 6082
rect 7300 6024 7562 6080
rect 7618 6024 7623 6080
rect 7300 6022 7623 6024
rect 7300 6020 7306 6022
rect 7557 6019 7623 6022
rect 11513 6082 11579 6085
rect 11830 6082 11836 6084
rect 11513 6080 11836 6082
rect 11513 6024 11518 6080
rect 11574 6024 11836 6080
rect 11513 6022 11836 6024
rect 11513 6019 11579 6022
rect 11830 6020 11836 6022
rect 11900 6020 11906 6084
rect 15561 6082 15627 6085
rect 17726 6082 17786 6294
rect 18505 6291 18571 6294
rect 18781 6354 18847 6357
rect 22200 6354 23000 6384
rect 18781 6352 23000 6354
rect 18781 6296 18786 6352
rect 18842 6296 23000 6352
rect 18781 6294 23000 6296
rect 18781 6291 18847 6294
rect 22200 6264 23000 6294
rect 18321 6218 18387 6221
rect 18689 6218 18755 6221
rect 18321 6216 18755 6218
rect 18321 6160 18326 6216
rect 18382 6160 18694 6216
rect 18750 6160 18755 6216
rect 18321 6158 18755 6160
rect 18321 6155 18387 6158
rect 18689 6155 18755 6158
rect 15561 6080 17786 6082
rect 15561 6024 15566 6080
rect 15622 6024 17786 6080
rect 15561 6022 17786 6024
rect 18321 6082 18387 6085
rect 18873 6082 18939 6085
rect 18321 6080 18939 6082
rect 18321 6024 18326 6080
rect 18382 6024 18878 6080
rect 18934 6024 18939 6080
rect 18321 6022 18939 6024
rect 15561 6019 15627 6022
rect 18321 6019 18387 6022
rect 18873 6019 18939 6022
rect 3545 6016 3861 6017
rect 0 5946 800 5976
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 1117 5946 1183 5949
rect 2814 5946 2820 5948
rect 0 5944 2820 5946
rect 0 5888 1122 5944
rect 1178 5888 2820 5944
rect 0 5886 2820 5888
rect 0 5856 800 5886
rect 1117 5883 1183 5886
rect 2814 5884 2820 5886
rect 2884 5884 2890 5948
rect 4889 5946 4955 5949
rect 8334 5946 8340 5948
rect 4889 5944 8340 5946
rect 4889 5888 4894 5944
rect 4950 5888 8340 5944
rect 4889 5886 8340 5888
rect 4889 5883 4955 5886
rect 8334 5884 8340 5886
rect 8404 5884 8410 5948
rect 9305 5946 9371 5949
rect 11329 5946 11395 5949
rect 9305 5944 11395 5946
rect 9305 5888 9310 5944
rect 9366 5888 11334 5944
rect 11390 5888 11395 5944
rect 9305 5886 11395 5888
rect 9305 5883 9371 5886
rect 11329 5883 11395 5886
rect 11830 5884 11836 5948
rect 11900 5946 11906 5948
rect 11973 5946 12039 5949
rect 11900 5944 12039 5946
rect 11900 5888 11978 5944
rect 12034 5888 12039 5944
rect 11900 5886 12039 5888
rect 11900 5884 11906 5886
rect 11973 5883 12039 5886
rect 15561 5946 15627 5949
rect 15694 5946 15700 5948
rect 15561 5944 15700 5946
rect 15561 5888 15566 5944
rect 15622 5888 15700 5944
rect 15561 5886 15700 5888
rect 15561 5883 15627 5886
rect 15694 5884 15700 5886
rect 15764 5884 15770 5948
rect 16941 5946 17007 5949
rect 18321 5946 18387 5949
rect 22200 5946 23000 5976
rect 16941 5944 18387 5946
rect 16941 5888 16946 5944
rect 17002 5888 18326 5944
rect 18382 5888 18387 5944
rect 16941 5886 18387 5888
rect 16941 5883 17007 5886
rect 18321 5883 18387 5886
rect 19566 5886 23000 5946
rect 1485 5810 1551 5813
rect 4245 5810 4311 5813
rect 1485 5808 4311 5810
rect 1485 5752 1490 5808
rect 1546 5752 4250 5808
rect 4306 5752 4311 5808
rect 1485 5750 4311 5752
rect 1485 5747 1551 5750
rect 4245 5747 4311 5750
rect 5165 5810 5231 5813
rect 9121 5810 9187 5813
rect 14549 5810 14615 5813
rect 16113 5812 16179 5813
rect 5165 5808 14615 5810
rect 5165 5752 5170 5808
rect 5226 5752 9126 5808
rect 9182 5752 14554 5808
rect 14610 5752 14615 5808
rect 5165 5750 14615 5752
rect 5165 5747 5231 5750
rect 9121 5747 9187 5750
rect 14549 5747 14615 5750
rect 16062 5748 16068 5812
rect 16132 5810 16179 5812
rect 16297 5810 16363 5813
rect 18965 5810 19031 5813
rect 19566 5810 19626 5886
rect 22200 5856 23000 5886
rect 16132 5808 16224 5810
rect 16174 5752 16224 5808
rect 16132 5750 16224 5752
rect 16297 5808 19626 5810
rect 16297 5752 16302 5808
rect 16358 5752 18970 5808
rect 19026 5752 19626 5808
rect 16297 5750 19626 5752
rect 16132 5748 16179 5750
rect 16113 5747 16179 5748
rect 16297 5747 16363 5750
rect 18965 5747 19031 5750
rect 3366 5612 3372 5676
rect 3436 5674 3442 5676
rect 3785 5674 3851 5677
rect 3918 5674 3924 5676
rect 3436 5672 3924 5674
rect 3436 5616 3790 5672
rect 3846 5616 3924 5672
rect 3436 5614 3924 5616
rect 3436 5612 3442 5614
rect 3785 5611 3851 5614
rect 3918 5612 3924 5614
rect 3988 5612 3994 5676
rect 6361 5674 6427 5677
rect 10685 5674 10751 5677
rect 12433 5674 12499 5677
rect 12617 5674 12683 5677
rect 6361 5672 10751 5674
rect 6361 5616 6366 5672
rect 6422 5616 10690 5672
rect 10746 5616 10751 5672
rect 6361 5614 10751 5616
rect 6361 5611 6427 5614
rect 10685 5611 10751 5614
rect 11838 5672 12499 5674
rect 11838 5616 12438 5672
rect 12494 5616 12499 5672
rect 11838 5614 12499 5616
rect 0 5538 800 5568
rect 3182 5538 3188 5540
rect 0 5478 3188 5538
rect 0 5448 800 5478
rect 3182 5476 3188 5478
rect 3252 5476 3258 5540
rect 3509 5538 3575 5541
rect 5717 5538 5783 5541
rect 7649 5538 7715 5541
rect 3509 5536 5783 5538
rect 3509 5480 3514 5536
rect 3570 5480 5722 5536
rect 5778 5480 5783 5536
rect 3509 5478 5783 5480
rect 3509 5475 3575 5478
rect 5717 5475 5783 5478
rect 6548 5536 7715 5538
rect 6548 5480 7654 5536
rect 7710 5480 7715 5536
rect 6548 5478 7715 5480
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 1945 5402 2011 5405
rect 5809 5402 5875 5405
rect 1945 5400 5875 5402
rect 1945 5344 1950 5400
rect 2006 5344 5814 5400
rect 5870 5344 5875 5400
rect 1945 5342 5875 5344
rect 1945 5339 2011 5342
rect 5809 5339 5875 5342
rect 974 5204 980 5268
rect 1044 5266 1050 5268
rect 1209 5266 1275 5269
rect 1044 5264 1275 5266
rect 1044 5208 1214 5264
rect 1270 5208 1275 5264
rect 1044 5206 1275 5208
rect 1044 5204 1050 5206
rect 1209 5203 1275 5206
rect 3417 5266 3483 5269
rect 6548 5266 6608 5478
rect 7649 5475 7715 5478
rect 8753 5538 8819 5541
rect 11053 5538 11119 5541
rect 8753 5536 11119 5538
rect 8753 5480 8758 5536
rect 8814 5480 11058 5536
rect 11114 5480 11119 5536
rect 8753 5478 11119 5480
rect 8753 5475 8819 5478
rect 11053 5475 11119 5478
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 7557 5404 7623 5405
rect 7557 5402 7604 5404
rect 7512 5400 7604 5402
rect 7512 5344 7562 5400
rect 7512 5342 7604 5344
rect 7557 5340 7604 5342
rect 7668 5340 7674 5404
rect 9673 5402 9739 5405
rect 7974 5400 9739 5402
rect 7974 5344 9678 5400
rect 9734 5344 9739 5400
rect 7974 5342 9739 5344
rect 7557 5339 7623 5340
rect 7974 5266 8034 5342
rect 9673 5339 9739 5342
rect 3417 5264 6608 5266
rect 3417 5208 3422 5264
rect 3478 5208 6608 5264
rect 3417 5206 6608 5208
rect 7606 5206 8034 5266
rect 3417 5203 3483 5206
rect 0 5130 800 5160
rect 2221 5130 2287 5133
rect 0 5128 2287 5130
rect 0 5072 2226 5128
rect 2282 5072 2287 5128
rect 0 5070 2287 5072
rect 0 5040 800 5070
rect 2221 5067 2287 5070
rect 2405 5130 2471 5133
rect 3182 5130 3188 5132
rect 2405 5128 3188 5130
rect 2405 5072 2410 5128
rect 2466 5072 3188 5128
rect 2405 5070 3188 5072
rect 2405 5067 2471 5070
rect 3182 5068 3188 5070
rect 3252 5068 3258 5132
rect 3785 5130 3851 5133
rect 3785 5128 5458 5130
rect 3785 5072 3790 5128
rect 3846 5072 5458 5128
rect 3785 5070 5458 5072
rect 3785 5067 3851 5070
rect 1945 4994 2011 4997
rect 2446 4994 2452 4996
rect 1945 4992 2452 4994
rect 1945 4936 1950 4992
rect 2006 4936 2452 4992
rect 1945 4934 2452 4936
rect 1945 4931 2011 4934
rect 2446 4932 2452 4934
rect 2516 4932 2522 4996
rect 4838 4932 4844 4996
rect 4908 4994 4914 4996
rect 5257 4994 5323 4997
rect 4908 4992 5323 4994
rect 4908 4936 5262 4992
rect 5318 4936 5323 4992
rect 4908 4934 5323 4936
rect 5398 4994 5458 5070
rect 5574 5068 5580 5132
rect 5644 5130 5650 5132
rect 6453 5130 6519 5133
rect 7606 5130 7666 5206
rect 8150 5204 8156 5268
rect 8220 5266 8226 5268
rect 11838 5266 11898 5614
rect 12433 5611 12499 5614
rect 12574 5672 12683 5674
rect 12574 5616 12622 5672
rect 12678 5616 12683 5672
rect 12574 5611 12683 5616
rect 12893 5674 12959 5677
rect 19793 5674 19859 5677
rect 12893 5672 19859 5674
rect 12893 5616 12898 5672
rect 12954 5616 19798 5672
rect 19854 5616 19859 5672
rect 12893 5614 19859 5616
rect 12893 5611 12959 5614
rect 19793 5611 19859 5614
rect 21590 5614 22202 5674
rect 12014 5476 12020 5540
rect 12084 5538 12090 5540
rect 12574 5538 12634 5611
rect 12084 5478 12634 5538
rect 13353 5538 13419 5541
rect 16297 5538 16363 5541
rect 13353 5536 16363 5538
rect 13353 5480 13358 5536
rect 13414 5480 16302 5536
rect 16358 5480 16363 5536
rect 13353 5478 16363 5480
rect 12084 5476 12090 5478
rect 13353 5475 13419 5478
rect 16297 5475 16363 5478
rect 18413 5538 18479 5541
rect 21449 5538 21515 5541
rect 21590 5538 21650 5614
rect 18413 5536 21650 5538
rect 18413 5480 18418 5536
rect 18474 5480 21454 5536
rect 21510 5480 21650 5536
rect 18413 5478 21650 5480
rect 22142 5568 22202 5614
rect 22142 5478 23000 5568
rect 18413 5475 18479 5478
rect 21449 5475 21515 5478
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 22200 5448 23000 5478
rect 21738 5407 22054 5408
rect 11973 5402 12039 5405
rect 14089 5402 14155 5405
rect 15193 5404 15259 5405
rect 11973 5400 14155 5402
rect 11973 5344 11978 5400
rect 12034 5344 14094 5400
rect 14150 5344 14155 5400
rect 11973 5342 14155 5344
rect 11973 5339 12039 5342
rect 14089 5339 14155 5342
rect 15142 5340 15148 5404
rect 15212 5402 15259 5404
rect 15212 5400 15394 5402
rect 15254 5344 15394 5400
rect 15212 5342 15394 5344
rect 15212 5340 15259 5342
rect 15193 5339 15259 5340
rect 15193 5266 15259 5269
rect 8220 5206 11898 5266
rect 11976 5264 15259 5266
rect 11976 5208 15198 5264
rect 15254 5208 15259 5264
rect 11976 5206 15259 5208
rect 15334 5266 15394 5342
rect 16297 5266 16363 5269
rect 16941 5266 17007 5269
rect 15334 5264 17007 5266
rect 15334 5208 16302 5264
rect 16358 5208 16946 5264
rect 17002 5208 17007 5264
rect 15334 5206 17007 5208
rect 8220 5204 8226 5206
rect 5644 5128 7666 5130
rect 5644 5072 6458 5128
rect 6514 5072 7666 5128
rect 5644 5070 7666 5072
rect 8109 5130 8175 5133
rect 11329 5130 11395 5133
rect 8109 5128 11395 5130
rect 8109 5072 8114 5128
rect 8170 5072 11334 5128
rect 11390 5072 11395 5128
rect 8109 5070 11395 5072
rect 5644 5068 5650 5070
rect 6453 5067 6519 5070
rect 8109 5067 8175 5070
rect 11329 5067 11395 5070
rect 7598 4994 7604 4996
rect 5398 4934 7604 4994
rect 4908 4932 4914 4934
rect 5257 4931 5323 4934
rect 7598 4932 7604 4934
rect 7668 4994 7674 4996
rect 8477 4994 8543 4997
rect 7668 4992 8543 4994
rect 7668 4936 8482 4992
rect 8538 4936 8543 4992
rect 7668 4934 8543 4936
rect 7668 4932 7674 4934
rect 8477 4931 8543 4934
rect 9673 4994 9739 4997
rect 11976 4994 12036 5206
rect 15193 5203 15259 5206
rect 16297 5203 16363 5206
rect 16941 5203 17007 5206
rect 12433 5130 12499 5133
rect 12985 5130 13051 5133
rect 17309 5130 17375 5133
rect 21081 5130 21147 5133
rect 12433 5128 17375 5130
rect 12433 5072 12438 5128
rect 12494 5072 12990 5128
rect 13046 5072 17314 5128
rect 17370 5072 17375 5128
rect 12433 5070 17375 5072
rect 12433 5067 12499 5070
rect 12985 5067 13051 5070
rect 17309 5067 17375 5070
rect 19014 5128 21147 5130
rect 19014 5072 21086 5128
rect 21142 5072 21147 5128
rect 19014 5070 21147 5072
rect 9673 4992 12036 4994
rect 9673 4936 9678 4992
rect 9734 4936 12036 4992
rect 9673 4934 12036 4936
rect 12341 4994 12407 4997
rect 13353 4994 13419 4997
rect 12341 4992 13419 4994
rect 12341 4936 12346 4992
rect 12402 4936 13358 4992
rect 13414 4936 13419 4992
rect 12341 4934 13419 4936
rect 9673 4931 9739 4934
rect 12341 4931 12407 4934
rect 13353 4931 13419 4934
rect 14365 4994 14431 4997
rect 15285 4994 15351 4997
rect 17585 4994 17651 4997
rect 14365 4992 17651 4994
rect 14365 4936 14370 4992
rect 14426 4936 15290 4992
rect 15346 4936 17590 4992
rect 17646 4936 17651 4992
rect 14365 4934 17651 4936
rect 14365 4931 14431 4934
rect 15285 4931 15351 4934
rect 17585 4931 17651 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 1301 4858 1367 4861
rect 4337 4858 4403 4861
rect 7281 4858 7347 4861
rect 8150 4858 8156 4860
rect 1301 4856 2790 4858
rect 1301 4800 1306 4856
rect 1362 4800 2790 4856
rect 1301 4798 2790 4800
rect 1301 4795 1367 4798
rect 0 4722 800 4752
rect 974 4722 980 4724
rect 0 4662 980 4722
rect 0 4632 800 4662
rect 974 4660 980 4662
rect 1044 4660 1050 4724
rect 2730 4722 2790 4798
rect 4337 4856 8156 4858
rect 4337 4800 4342 4856
rect 4398 4800 7286 4856
rect 7342 4800 8156 4856
rect 4337 4798 8156 4800
rect 4337 4795 4403 4798
rect 7281 4795 7347 4798
rect 8150 4796 8156 4798
rect 8220 4796 8226 4860
rect 10501 4858 10567 4861
rect 11789 4858 11855 4861
rect 10501 4856 11855 4858
rect 10501 4800 10506 4856
rect 10562 4800 11794 4856
rect 11850 4800 11855 4856
rect 10501 4798 11855 4800
rect 10501 4795 10567 4798
rect 11789 4795 11855 4798
rect 15193 4858 15259 4861
rect 19014 4858 19074 5070
rect 21081 5067 21147 5070
rect 21541 5130 21607 5133
rect 22200 5130 23000 5160
rect 21541 5128 23000 5130
rect 21541 5072 21546 5128
rect 21602 5072 23000 5128
rect 21541 5070 23000 5072
rect 21541 5067 21607 5070
rect 22200 5040 23000 5070
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 15193 4856 19074 4858
rect 15193 4800 15198 4856
rect 15254 4800 19074 4856
rect 15193 4798 19074 4800
rect 15193 4795 15259 4798
rect 4245 4722 4311 4725
rect 2730 4720 4311 4722
rect 2730 4664 4250 4720
rect 4306 4664 4311 4720
rect 2730 4662 4311 4664
rect 4245 4659 4311 4662
rect 4797 4722 4863 4725
rect 5257 4722 5323 4725
rect 4797 4720 5323 4722
rect 4797 4664 4802 4720
rect 4858 4664 5262 4720
rect 5318 4664 5323 4720
rect 4797 4662 5323 4664
rect 4797 4659 4863 4662
rect 5257 4659 5323 4662
rect 6085 4722 6151 4725
rect 12934 4722 12940 4724
rect 6085 4720 12940 4722
rect 6085 4664 6090 4720
rect 6146 4664 12940 4720
rect 6085 4662 12940 4664
rect 6085 4659 6151 4662
rect 12934 4660 12940 4662
rect 13004 4660 13010 4724
rect 20437 4722 20503 4725
rect 21081 4722 21147 4725
rect 22200 4722 23000 4752
rect 20437 4720 23000 4722
rect 20437 4664 20442 4720
rect 20498 4664 21086 4720
rect 21142 4664 23000 4720
rect 20437 4662 23000 4664
rect 20437 4659 20503 4662
rect 21081 4659 21147 4662
rect 22200 4632 23000 4662
rect 2405 4586 2471 4589
rect 5717 4586 5783 4589
rect 6678 4586 6684 4588
rect 2405 4584 6684 4586
rect 2405 4528 2410 4584
rect 2466 4528 5722 4584
rect 5778 4528 6684 4584
rect 2405 4526 6684 4528
rect 2405 4523 2471 4526
rect 5717 4523 5783 4526
rect 6678 4524 6684 4526
rect 6748 4524 6754 4588
rect 6913 4586 6979 4589
rect 13353 4586 13419 4589
rect 13486 4586 13492 4588
rect 6913 4584 13492 4586
rect 6913 4528 6918 4584
rect 6974 4528 13358 4584
rect 13414 4528 13492 4584
rect 6913 4526 13492 4528
rect 6913 4523 6979 4526
rect 13353 4523 13419 4526
rect 13486 4524 13492 4526
rect 13556 4524 13562 4588
rect 2497 4450 2563 4453
rect 4102 4450 4108 4452
rect 2497 4448 4108 4450
rect 2497 4392 2502 4448
rect 2558 4392 4108 4448
rect 2497 4390 4108 4392
rect 2497 4387 2563 4390
rect 4102 4388 4108 4390
rect 4172 4388 4178 4452
rect 4797 4450 4863 4453
rect 5390 4450 5396 4452
rect 4797 4448 5396 4450
rect 4797 4392 4802 4448
rect 4858 4392 5396 4448
rect 4797 4390 5396 4392
rect 4797 4387 4863 4390
rect 5390 4388 5396 4390
rect 5460 4388 5466 4452
rect 17534 4388 17540 4452
rect 17604 4450 17610 4452
rect 18505 4450 18571 4453
rect 17604 4448 18571 4450
rect 17604 4392 18510 4448
rect 18566 4392 18571 4448
rect 17604 4390 18571 4392
rect 17604 4388 17610 4390
rect 18505 4387 18571 4390
rect 6144 4384 6460 4385
rect 0 4314 800 4344
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 3417 4314 3483 4317
rect 0 4312 3483 4314
rect 0 4256 3422 4312
rect 3478 4256 3483 4312
rect 0 4254 3483 4256
rect 0 4224 800 4254
rect 3417 4251 3483 4254
rect 4102 4252 4108 4316
rect 4172 4314 4178 4316
rect 4889 4314 4955 4317
rect 4172 4312 4955 4314
rect 4172 4256 4894 4312
rect 4950 4256 4955 4312
rect 4172 4254 4955 4256
rect 4172 4252 4178 4254
rect 4889 4251 4955 4254
rect 7281 4314 7347 4317
rect 9305 4314 9371 4317
rect 7281 4312 9371 4314
rect 7281 4256 7286 4312
rect 7342 4256 9310 4312
rect 9366 4256 9371 4312
rect 7281 4254 9371 4256
rect 7281 4251 7347 4254
rect 9305 4251 9371 4254
rect 11881 4314 11947 4317
rect 15193 4314 15259 4317
rect 22200 4314 23000 4344
rect 11881 4312 15259 4314
rect 11881 4256 11886 4312
rect 11942 4256 15198 4312
rect 15254 4256 15259 4312
rect 11881 4254 15259 4256
rect 11881 4251 11947 4254
rect 15193 4251 15259 4254
rect 2221 4178 2287 4181
rect 14406 4178 14412 4180
rect 2221 4176 14412 4178
rect 2221 4120 2226 4176
rect 2282 4120 14412 4176
rect 2221 4118 14412 4120
rect 2221 4115 2287 4118
rect 14406 4116 14412 4118
rect 14476 4116 14482 4180
rect 15196 4178 15256 4251
rect 22142 4224 23000 4314
rect 16941 4178 17007 4181
rect 15196 4176 17007 4178
rect 15196 4120 16946 4176
rect 17002 4120 17007 4176
rect 15196 4118 17007 4120
rect 16941 4115 17007 4118
rect 22001 4178 22067 4181
rect 22142 4178 22202 4224
rect 22001 4176 22202 4178
rect 22001 4120 22006 4176
rect 22062 4120 22202 4176
rect 22001 4118 22202 4120
rect 22001 4115 22067 4118
rect 5022 4042 5028 4044
rect 2454 3982 5028 4042
rect 0 3906 800 3936
rect 2454 3906 2514 3982
rect 5022 3980 5028 3982
rect 5092 3980 5098 4044
rect 5942 3980 5948 4044
rect 6012 4042 6018 4044
rect 6361 4042 6427 4045
rect 6012 4040 6427 4042
rect 6012 3984 6366 4040
rect 6422 3984 6427 4040
rect 6012 3982 6427 3984
rect 6012 3980 6018 3982
rect 6361 3979 6427 3982
rect 6678 3980 6684 4044
rect 6748 4042 6754 4044
rect 10133 4042 10199 4045
rect 6748 4040 10199 4042
rect 6748 3984 10138 4040
rect 10194 3984 10199 4040
rect 6748 3982 10199 3984
rect 6748 3980 6754 3982
rect 10133 3979 10199 3982
rect 11881 4042 11947 4045
rect 12566 4042 12572 4044
rect 11881 4040 12572 4042
rect 11881 3984 11886 4040
rect 11942 3984 12572 4040
rect 11881 3982 12572 3984
rect 11881 3979 11947 3982
rect 12566 3980 12572 3982
rect 12636 3980 12642 4044
rect 15561 4042 15627 4045
rect 19425 4042 19491 4045
rect 13724 4040 19491 4042
rect 13724 3984 15566 4040
rect 15622 3984 19430 4040
rect 19486 3984 19491 4040
rect 13724 3982 19491 3984
rect 0 3846 2514 3906
rect 0 3816 800 3846
rect 2630 3844 2636 3908
rect 2700 3906 2706 3908
rect 3325 3906 3391 3909
rect 7782 3906 7788 3908
rect 2700 3904 3391 3906
rect 2700 3848 3330 3904
rect 3386 3848 3391 3904
rect 2700 3846 3391 3848
rect 2700 3844 2706 3846
rect 3325 3843 3391 3846
rect 5950 3846 7788 3906
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 974 3708 980 3772
rect 1044 3770 1050 3772
rect 1485 3770 1551 3773
rect 1044 3768 1551 3770
rect 1044 3712 1490 3768
rect 1546 3712 1551 3768
rect 1044 3710 1551 3712
rect 1044 3708 1050 3710
rect 1485 3707 1551 3710
rect 4470 3634 4476 3636
rect 2270 3574 4476 3634
rect 0 3498 800 3528
rect 2270 3498 2330 3574
rect 4470 3572 4476 3574
rect 4540 3572 4546 3636
rect 0 3438 2330 3498
rect 2589 3498 2655 3501
rect 4654 3498 4660 3500
rect 2589 3496 4660 3498
rect 2589 3440 2594 3496
rect 2650 3440 4660 3496
rect 2589 3438 4660 3440
rect 0 3408 800 3438
rect 2589 3435 2655 3438
rect 4654 3436 4660 3438
rect 4724 3436 4730 3500
rect 3141 3362 3207 3365
rect 5950 3362 6010 3846
rect 7782 3844 7788 3846
rect 7852 3844 7858 3908
rect 10869 3906 10935 3909
rect 13169 3906 13235 3909
rect 10869 3904 13235 3906
rect 10869 3848 10874 3904
rect 10930 3848 13174 3904
rect 13230 3848 13235 3904
rect 10869 3846 13235 3848
rect 10869 3843 10935 3846
rect 13169 3843 13235 3846
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 6269 3770 6335 3773
rect 7966 3770 7972 3772
rect 6269 3768 7972 3770
rect 6269 3712 6274 3768
rect 6330 3712 7972 3768
rect 6269 3710 7972 3712
rect 6269 3707 6335 3710
rect 7966 3708 7972 3710
rect 8036 3708 8042 3772
rect 9254 3708 9260 3772
rect 9324 3770 9330 3772
rect 13724 3770 13784 3982
rect 15561 3979 15627 3982
rect 19425 3979 19491 3982
rect 20253 4044 20319 4045
rect 20253 4040 20300 4044
rect 20364 4042 20370 4044
rect 20253 3984 20258 4040
rect 20253 3980 20300 3984
rect 20364 3982 20410 4042
rect 20364 3980 20370 3982
rect 20253 3979 20319 3980
rect 14457 3906 14523 3909
rect 14457 3904 14658 3906
rect 14457 3848 14462 3904
rect 14518 3848 14658 3904
rect 14457 3846 14658 3848
rect 14457 3843 14523 3846
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 9324 3710 13784 3770
rect 14598 3770 14658 3846
rect 18822 3844 18828 3908
rect 18892 3906 18898 3908
rect 18965 3906 19031 3909
rect 18892 3904 19031 3906
rect 18892 3848 18970 3904
rect 19026 3848 19031 3904
rect 18892 3846 19031 3848
rect 18892 3844 18898 3846
rect 18965 3843 19031 3846
rect 20345 3906 20411 3909
rect 20478 3906 20484 3908
rect 20345 3904 20484 3906
rect 20345 3848 20350 3904
rect 20406 3848 20484 3904
rect 20345 3846 20484 3848
rect 20345 3843 20411 3846
rect 20478 3844 20484 3846
rect 20548 3844 20554 3908
rect 22001 3906 22067 3909
rect 22200 3906 23000 3936
rect 22001 3904 23000 3906
rect 22001 3848 22006 3904
rect 22062 3848 23000 3904
rect 22001 3846 23000 3848
rect 22001 3843 22067 3846
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 22200 3816 23000 3846
rect 19139 3775 19455 3776
rect 14733 3770 14799 3773
rect 14598 3768 14799 3770
rect 14598 3712 14738 3768
rect 14794 3712 14799 3768
rect 14598 3710 14799 3712
rect 9324 3708 9330 3710
rect 14733 3707 14799 3710
rect 19742 3708 19748 3772
rect 19812 3770 19818 3772
rect 19885 3770 19951 3773
rect 19812 3768 19951 3770
rect 19812 3712 19890 3768
rect 19946 3712 19951 3768
rect 19812 3710 19951 3712
rect 19812 3708 19818 3710
rect 19885 3707 19951 3710
rect 20621 3770 20687 3773
rect 22001 3770 22067 3773
rect 20621 3768 22067 3770
rect 20621 3712 20626 3768
rect 20682 3712 22006 3768
rect 22062 3712 22067 3768
rect 20621 3710 22067 3712
rect 20621 3707 20687 3710
rect 22001 3707 22067 3710
rect 6453 3634 6519 3637
rect 6913 3634 6979 3637
rect 11830 3634 11836 3636
rect 6453 3632 11836 3634
rect 6453 3576 6458 3632
rect 6514 3576 6918 3632
rect 6974 3576 11836 3632
rect 6453 3574 11836 3576
rect 6453 3571 6519 3574
rect 6913 3571 6979 3574
rect 11830 3572 11836 3574
rect 11900 3572 11906 3636
rect 12709 3634 12775 3637
rect 21357 3634 21423 3637
rect 12709 3632 21423 3634
rect 12709 3576 12714 3632
rect 12770 3576 21362 3632
rect 21418 3576 21423 3632
rect 12709 3574 21423 3576
rect 12709 3571 12775 3574
rect 21357 3571 21423 3574
rect 6085 3498 6151 3501
rect 6085 3496 7298 3498
rect 6085 3440 6090 3496
rect 6146 3440 7298 3496
rect 6085 3438 7298 3440
rect 6085 3435 6151 3438
rect 3141 3360 6010 3362
rect 3141 3304 3146 3360
rect 3202 3304 6010 3360
rect 3141 3302 6010 3304
rect 3141 3299 3207 3302
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 1393 3226 1459 3229
rect 2497 3226 2563 3229
rect 5533 3226 5599 3229
rect 1393 3224 5599 3226
rect 1393 3168 1398 3224
rect 1454 3168 2502 3224
rect 2558 3168 5538 3224
rect 5594 3168 5599 3224
rect 1393 3166 5599 3168
rect 1393 3163 1459 3166
rect 2497 3163 2563 3166
rect 5533 3163 5599 3166
rect 0 3090 800 3120
rect 3785 3090 3851 3093
rect 0 3088 3851 3090
rect 0 3032 3790 3088
rect 3846 3032 3851 3088
rect 0 3030 3851 3032
rect 0 3000 800 3030
rect 3785 3027 3851 3030
rect 3325 2956 3391 2957
rect 3325 2954 3372 2956
rect 3280 2952 3372 2954
rect 3280 2896 3330 2952
rect 3280 2894 3372 2896
rect 3325 2892 3372 2894
rect 3436 2892 3442 2956
rect 3509 2954 3575 2957
rect 4521 2954 4587 2957
rect 3509 2952 4587 2954
rect 3509 2896 3514 2952
rect 3570 2896 4526 2952
rect 4582 2896 4587 2952
rect 3509 2894 4587 2896
rect 3325 2891 3391 2892
rect 3509 2891 3575 2894
rect 4521 2891 4587 2894
rect 4981 2954 5047 2957
rect 5206 2954 5212 2956
rect 4981 2952 5212 2954
rect 4981 2896 4986 2952
rect 5042 2896 5212 2952
rect 4981 2894 5212 2896
rect 4981 2891 5047 2894
rect 5206 2892 5212 2894
rect 5276 2892 5282 2956
rect 7238 2818 7298 3438
rect 7966 3436 7972 3500
rect 8036 3498 8042 3500
rect 9254 3498 9260 3500
rect 8036 3438 9260 3498
rect 8036 3436 8042 3438
rect 9254 3436 9260 3438
rect 9324 3436 9330 3500
rect 10133 3498 10199 3501
rect 12157 3498 12223 3501
rect 14733 3498 14799 3501
rect 10133 3496 11898 3498
rect 10133 3440 10138 3496
rect 10194 3440 11898 3496
rect 10133 3438 11898 3440
rect 10133 3435 10199 3438
rect 7373 3362 7439 3365
rect 11838 3362 11898 3438
rect 12157 3496 14799 3498
rect 12157 3440 12162 3496
rect 12218 3440 14738 3496
rect 14794 3440 14799 3496
rect 12157 3438 14799 3440
rect 12157 3435 12223 3438
rect 14733 3435 14799 3438
rect 18965 3498 19031 3501
rect 22200 3498 23000 3528
rect 18965 3496 23000 3498
rect 18965 3440 18970 3496
rect 19026 3440 23000 3496
rect 18965 3438 23000 3440
rect 18965 3435 19031 3438
rect 22200 3408 23000 3438
rect 15694 3362 15700 3364
rect 7373 3360 11162 3362
rect 7373 3304 7378 3360
rect 7434 3304 11162 3360
rect 7373 3302 11162 3304
rect 11838 3302 15700 3362
rect 7373 3299 7439 3302
rect 11102 3229 11162 3302
rect 15694 3300 15700 3302
rect 15764 3300 15770 3364
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 9990 3164 9996 3228
rect 10060 3226 10066 3228
rect 10133 3226 10199 3229
rect 10060 3224 10199 3226
rect 10060 3168 10138 3224
rect 10194 3168 10199 3224
rect 10060 3166 10199 3168
rect 11102 3224 11211 3229
rect 11102 3168 11150 3224
rect 11206 3168 11211 3224
rect 11102 3166 11211 3168
rect 10060 3164 10066 3166
rect 10133 3163 10199 3166
rect 11145 3163 11211 3166
rect 12433 3226 12499 3229
rect 14181 3226 14247 3229
rect 12433 3224 14247 3226
rect 12433 3168 12438 3224
rect 12494 3168 14186 3224
rect 14242 3168 14247 3224
rect 12433 3166 14247 3168
rect 12433 3163 12499 3166
rect 14181 3163 14247 3166
rect 7741 3090 7807 3093
rect 8569 3090 8635 3093
rect 17401 3090 17467 3093
rect 7741 3088 8172 3090
rect 7741 3032 7746 3088
rect 7802 3032 8172 3088
rect 7741 3030 8172 3032
rect 7741 3027 7807 3030
rect 8112 2957 8172 3030
rect 8569 3088 17467 3090
rect 8569 3032 8574 3088
rect 8630 3032 17406 3088
rect 17462 3032 17467 3088
rect 8569 3030 17467 3032
rect 8569 3027 8635 3030
rect 17401 3027 17467 3030
rect 17902 3028 17908 3092
rect 17972 3090 17978 3092
rect 18045 3090 18111 3093
rect 17972 3088 18111 3090
rect 17972 3032 18050 3088
rect 18106 3032 18111 3088
rect 17972 3030 18111 3032
rect 17972 3028 17978 3030
rect 18045 3027 18111 3030
rect 19701 3090 19767 3093
rect 22200 3090 23000 3120
rect 19701 3088 23000 3090
rect 19701 3032 19706 3088
rect 19762 3032 23000 3088
rect 19701 3030 23000 3032
rect 19701 3027 19767 3030
rect 22200 3000 23000 3030
rect 8109 2952 8175 2957
rect 10726 2954 10732 2956
rect 8109 2896 8114 2952
rect 8170 2896 8175 2952
rect 8109 2891 8175 2896
rect 8526 2894 10732 2954
rect 8526 2818 8586 2894
rect 10726 2892 10732 2894
rect 10796 2892 10802 2956
rect 12065 2954 12131 2957
rect 13905 2954 13971 2957
rect 12065 2952 13971 2954
rect 12065 2896 12070 2952
rect 12126 2896 13910 2952
rect 13966 2896 13971 2952
rect 12065 2894 13971 2896
rect 12065 2891 12131 2894
rect 13905 2891 13971 2894
rect 14365 2954 14431 2957
rect 14590 2954 14596 2956
rect 14365 2952 14596 2954
rect 14365 2896 14370 2952
rect 14426 2896 14596 2952
rect 14365 2894 14596 2896
rect 14365 2891 14431 2894
rect 14590 2892 14596 2894
rect 14660 2954 14666 2956
rect 17217 2954 17283 2957
rect 14660 2952 17283 2954
rect 14660 2896 17222 2952
rect 17278 2896 17283 2952
rect 14660 2894 17283 2896
rect 14660 2892 14666 2894
rect 17217 2891 17283 2894
rect 17401 2954 17467 2957
rect 19701 2954 19767 2957
rect 17401 2952 19767 2954
rect 17401 2896 17406 2952
rect 17462 2896 19706 2952
rect 19762 2896 19767 2952
rect 17401 2894 19767 2896
rect 17401 2891 17467 2894
rect 19701 2891 19767 2894
rect 7238 2758 8586 2818
rect 15561 2818 15627 2821
rect 16113 2818 16179 2821
rect 15561 2816 16179 2818
rect 15561 2760 15566 2816
rect 15622 2760 16118 2816
rect 16174 2760 16179 2816
rect 15561 2758 16179 2760
rect 15561 2755 15627 2758
rect 16113 2755 16179 2758
rect 3545 2752 3861 2753
rect 0 2682 800 2712
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 2865 2682 2931 2685
rect 4705 2682 4771 2685
rect 5574 2682 5580 2684
rect 0 2680 3434 2682
rect 0 2624 2870 2680
rect 2926 2624 3434 2680
rect 0 2622 3434 2624
rect 0 2592 800 2622
rect 2865 2619 2931 2622
rect 1158 2484 1164 2548
rect 1228 2546 1234 2548
rect 2221 2546 2287 2549
rect 3141 2546 3207 2549
rect 1228 2544 3207 2546
rect 1228 2488 2226 2544
rect 2282 2488 3146 2544
rect 3202 2488 3207 2544
rect 1228 2486 3207 2488
rect 3374 2546 3434 2622
rect 4705 2680 5580 2682
rect 4705 2624 4710 2680
rect 4766 2624 5580 2680
rect 4705 2622 5580 2624
rect 4705 2619 4771 2622
rect 5574 2620 5580 2622
rect 5644 2620 5650 2684
rect 6862 2620 6868 2684
rect 6932 2682 6938 2684
rect 8201 2682 8267 2685
rect 6932 2680 8267 2682
rect 6932 2624 8206 2680
rect 8262 2624 8267 2680
rect 6932 2622 8267 2624
rect 6932 2620 6938 2622
rect 8201 2619 8267 2622
rect 10174 2620 10180 2684
rect 10244 2682 10250 2684
rect 13721 2682 13787 2685
rect 10244 2680 13787 2682
rect 10244 2624 13726 2680
rect 13782 2624 13787 2680
rect 10244 2622 13787 2624
rect 10244 2620 10250 2622
rect 13721 2619 13787 2622
rect 20069 2682 20135 2685
rect 22200 2682 23000 2712
rect 20069 2680 23000 2682
rect 20069 2624 20074 2680
rect 20130 2624 23000 2680
rect 20069 2622 23000 2624
rect 20069 2619 20135 2622
rect 22200 2592 23000 2622
rect 3374 2486 6746 2546
rect 1228 2484 1234 2486
rect 2221 2483 2287 2486
rect 3141 2483 3207 2486
rect 3417 2410 3483 2413
rect 1166 2408 3483 2410
rect 1166 2352 3422 2408
rect 3478 2352 3483 2408
rect 1166 2350 3483 2352
rect 0 2274 800 2304
rect 1166 2274 1226 2350
rect 3417 2347 3483 2350
rect 0 2214 1226 2274
rect 0 2184 800 2214
rect 1342 2212 1348 2276
rect 1412 2274 1418 2276
rect 3693 2274 3759 2277
rect 1412 2272 3759 2274
rect 1412 2216 3698 2272
rect 3754 2216 3759 2272
rect 1412 2214 3759 2216
rect 6686 2274 6746 2486
rect 7230 2484 7236 2548
rect 7300 2546 7306 2548
rect 7373 2546 7439 2549
rect 7557 2548 7623 2549
rect 7557 2546 7604 2548
rect 7300 2544 7439 2546
rect 7300 2488 7378 2544
rect 7434 2488 7439 2544
rect 7300 2486 7439 2488
rect 7512 2544 7604 2546
rect 7512 2488 7562 2544
rect 7512 2486 7604 2488
rect 7300 2484 7306 2486
rect 7373 2483 7439 2486
rect 7557 2484 7604 2486
rect 7668 2484 7674 2548
rect 10133 2546 10199 2549
rect 11094 2546 11100 2548
rect 10133 2544 11100 2546
rect 10133 2488 10138 2544
rect 10194 2488 11100 2544
rect 10133 2486 11100 2488
rect 7557 2483 7623 2484
rect 10133 2483 10199 2486
rect 11094 2484 11100 2486
rect 11164 2484 11170 2548
rect 7414 2348 7420 2412
rect 7484 2410 7490 2412
rect 10685 2410 10751 2413
rect 12198 2410 12204 2412
rect 7484 2408 10751 2410
rect 7484 2352 10690 2408
rect 10746 2352 10751 2408
rect 7484 2350 10751 2352
rect 7484 2348 7490 2350
rect 10685 2347 10751 2350
rect 10918 2350 12204 2410
rect 10918 2274 10978 2350
rect 12198 2348 12204 2350
rect 12268 2348 12274 2412
rect 20713 2410 20779 2413
rect 20713 2408 22202 2410
rect 20713 2352 20718 2408
rect 20774 2352 22202 2408
rect 20713 2350 22202 2352
rect 20713 2347 20779 2350
rect 6686 2214 10978 2274
rect 22142 2304 22202 2350
rect 22142 2214 23000 2304
rect 1412 2212 1418 2214
rect 3693 2211 3759 2214
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 22200 2184 23000 2214
rect 21738 2143 22054 2144
rect 7373 2002 7439 2005
rect 17350 2002 17356 2004
rect 7373 2000 17356 2002
rect 7373 1944 7378 2000
rect 7434 1944 17356 2000
rect 7373 1942 17356 1944
rect 7373 1939 7439 1942
rect 17350 1940 17356 1942
rect 17420 1940 17426 2004
rect 0 1866 800 1896
rect 3785 1866 3851 1869
rect 0 1864 3851 1866
rect 0 1808 3790 1864
rect 3846 1808 3851 1864
rect 0 1806 3851 1808
rect 0 1776 800 1806
rect 3785 1803 3851 1806
rect 3969 1866 4035 1869
rect 10593 1866 10659 1869
rect 3969 1864 10659 1866
rect 3969 1808 3974 1864
rect 4030 1808 10598 1864
rect 10654 1808 10659 1864
rect 3969 1806 10659 1808
rect 3969 1803 4035 1806
rect 10593 1803 10659 1806
rect 19793 1866 19859 1869
rect 22200 1866 23000 1896
rect 19793 1864 23000 1866
rect 19793 1808 19798 1864
rect 19854 1808 23000 1864
rect 19793 1806 23000 1808
rect 19793 1803 19859 1806
rect 22200 1776 23000 1806
rect 6637 1730 6703 1733
rect 10358 1730 10364 1732
rect 6637 1728 10364 1730
rect 6637 1672 6642 1728
rect 6698 1672 10364 1728
rect 6637 1670 10364 1672
rect 6637 1667 6703 1670
rect 10358 1668 10364 1670
rect 10428 1668 10434 1732
rect 0 1458 800 1488
rect 9438 1458 9444 1460
rect 0 1398 9444 1458
rect 0 1368 800 1398
rect 9438 1396 9444 1398
rect 9508 1396 9514 1460
rect 20805 1458 20871 1461
rect 22200 1458 23000 1488
rect 20805 1456 23000 1458
rect 20805 1400 20810 1456
rect 20866 1400 23000 1456
rect 20805 1398 23000 1400
rect 20805 1395 20871 1398
rect 22200 1368 23000 1398
rect 5390 1260 5396 1324
rect 5460 1322 5466 1324
rect 12014 1322 12020 1324
rect 5460 1262 12020 1322
rect 5460 1260 5466 1262
rect 12014 1260 12020 1262
rect 12084 1260 12090 1324
rect 17718 1260 17724 1324
rect 17788 1322 17794 1324
rect 20529 1322 20595 1325
rect 17788 1320 20595 1322
rect 17788 1264 20534 1320
rect 20590 1264 20595 1320
rect 17788 1262 20595 1264
rect 17788 1260 17794 1262
rect 20529 1259 20595 1262
rect 2773 1186 2839 1189
rect 13670 1186 13676 1188
rect 2730 1184 13676 1186
rect 2730 1128 2778 1184
rect 2834 1128 13676 1184
rect 2730 1126 13676 1128
rect 2730 1123 2839 1126
rect 13670 1124 13676 1126
rect 13740 1124 13746 1188
rect 0 1050 800 1080
rect 2730 1050 2790 1123
rect 0 990 2790 1050
rect 0 960 800 990
rect 4102 988 4108 1052
rect 4172 1050 4178 1052
rect 15009 1050 15075 1053
rect 4172 1048 15075 1050
rect 4172 992 15014 1048
rect 15070 992 15075 1048
rect 4172 990 15075 992
rect 4172 988 4178 990
rect 15009 987 15075 990
rect 20529 1050 20595 1053
rect 22200 1050 23000 1080
rect 20529 1048 23000 1050
rect 20529 992 20534 1048
rect 20590 992 23000 1048
rect 20529 990 23000 992
rect 20529 987 20595 990
rect 22200 960 23000 990
rect 0 642 800 672
rect 2998 642 3004 644
rect 0 582 3004 642
rect 0 552 800 582
rect 2998 580 3004 582
rect 3068 580 3074 644
rect 21633 642 21699 645
rect 22200 642 23000 672
rect 21633 640 23000 642
rect 21633 584 21638 640
rect 21694 584 23000 640
rect 21633 582 23000 584
rect 21633 579 21699 582
rect 22200 552 23000 582
rect 3877 98 3943 101
rect 12750 98 12756 100
rect 3877 96 12756 98
rect 3877 40 3882 96
rect 3938 40 12756 96
rect 3877 38 12756 40
rect 3877 35 3943 38
rect 12750 36 12756 38
rect 12820 36 12826 100
<< via3 >>
rect 14596 22476 14660 22540
rect 1164 21660 1228 21724
rect 12940 21660 13004 21724
rect 1716 21524 1780 21588
rect 13308 21252 13372 21316
rect 14412 21116 14476 21180
rect 7420 20980 7484 21044
rect 7236 20844 7300 20908
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 10180 20300 10244 20364
rect 11100 20360 11164 20364
rect 11100 20304 11114 20360
rect 11114 20304 11164 20360
rect 11100 20300 11164 20304
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 10548 19756 10612 19820
rect 5948 19620 6012 19684
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3004 19544 3068 19548
rect 3004 19488 3018 19544
rect 3018 19488 3068 19544
rect 3004 19484 3068 19488
rect 9812 19484 9876 19548
rect 19564 19348 19628 19412
rect 3372 19212 3436 19276
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 3924 18864 3988 18868
rect 3924 18808 3938 18864
rect 3938 18808 3988 18864
rect 3924 18804 3988 18808
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 5028 18260 5092 18324
rect 9260 17988 9324 18052
rect 12020 17988 12084 18052
rect 20484 17988 20548 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 5212 17852 5276 17916
rect 17172 17852 17236 17916
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 7604 17232 7668 17236
rect 7604 17176 7654 17232
rect 7654 17176 7668 17232
rect 7604 17172 7668 17176
rect 6684 16900 6748 16964
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 1900 16628 1964 16692
rect 19748 16628 19812 16692
rect 20300 16688 20364 16692
rect 20300 16632 20350 16688
rect 20350 16632 20364 16688
rect 20300 16628 20364 16632
rect 980 16356 1044 16420
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 15700 16552 15764 16556
rect 15700 16496 15750 16552
rect 15750 16496 15764 16552
rect 15700 16492 15764 16496
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 17540 15948 17604 16012
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 4844 15676 4908 15740
rect 3924 15404 3988 15468
rect 19564 15404 19628 15468
rect 3004 15328 3068 15332
rect 3004 15272 3054 15328
rect 3054 15272 3068 15328
rect 3004 15268 3068 15272
rect 4292 15268 4356 15332
rect 8340 15328 8404 15332
rect 8340 15272 8354 15328
rect 8354 15272 8404 15328
rect 8340 15268 8404 15272
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 5948 15192 6012 15196
rect 5948 15136 5962 15192
rect 5962 15136 6012 15192
rect 5948 15132 6012 15136
rect 7052 15132 7116 15196
rect 11836 15268 11900 15332
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 8156 14648 8220 14652
rect 8156 14592 8206 14648
rect 8206 14592 8220 14648
rect 8156 14588 8220 14592
rect 3372 14452 3436 14516
rect 7604 14452 7668 14516
rect 2268 14180 2332 14244
rect 14412 14240 14476 14244
rect 14412 14184 14426 14240
rect 14426 14184 14476 14240
rect 14412 14180 14476 14184
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 14412 14044 14476 14108
rect 19564 14104 19628 14108
rect 19564 14048 19578 14104
rect 19578 14048 19628 14104
rect 19564 14044 19628 14048
rect 9444 13772 9508 13836
rect 5580 13636 5644 13700
rect 11100 13772 11164 13836
rect 12204 13832 12268 13836
rect 12204 13776 12254 13832
rect 12254 13776 12268 13832
rect 12204 13772 12268 13776
rect 13492 13832 13556 13836
rect 13492 13776 13506 13832
rect 13506 13776 13556 13832
rect 13492 13772 13556 13776
rect 14964 13772 15028 13836
rect 19932 13772 19996 13836
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 1348 13500 1412 13564
rect 4108 13500 4172 13564
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 21036 13500 21100 13564
rect 2820 13228 2884 13292
rect 12572 13364 12636 13428
rect 10180 13228 10244 13292
rect 16068 13228 16132 13292
rect 19564 13228 19628 13292
rect 7788 13092 7852 13156
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 3188 12956 3252 13020
rect 4108 12956 4172 13020
rect 6868 12956 6932 13020
rect 10364 12956 10428 13020
rect 12940 12956 13004 13020
rect 13676 12880 13740 12884
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 13676 12824 13690 12880
rect 13690 12824 13740 12880
rect 13676 12820 13740 12824
rect 16988 12820 17052 12884
rect 980 12684 1044 12748
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 7604 12684 7668 12748
rect 17724 12548 17788 12612
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 9628 12412 9692 12476
rect 10548 12472 10612 12476
rect 10548 12416 10598 12472
rect 10598 12416 10612 12472
rect 10548 12412 10612 12416
rect 12020 12472 12084 12476
rect 12020 12416 12034 12472
rect 12034 12416 12084 12472
rect 7236 12276 7300 12340
rect 7420 12276 7484 12340
rect 7972 12276 8036 12340
rect 9996 12276 10060 12340
rect 12020 12412 12084 12416
rect 12940 12276 13004 12340
rect 15884 12276 15948 12340
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 7052 11928 7116 11932
rect 7052 11872 7066 11928
rect 7066 11872 7116 11928
rect 7052 11868 7116 11872
rect 7236 11868 7300 11932
rect 8524 11928 8588 11932
rect 8524 11872 8574 11928
rect 8574 11872 8588 11928
rect 8524 11868 8588 11872
rect 9260 11868 9324 11932
rect 10548 11868 10612 11932
rect 14412 12004 14476 12068
rect 14780 12004 14844 12068
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 14412 11868 14476 11932
rect 15332 11868 15396 11932
rect 12020 11732 12084 11796
rect 12388 11732 12452 11796
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 1716 11384 1780 11388
rect 1716 11328 1730 11384
rect 1730 11328 1780 11384
rect 1716 11324 1780 11328
rect 5580 11596 5644 11660
rect 14596 11596 14660 11660
rect 17172 11596 17236 11660
rect 18644 11596 18708 11660
rect 4476 11460 4540 11524
rect 7972 11460 8036 11524
rect 12020 11460 12084 11524
rect 15332 11460 15396 11524
rect 17172 11460 17236 11524
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6684 11324 6748 11388
rect 7972 11324 8036 11388
rect 9628 11324 9692 11388
rect 12940 11324 13004 11388
rect 13308 11384 13372 11388
rect 13308 11328 13358 11384
rect 13358 11328 13372 11384
rect 13308 11324 13372 11328
rect 3924 11188 3988 11252
rect 4108 11188 4172 11252
rect 8340 11188 8404 11252
rect 10732 11188 10796 11252
rect 12388 11188 12452 11252
rect 15148 11188 15212 11252
rect 19748 11188 19812 11252
rect 5396 11052 5460 11116
rect 12756 11052 12820 11116
rect 19932 11052 19996 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 8340 10916 8404 10980
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 5948 10704 6012 10708
rect 5948 10648 5998 10704
rect 5998 10648 6012 10704
rect 5948 10644 6012 10648
rect 7420 10644 7484 10708
rect 7788 10644 7852 10708
rect 14596 10780 14660 10844
rect 21036 10780 21100 10844
rect 5580 10372 5644 10436
rect 7052 10432 7116 10436
rect 7052 10376 7066 10432
rect 7066 10376 7116 10432
rect 7052 10372 7116 10376
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 7788 10296 7852 10300
rect 7788 10240 7838 10296
rect 7838 10240 7852 10296
rect 7788 10236 7852 10240
rect 4844 10100 4908 10164
rect 7236 10100 7300 10164
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 10364 10236 10428 10300
rect 17540 10508 17604 10572
rect 17540 10372 17604 10436
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 18828 10236 18892 10300
rect 20116 10100 20180 10164
rect 5580 9888 5644 9892
rect 5580 9832 5594 9888
rect 5594 9832 5644 9888
rect 5580 9828 5644 9832
rect 7052 9828 7116 9892
rect 9260 9828 9324 9892
rect 11100 9964 11164 10028
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 12572 9828 12636 9892
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 10180 9752 10244 9756
rect 10180 9696 10194 9752
rect 10194 9696 10244 9752
rect 10180 9692 10244 9696
rect 12572 9692 12636 9756
rect 3004 9556 3068 9620
rect 5212 9556 5276 9620
rect 6868 9420 6932 9484
rect 4660 9284 4724 9348
rect 9996 9284 10060 9348
rect 14780 9284 14844 9348
rect 17356 9284 17420 9348
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 9444 9148 9508 9212
rect 5212 9012 5276 9076
rect 9812 9012 9876 9076
rect 16988 9012 17052 9076
rect 5028 8876 5092 8940
rect 5948 8740 6012 8804
rect 6684 8740 6748 8804
rect 1900 8604 1964 8668
rect 2452 8664 2516 8668
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 2452 8608 2502 8664
rect 2502 8608 2516 8664
rect 2452 8604 2516 8608
rect 1716 8468 1780 8532
rect 8156 8604 8220 8668
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 7420 8528 7484 8532
rect 7420 8472 7470 8528
rect 7470 8472 7484 8528
rect 7420 8468 7484 8472
rect 17908 8332 17972 8396
rect 19932 8196 19996 8260
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 5396 8060 5460 8124
rect 10364 7924 10428 7988
rect 15332 7924 15396 7988
rect 4108 7788 4172 7852
rect 5212 7788 5276 7852
rect 5948 7788 6012 7852
rect 4292 7652 4356 7716
rect 5028 7652 5092 7716
rect 7236 7652 7300 7716
rect 10548 7652 10612 7716
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 5580 7516 5644 7580
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 17540 7380 17604 7444
rect 6684 7108 6748 7172
rect 7420 7168 7484 7172
rect 7420 7112 7434 7168
rect 7434 7112 7484 7168
rect 7420 7108 7484 7112
rect 9996 7168 10060 7172
rect 9996 7112 10046 7168
rect 10046 7112 10060 7168
rect 9996 7108 10060 7112
rect 17172 7108 17236 7172
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 4844 6972 4908 7036
rect 8524 6972 8588 7036
rect 9444 6972 9508 7036
rect 1716 6836 1780 6900
rect 3924 6836 3988 6900
rect 15884 6836 15948 6900
rect 18644 6836 18708 6900
rect 2636 6624 2700 6628
rect 2636 6568 2686 6624
rect 2686 6568 2700 6624
rect 2636 6564 2700 6568
rect 4660 6624 4724 6628
rect 4660 6568 4710 6624
rect 4710 6568 4724 6624
rect 4660 6564 4724 6568
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 2268 6428 2332 6492
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 4108 6292 4172 6356
rect 14964 6156 15028 6220
rect 4476 6020 4540 6084
rect 7052 6020 7116 6084
rect 7236 6020 7300 6084
rect 11836 6020 11900 6084
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 2820 5884 2884 5948
rect 8340 5884 8404 5948
rect 11836 5884 11900 5948
rect 15700 5884 15764 5948
rect 16068 5808 16132 5812
rect 16068 5752 16118 5808
rect 16118 5752 16132 5808
rect 16068 5748 16132 5752
rect 3372 5612 3436 5676
rect 3924 5612 3988 5676
rect 3188 5476 3252 5540
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 980 5204 1044 5268
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 7604 5400 7668 5404
rect 7604 5344 7618 5400
rect 7618 5344 7668 5400
rect 7604 5340 7668 5344
rect 3188 5068 3252 5132
rect 2452 4932 2516 4996
rect 4844 4932 4908 4996
rect 5580 5068 5644 5132
rect 8156 5204 8220 5268
rect 12020 5476 12084 5540
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 15148 5400 15212 5404
rect 15148 5344 15198 5400
rect 15198 5344 15212 5400
rect 15148 5340 15212 5344
rect 7604 4932 7668 4996
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 980 4660 1044 4724
rect 8156 4796 8220 4860
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 12940 4660 13004 4724
rect 6684 4524 6748 4588
rect 13492 4524 13556 4588
rect 4108 4388 4172 4452
rect 5396 4388 5460 4452
rect 17540 4388 17604 4452
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 4108 4252 4172 4316
rect 14412 4116 14476 4180
rect 5028 3980 5092 4044
rect 5948 3980 6012 4044
rect 6684 3980 6748 4044
rect 12572 3980 12636 4044
rect 2636 3844 2700 3908
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 980 3708 1044 3772
rect 4476 3572 4540 3636
rect 4660 3436 4724 3500
rect 7788 3844 7852 3908
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 7972 3708 8036 3772
rect 9260 3708 9324 3772
rect 20300 4040 20364 4044
rect 20300 3984 20314 4040
rect 20314 3984 20364 4040
rect 20300 3980 20364 3984
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 18828 3844 18892 3908
rect 20484 3844 20548 3908
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 19748 3708 19812 3772
rect 11836 3572 11900 3636
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 3372 2952 3436 2956
rect 3372 2896 3386 2952
rect 3386 2896 3436 2952
rect 3372 2892 3436 2896
rect 5212 2892 5276 2956
rect 7972 3436 8036 3500
rect 9260 3436 9324 3500
rect 15700 3300 15764 3364
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 9996 3164 10060 3228
rect 17908 3028 17972 3092
rect 10732 2892 10796 2956
rect 14596 2892 14660 2956
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 1164 2484 1228 2548
rect 5580 2620 5644 2684
rect 6868 2620 6932 2684
rect 10180 2620 10244 2684
rect 1348 2212 1412 2276
rect 7236 2484 7300 2548
rect 7604 2544 7668 2548
rect 7604 2488 7618 2544
rect 7618 2488 7668 2544
rect 7604 2484 7668 2488
rect 11100 2484 11164 2548
rect 7420 2348 7484 2412
rect 12204 2348 12268 2412
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
rect 17356 1940 17420 2004
rect 10364 1668 10428 1732
rect 9444 1396 9508 1460
rect 5396 1260 5460 1324
rect 12020 1260 12084 1324
rect 17724 1260 17788 1324
rect 13676 1124 13740 1188
rect 4108 988 4172 1052
rect 3004 580 3068 644
rect 12756 36 12820 100
<< metal4 >>
rect 14595 22540 14661 22541
rect 14595 22476 14596 22540
rect 14660 22476 14661 22540
rect 14595 22475 14661 22476
rect 1163 21724 1229 21725
rect 1163 21660 1164 21724
rect 1228 21660 1229 21724
rect 1163 21659 1229 21660
rect 12939 21724 13005 21725
rect 12939 21660 12940 21724
rect 13004 21660 13005 21724
rect 12939 21659 13005 21660
rect 979 16420 1045 16421
rect 979 16356 980 16420
rect 1044 16356 1045 16420
rect 979 16355 1045 16356
rect 982 13290 1042 16355
rect 614 13230 1042 13290
rect 614 5130 674 13230
rect 979 12748 1045 12749
rect 979 12684 980 12748
rect 1044 12684 1045 12748
rect 979 12683 1045 12684
rect 982 5269 1042 12683
rect 979 5268 1045 5269
rect 979 5204 980 5268
rect 1044 5204 1045 5268
rect 979 5203 1045 5204
rect 614 5070 1042 5130
rect 982 4725 1042 5070
rect 979 4724 1045 4725
rect 979 4660 980 4724
rect 1044 4660 1045 4724
rect 979 4659 1045 4660
rect 982 3773 1042 4659
rect 979 3772 1045 3773
rect 979 3708 980 3772
rect 1044 3708 1045 3772
rect 979 3707 1045 3708
rect 1166 2549 1226 21659
rect 1715 21588 1781 21589
rect 1715 21524 1716 21588
rect 1780 21524 1781 21588
rect 1715 21523 1781 21524
rect 1347 13564 1413 13565
rect 1347 13500 1348 13564
rect 1412 13500 1413 13564
rect 1347 13499 1413 13500
rect 1163 2548 1229 2549
rect 1163 2484 1164 2548
rect 1228 2484 1229 2548
rect 1163 2483 1229 2484
rect 1350 2277 1410 13499
rect 1718 11389 1778 21523
rect 7419 21044 7485 21045
rect 7419 20980 7420 21044
rect 7484 20980 7485 21044
rect 7419 20979 7485 20980
rect 7235 20908 7301 20909
rect 7235 20844 7236 20908
rect 7300 20844 7301 20908
rect 7235 20843 7301 20844
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3003 19548 3069 19549
rect 3003 19484 3004 19548
rect 3068 19484 3069 19548
rect 3003 19483 3069 19484
rect 1899 16692 1965 16693
rect 1899 16628 1900 16692
rect 1964 16628 1965 16692
rect 1899 16627 1965 16628
rect 1715 11388 1781 11389
rect 1715 11324 1716 11388
rect 1780 11324 1781 11388
rect 1715 11323 1781 11324
rect 1902 8669 1962 16627
rect 3006 15333 3066 19483
rect 3371 19276 3437 19277
rect 3371 19212 3372 19276
rect 3436 19212 3437 19276
rect 3371 19211 3437 19212
rect 3003 15332 3069 15333
rect 3003 15268 3004 15332
rect 3068 15268 3069 15332
rect 3003 15267 3069 15268
rect 3374 14517 3434 19211
rect 3543 19072 3863 20096
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 5947 19684 6013 19685
rect 5947 19620 5948 19684
rect 6012 19620 6013 19684
rect 5947 19619 6013 19620
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3923 18868 3989 18869
rect 3923 18804 3924 18868
rect 3988 18804 3989 18868
rect 3923 18803 3989 18804
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3926 15469 3986 18803
rect 5027 18324 5093 18325
rect 5027 18260 5028 18324
rect 5092 18260 5093 18324
rect 5027 18259 5093 18260
rect 4843 15740 4909 15741
rect 4843 15676 4844 15740
rect 4908 15676 4909 15740
rect 4843 15675 4909 15676
rect 3923 15468 3989 15469
rect 3923 15404 3924 15468
rect 3988 15404 3989 15468
rect 3923 15403 3989 15404
rect 4291 15332 4357 15333
rect 4291 15268 4292 15332
rect 4356 15268 4357 15332
rect 4291 15267 4357 15268
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3371 14516 3437 14517
rect 3371 14452 3372 14516
rect 3436 14452 3437 14516
rect 3371 14451 3437 14452
rect 2267 14244 2333 14245
rect 2267 14180 2268 14244
rect 2332 14180 2333 14244
rect 2267 14179 2333 14180
rect 1899 8668 1965 8669
rect 1899 8604 1900 8668
rect 1964 8604 1965 8668
rect 1899 8603 1965 8604
rect 1715 8532 1781 8533
rect 1715 8468 1716 8532
rect 1780 8468 1781 8532
rect 1715 8467 1781 8468
rect 1718 6901 1778 8467
rect 1715 6900 1781 6901
rect 1715 6836 1716 6900
rect 1780 6836 1781 6900
rect 1715 6835 1781 6836
rect 2270 6493 2330 14179
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 2819 13292 2885 13293
rect 2819 13228 2820 13292
rect 2884 13228 2885 13292
rect 2819 13227 2885 13228
rect 2451 8668 2517 8669
rect 2451 8604 2452 8668
rect 2516 8604 2517 8668
rect 2451 8603 2517 8604
rect 2267 6492 2333 6493
rect 2267 6428 2268 6492
rect 2332 6428 2333 6492
rect 2267 6427 2333 6428
rect 2454 4997 2514 8603
rect 2635 6628 2701 6629
rect 2635 6564 2636 6628
rect 2700 6564 2701 6628
rect 2635 6563 2701 6564
rect 2451 4996 2517 4997
rect 2451 4932 2452 4996
rect 2516 4932 2517 4996
rect 2451 4931 2517 4932
rect 2638 3909 2698 6563
rect 2822 5949 2882 13227
rect 3187 13020 3253 13021
rect 3187 12956 3188 13020
rect 3252 12956 3253 13020
rect 3187 12955 3253 12956
rect 3003 9620 3069 9621
rect 3003 9556 3004 9620
rect 3068 9556 3069 9620
rect 3003 9555 3069 9556
rect 2819 5948 2885 5949
rect 2819 5884 2820 5948
rect 2884 5884 2885 5948
rect 2819 5883 2885 5884
rect 2635 3908 2701 3909
rect 2635 3844 2636 3908
rect 2700 3844 2701 3908
rect 2635 3843 2701 3844
rect 1347 2276 1413 2277
rect 1347 2212 1348 2276
rect 1412 2212 1413 2276
rect 1347 2211 1413 2212
rect 3006 645 3066 9555
rect 3190 5541 3250 12955
rect 3543 12544 3863 13568
rect 4107 13564 4173 13565
rect 4107 13500 4108 13564
rect 4172 13500 4173 13564
rect 4107 13499 4173 13500
rect 4110 13021 4170 13499
rect 4107 13020 4173 13021
rect 4107 12956 4108 13020
rect 4172 12956 4173 13020
rect 4107 12955 4173 12956
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3923 11252 3989 11253
rect 3923 11188 3924 11252
rect 3988 11188 3989 11252
rect 3923 11187 3989 11188
rect 4107 11252 4173 11253
rect 4107 11188 4108 11252
rect 4172 11188 4173 11252
rect 4107 11187 4173 11188
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3926 6901 3986 11187
rect 4110 7853 4170 11187
rect 4107 7852 4173 7853
rect 4107 7788 4108 7852
rect 4172 7788 4173 7852
rect 4107 7787 4173 7788
rect 4294 7717 4354 15267
rect 4475 11524 4541 11525
rect 4475 11460 4476 11524
rect 4540 11460 4541 11524
rect 4475 11459 4541 11460
rect 4291 7716 4357 7717
rect 4291 7652 4292 7716
rect 4356 7652 4357 7716
rect 4291 7651 4357 7652
rect 4478 7170 4538 11459
rect 4846 10165 4906 15675
rect 4843 10164 4909 10165
rect 4843 10100 4844 10164
rect 4908 10100 4909 10164
rect 4843 10099 4909 10100
rect 4659 9348 4725 9349
rect 4659 9284 4660 9348
rect 4724 9284 4725 9348
rect 4659 9283 4725 9284
rect 4110 7110 4538 7170
rect 3923 6900 3989 6901
rect 3923 6836 3924 6900
rect 3988 6836 3989 6900
rect 3923 6835 3989 6836
rect 4110 6490 4170 7110
rect 4662 6629 4722 9283
rect 5030 8941 5090 18259
rect 5211 17916 5277 17917
rect 5211 17852 5212 17916
rect 5276 17852 5277 17916
rect 5211 17851 5277 17852
rect 5214 9621 5274 17851
rect 5950 15197 6010 19619
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6683 16964 6749 16965
rect 6683 16900 6684 16964
rect 6748 16900 6749 16964
rect 6683 16899 6749 16900
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 5947 15196 6013 15197
rect 5947 15132 5948 15196
rect 6012 15132 6013 15196
rect 5947 15131 6013 15132
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 5579 13700 5645 13701
rect 5579 13636 5580 13700
rect 5644 13636 5645 13700
rect 5579 13635 5645 13636
rect 5582 12450 5642 13635
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 5582 12390 5826 12450
rect 5579 11660 5645 11661
rect 5579 11596 5580 11660
rect 5644 11596 5645 11660
rect 5579 11595 5645 11596
rect 5395 11116 5461 11117
rect 5395 11052 5396 11116
rect 5460 11052 5461 11116
rect 5395 11051 5461 11052
rect 5211 9620 5277 9621
rect 5211 9556 5212 9620
rect 5276 9556 5277 9620
rect 5211 9555 5277 9556
rect 5214 9077 5274 9555
rect 5211 9076 5277 9077
rect 5211 9012 5212 9076
rect 5276 9012 5277 9076
rect 5211 9011 5277 9012
rect 5027 8940 5093 8941
rect 5027 8876 5028 8940
rect 5092 8876 5093 8940
rect 5027 8875 5093 8876
rect 5398 8125 5458 11051
rect 5582 10437 5642 11595
rect 5579 10436 5645 10437
rect 5579 10372 5580 10436
rect 5644 10372 5645 10436
rect 5579 10371 5645 10372
rect 5579 9892 5645 9893
rect 5579 9828 5580 9892
rect 5644 9828 5645 9892
rect 5579 9827 5645 9828
rect 5395 8124 5461 8125
rect 5395 8060 5396 8124
rect 5460 8060 5461 8124
rect 5395 8059 5461 8060
rect 5211 7852 5277 7853
rect 5211 7788 5212 7852
rect 5276 7788 5277 7852
rect 5211 7787 5277 7788
rect 5027 7716 5093 7717
rect 5027 7652 5028 7716
rect 5092 7652 5093 7716
rect 5027 7651 5093 7652
rect 4843 7036 4909 7037
rect 4843 6972 4844 7036
rect 4908 6972 4909 7036
rect 4843 6971 4909 6972
rect 4659 6628 4725 6629
rect 4659 6564 4660 6628
rect 4724 6564 4725 6628
rect 4659 6563 4725 6564
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3371 5676 3437 5677
rect 3371 5612 3372 5676
rect 3436 5612 3437 5676
rect 3371 5611 3437 5612
rect 3187 5540 3253 5541
rect 3187 5476 3188 5540
rect 3252 5476 3253 5540
rect 3187 5475 3253 5476
rect 3190 5133 3250 5475
rect 3187 5132 3253 5133
rect 3187 5068 3188 5132
rect 3252 5068 3253 5132
rect 3187 5067 3253 5068
rect 3374 2957 3434 5611
rect 3543 4928 3863 5952
rect 3926 6430 4170 6490
rect 3926 5677 3986 6430
rect 4107 6356 4173 6357
rect 4107 6292 4108 6356
rect 4172 6292 4173 6356
rect 4107 6291 4173 6292
rect 3923 5676 3989 5677
rect 3923 5612 3924 5676
rect 3988 5612 3989 5676
rect 3923 5611 3989 5612
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 4110 4453 4170 6291
rect 4475 6084 4541 6085
rect 4475 6020 4476 6084
rect 4540 6020 4541 6084
rect 4475 6019 4541 6020
rect 4107 4452 4173 4453
rect 4107 4388 4108 4452
rect 4172 4388 4173 4452
rect 4107 4387 4173 4388
rect 4107 4316 4173 4317
rect 4107 4252 4108 4316
rect 4172 4252 4173 4316
rect 4107 4251 4173 4252
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3371 2956 3437 2957
rect 3371 2892 3372 2956
rect 3436 2892 3437 2956
rect 3371 2891 3437 2892
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 4110 1053 4170 4251
rect 4478 3637 4538 6019
rect 4475 3636 4541 3637
rect 4475 3572 4476 3636
rect 4540 3572 4541 3636
rect 4475 3571 4541 3572
rect 4662 3501 4722 6563
rect 4846 4997 4906 6971
rect 4843 4996 4909 4997
rect 4843 4932 4844 4996
rect 4908 4932 4909 4996
rect 4843 4931 4909 4932
rect 5030 4045 5090 7651
rect 5027 4044 5093 4045
rect 5027 3980 5028 4044
rect 5092 3980 5093 4044
rect 5027 3979 5093 3980
rect 4659 3500 4725 3501
rect 4659 3436 4660 3500
rect 4724 3436 4725 3500
rect 4659 3435 4725 3436
rect 5214 2957 5274 7787
rect 5582 7581 5642 9827
rect 5579 7580 5645 7581
rect 5579 7516 5580 7580
rect 5644 7516 5645 7580
rect 5579 7515 5645 7516
rect 5766 6490 5826 12390
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6686 11389 6746 16899
rect 7051 15196 7117 15197
rect 7051 15132 7052 15196
rect 7116 15132 7117 15196
rect 7051 15131 7117 15132
rect 6867 13020 6933 13021
rect 6867 12956 6868 13020
rect 6932 12956 6933 13020
rect 6867 12955 6933 12956
rect 6683 11388 6749 11389
rect 6683 11324 6684 11388
rect 6748 11324 6749 11388
rect 6683 11323 6749 11324
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 5947 10708 6013 10709
rect 5947 10644 5948 10708
rect 6012 10644 6013 10708
rect 5947 10643 6013 10644
rect 5950 8805 6010 10643
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 5947 8804 6013 8805
rect 5947 8740 5948 8804
rect 6012 8740 6013 8804
rect 5947 8739 6013 8740
rect 6142 8736 6462 9760
rect 6870 9485 6930 12955
rect 7054 12066 7114 15131
rect 7238 12341 7298 20843
rect 7422 12341 7482 20979
rect 8741 20160 9061 20720
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 10179 20364 10245 20365
rect 10179 20300 10180 20364
rect 10244 20300 10245 20364
rect 10179 20299 10245 20300
rect 11099 20364 11165 20365
rect 11099 20300 11100 20364
rect 11164 20300 11165 20364
rect 11099 20299 11165 20300
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 9811 19548 9877 19549
rect 9811 19484 9812 19548
rect 9876 19484 9877 19548
rect 9811 19483 9877 19484
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 9259 18052 9325 18053
rect 9259 17988 9260 18052
rect 9324 17988 9325 18052
rect 9259 17987 9325 17988
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 7603 17236 7669 17237
rect 7603 17172 7604 17236
rect 7668 17172 7669 17236
rect 7603 17171 7669 17172
rect 7606 14517 7666 17171
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8339 15332 8405 15333
rect 8339 15268 8340 15332
rect 8404 15268 8405 15332
rect 8339 15267 8405 15268
rect 8155 14652 8221 14653
rect 8155 14588 8156 14652
rect 8220 14588 8221 14652
rect 8155 14587 8221 14588
rect 7603 14516 7669 14517
rect 7603 14452 7604 14516
rect 7668 14452 7669 14516
rect 7603 14451 7669 14452
rect 7787 13156 7853 13157
rect 7787 13092 7788 13156
rect 7852 13092 7853 13156
rect 7787 13091 7853 13092
rect 7603 12748 7669 12749
rect 7603 12684 7604 12748
rect 7668 12684 7669 12748
rect 7603 12683 7669 12684
rect 7235 12340 7301 12341
rect 7235 12276 7236 12340
rect 7300 12276 7301 12340
rect 7235 12275 7301 12276
rect 7419 12340 7485 12341
rect 7419 12276 7420 12340
rect 7484 12276 7485 12340
rect 7419 12275 7485 12276
rect 7054 12006 7482 12066
rect 7051 11932 7117 11933
rect 7051 11868 7052 11932
rect 7116 11868 7117 11932
rect 7051 11867 7117 11868
rect 7235 11932 7301 11933
rect 7235 11868 7236 11932
rect 7300 11868 7301 11932
rect 7235 11867 7301 11868
rect 7054 10437 7114 11867
rect 7051 10436 7117 10437
rect 7051 10372 7052 10436
rect 7116 10372 7117 10436
rect 7238 10434 7298 11867
rect 7422 10709 7482 12006
rect 7419 10708 7485 10709
rect 7419 10644 7420 10708
rect 7484 10644 7485 10708
rect 7419 10643 7485 10644
rect 7606 10570 7666 12683
rect 7790 10709 7850 13091
rect 7971 12340 8037 12341
rect 7971 12276 7972 12340
rect 8036 12276 8037 12340
rect 7971 12275 8037 12276
rect 7974 11525 8034 12275
rect 7971 11524 8037 11525
rect 7971 11460 7972 11524
rect 8036 11460 8037 11524
rect 7971 11459 8037 11460
rect 7971 11388 8037 11389
rect 7971 11324 7972 11388
rect 8036 11324 8037 11388
rect 7971 11323 8037 11324
rect 7787 10708 7853 10709
rect 7787 10644 7788 10708
rect 7852 10644 7853 10708
rect 7787 10643 7853 10644
rect 7606 10510 7712 10570
rect 7238 10374 7482 10434
rect 7051 10371 7117 10372
rect 7235 10164 7301 10165
rect 7235 10100 7236 10164
rect 7300 10100 7301 10164
rect 7235 10099 7301 10100
rect 7051 9892 7117 9893
rect 7051 9828 7052 9892
rect 7116 9828 7117 9892
rect 7051 9827 7117 9828
rect 6867 9484 6933 9485
rect 6867 9420 6868 9484
rect 6932 9420 6933 9484
rect 6867 9419 6933 9420
rect 6683 8804 6749 8805
rect 6683 8740 6684 8804
rect 6748 8740 6749 8804
rect 6683 8739 6749 8740
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 5947 7852 6013 7853
rect 5947 7788 5948 7852
rect 6012 7788 6013 7852
rect 5947 7787 6013 7788
rect 5582 6430 5826 6490
rect 5582 5133 5642 6430
rect 5579 5132 5645 5133
rect 5579 5068 5580 5132
rect 5644 5068 5645 5132
rect 5579 5067 5645 5068
rect 5395 4452 5461 4453
rect 5395 4388 5396 4452
rect 5460 4388 5461 4452
rect 5395 4387 5461 4388
rect 5211 2956 5277 2957
rect 5211 2892 5212 2956
rect 5276 2892 5277 2956
rect 5211 2891 5277 2892
rect 5398 1325 5458 4387
rect 5582 2685 5642 5067
rect 5950 4045 6010 7787
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6686 7173 6746 8739
rect 6683 7172 6749 7173
rect 6683 7108 6684 7172
rect 6748 7108 6749 7172
rect 6683 7107 6749 7108
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6683 4588 6749 4589
rect 6683 4524 6684 4588
rect 6748 4524 6749 4588
rect 6683 4523 6749 4524
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 5947 4044 6013 4045
rect 5947 3980 5948 4044
rect 6012 3980 6013 4044
rect 5947 3979 6013 3980
rect 6142 3296 6462 4320
rect 6686 4045 6746 4523
rect 6683 4044 6749 4045
rect 6683 3980 6684 4044
rect 6748 3980 6749 4044
rect 6683 3979 6749 3980
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 5579 2684 5645 2685
rect 5579 2620 5580 2684
rect 5644 2620 5645 2684
rect 5579 2619 5645 2620
rect 6142 2208 6462 3232
rect 6870 2685 6930 9419
rect 7054 6085 7114 9827
rect 7238 7717 7298 10099
rect 7422 8533 7482 10374
rect 7652 10298 7712 10510
rect 7606 10238 7712 10298
rect 7787 10300 7853 10301
rect 7419 8532 7485 8533
rect 7419 8468 7420 8532
rect 7484 8468 7485 8532
rect 7419 8467 7485 8468
rect 7235 7716 7301 7717
rect 7235 7652 7236 7716
rect 7300 7652 7301 7716
rect 7235 7651 7301 7652
rect 7419 7172 7485 7173
rect 7419 7108 7420 7172
rect 7484 7108 7485 7172
rect 7419 7107 7485 7108
rect 7051 6084 7117 6085
rect 7051 6020 7052 6084
rect 7116 6020 7117 6084
rect 7051 6019 7117 6020
rect 7235 6084 7301 6085
rect 7235 6020 7236 6084
rect 7300 6020 7301 6084
rect 7235 6019 7301 6020
rect 6867 2684 6933 2685
rect 6867 2620 6868 2684
rect 6932 2620 6933 2684
rect 6867 2619 6933 2620
rect 7238 2549 7298 6019
rect 7235 2548 7301 2549
rect 7235 2484 7236 2548
rect 7300 2484 7301 2548
rect 7235 2483 7301 2484
rect 7422 2413 7482 7107
rect 7606 5405 7666 10238
rect 7787 10236 7788 10300
rect 7852 10236 7853 10300
rect 7787 10235 7853 10236
rect 7603 5404 7669 5405
rect 7603 5340 7604 5404
rect 7668 5340 7669 5404
rect 7603 5339 7669 5340
rect 7603 4996 7669 4997
rect 7603 4932 7604 4996
rect 7668 4932 7669 4996
rect 7603 4931 7669 4932
rect 7606 2549 7666 4931
rect 7790 3909 7850 10235
rect 7787 3908 7853 3909
rect 7787 3844 7788 3908
rect 7852 3844 7853 3908
rect 7787 3843 7853 3844
rect 7974 3773 8034 11323
rect 8158 8669 8218 14587
rect 8342 11253 8402 15267
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8523 11932 8589 11933
rect 8523 11868 8524 11932
rect 8588 11868 8589 11932
rect 8523 11867 8589 11868
rect 8339 11252 8405 11253
rect 8339 11188 8340 11252
rect 8404 11188 8405 11252
rect 8339 11187 8405 11188
rect 8339 10980 8405 10981
rect 8339 10916 8340 10980
rect 8404 10916 8405 10980
rect 8339 10915 8405 10916
rect 8155 8668 8221 8669
rect 8155 8604 8156 8668
rect 8220 8604 8221 8668
rect 8155 8603 8221 8604
rect 8342 5949 8402 10915
rect 8526 7037 8586 11867
rect 8741 11456 9061 12480
rect 9262 11933 9322 17987
rect 9443 13836 9509 13837
rect 9443 13772 9444 13836
rect 9508 13772 9509 13836
rect 9443 13771 9509 13772
rect 9259 11932 9325 11933
rect 9259 11868 9260 11932
rect 9324 11868 9325 11932
rect 9259 11867 9325 11868
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 9262 9893 9322 11867
rect 9259 9892 9325 9893
rect 9259 9828 9260 9892
rect 9324 9828 9325 9892
rect 9259 9827 9325 9828
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 9446 9213 9506 13771
rect 9627 12476 9693 12477
rect 9627 12412 9628 12476
rect 9692 12412 9693 12476
rect 9627 12411 9693 12412
rect 9630 11389 9690 12411
rect 9627 11388 9693 11389
rect 9627 11324 9628 11388
rect 9692 11324 9693 11388
rect 9627 11323 9693 11324
rect 9443 9212 9509 9213
rect 9443 9148 9444 9212
rect 9508 9148 9509 9212
rect 9443 9147 9509 9148
rect 9814 9077 9874 19483
rect 10182 13293 10242 20299
rect 10547 19820 10613 19821
rect 10547 19756 10548 19820
rect 10612 19756 10613 19820
rect 10547 19755 10613 19756
rect 10179 13292 10245 13293
rect 10179 13228 10180 13292
rect 10244 13228 10245 13292
rect 10179 13227 10245 13228
rect 10363 13020 10429 13021
rect 10363 12956 10364 13020
rect 10428 12956 10429 13020
rect 10363 12955 10429 12956
rect 9995 12340 10061 12341
rect 9995 12276 9996 12340
rect 10060 12276 10061 12340
rect 9995 12275 10061 12276
rect 9998 9349 10058 12275
rect 10366 10301 10426 12955
rect 10550 12477 10610 19755
rect 11102 13837 11162 20299
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 12019 18052 12085 18053
rect 12019 17988 12020 18052
rect 12084 17988 12085 18052
rect 12019 17987 12085 17988
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11835 15332 11901 15333
rect 11835 15268 11836 15332
rect 11900 15268 11901 15332
rect 11835 15267 11901 15268
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11099 13836 11165 13837
rect 11099 13772 11100 13836
rect 11164 13772 11165 13836
rect 11099 13771 11165 13772
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 10547 12476 10613 12477
rect 10547 12412 10548 12476
rect 10612 12450 10613 12476
rect 10612 12412 10794 12450
rect 10547 12411 10794 12412
rect 10550 12390 10794 12411
rect 10547 11932 10613 11933
rect 10547 11868 10548 11932
rect 10612 11868 10613 11932
rect 10547 11867 10613 11868
rect 10363 10300 10429 10301
rect 10363 10236 10364 10300
rect 10428 10236 10429 10300
rect 10363 10235 10429 10236
rect 10179 9756 10245 9757
rect 10179 9692 10180 9756
rect 10244 9692 10245 9756
rect 10179 9691 10245 9692
rect 9995 9348 10061 9349
rect 9995 9284 9996 9348
rect 10060 9284 10061 9348
rect 9995 9283 10061 9284
rect 9811 9076 9877 9077
rect 9811 9012 9812 9076
rect 9876 9012 9877 9076
rect 9811 9011 9877 9012
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 9995 7172 10061 7173
rect 9995 7108 9996 7172
rect 10060 7108 10061 7172
rect 9995 7107 10061 7108
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8523 7036 8589 7037
rect 8523 6972 8524 7036
rect 8588 6972 8589 7036
rect 8523 6971 8589 6972
rect 8741 6016 9061 7040
rect 9443 7036 9509 7037
rect 9443 6972 9444 7036
rect 9508 6972 9509 7036
rect 9443 6971 9509 6972
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8339 5948 8405 5949
rect 8339 5884 8340 5948
rect 8404 5884 8405 5948
rect 8339 5883 8405 5884
rect 8155 5268 8221 5269
rect 8155 5204 8156 5268
rect 8220 5204 8221 5268
rect 8155 5203 8221 5204
rect 8158 4861 8218 5203
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8155 4860 8221 4861
rect 8155 4796 8156 4860
rect 8220 4796 8221 4860
rect 8155 4795 8221 4796
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 7971 3772 8037 3773
rect 7971 3708 7972 3772
rect 8036 3708 8037 3772
rect 7971 3707 8037 3708
rect 7974 3501 8034 3707
rect 7971 3500 8037 3501
rect 7971 3436 7972 3500
rect 8036 3436 8037 3500
rect 7971 3435 8037 3436
rect 8741 2752 9061 3776
rect 9259 3772 9325 3773
rect 9259 3708 9260 3772
rect 9324 3708 9325 3772
rect 9259 3707 9325 3708
rect 9262 3501 9322 3707
rect 9259 3500 9325 3501
rect 9259 3436 9260 3500
rect 9324 3436 9325 3500
rect 9259 3435 9325 3436
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 7603 2548 7669 2549
rect 7603 2484 7604 2548
rect 7668 2484 7669 2548
rect 7603 2483 7669 2484
rect 7419 2412 7485 2413
rect 7419 2348 7420 2412
rect 7484 2348 7485 2412
rect 7419 2347 7485 2348
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 2128 9061 2688
rect 9446 1461 9506 6971
rect 9998 3229 10058 7107
rect 9995 3228 10061 3229
rect 9995 3164 9996 3228
rect 10060 3164 10061 3228
rect 9995 3163 10061 3164
rect 10182 2685 10242 9691
rect 10363 7988 10429 7989
rect 10363 7924 10364 7988
rect 10428 7924 10429 7988
rect 10363 7923 10429 7924
rect 10179 2684 10245 2685
rect 10179 2620 10180 2684
rect 10244 2620 10245 2684
rect 10179 2619 10245 2620
rect 10366 1733 10426 7923
rect 10550 7717 10610 11867
rect 10734 11253 10794 12390
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 10731 11252 10797 11253
rect 10731 11188 10732 11252
rect 10796 11188 10797 11252
rect 10731 11187 10797 11188
rect 10547 7716 10613 7717
rect 10547 7652 10548 7716
rect 10612 7652 10613 7716
rect 10547 7651 10613 7652
rect 10734 2957 10794 11187
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11099 10028 11165 10029
rect 11099 9964 11100 10028
rect 11164 9964 11165 10028
rect 11099 9963 11165 9964
rect 10731 2956 10797 2957
rect 10731 2892 10732 2956
rect 10796 2892 10797 2956
rect 10731 2891 10797 2892
rect 11102 2549 11162 9963
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11838 6085 11898 15267
rect 12022 12477 12082 17987
rect 12203 13836 12269 13837
rect 12203 13772 12204 13836
rect 12268 13772 12269 13836
rect 12203 13771 12269 13772
rect 12019 12476 12085 12477
rect 12019 12412 12020 12476
rect 12084 12412 12085 12476
rect 12019 12411 12085 12412
rect 12019 11796 12085 11797
rect 12019 11732 12020 11796
rect 12084 11732 12085 11796
rect 12019 11731 12085 11732
rect 12022 11525 12082 11731
rect 12019 11524 12085 11525
rect 12019 11460 12020 11524
rect 12084 11460 12085 11524
rect 12019 11459 12085 11460
rect 11835 6084 11901 6085
rect 11835 6020 11836 6084
rect 11900 6020 11901 6084
rect 11835 6019 11901 6020
rect 11835 5948 11901 5949
rect 11835 5884 11836 5948
rect 11900 5884 11901 5948
rect 11835 5883 11901 5884
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11838 3637 11898 5883
rect 12022 5541 12082 11459
rect 12019 5540 12085 5541
rect 12019 5476 12020 5540
rect 12084 5476 12085 5540
rect 12019 5475 12085 5476
rect 11835 3636 11901 3637
rect 11835 3572 11836 3636
rect 11900 3572 11901 3636
rect 11835 3571 11901 3572
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11099 2548 11165 2549
rect 11099 2484 11100 2548
rect 11164 2484 11165 2548
rect 11099 2483 11165 2484
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 10363 1732 10429 1733
rect 10363 1668 10364 1732
rect 10428 1668 10429 1732
rect 10363 1667 10429 1668
rect 9443 1460 9509 1461
rect 9443 1396 9444 1460
rect 9508 1396 9509 1460
rect 9443 1395 9509 1396
rect 12022 1325 12082 5475
rect 12206 2413 12266 13771
rect 12571 13428 12637 13429
rect 12571 13364 12572 13428
rect 12636 13364 12637 13428
rect 12571 13363 12637 13364
rect 12387 11796 12453 11797
rect 12387 11732 12388 11796
rect 12452 11732 12453 11796
rect 12387 11731 12453 11732
rect 12390 11253 12450 11731
rect 12387 11252 12453 11253
rect 12387 11188 12388 11252
rect 12452 11188 12453 11252
rect 12387 11187 12453 11188
rect 12574 9893 12634 13363
rect 12942 13021 13002 21659
rect 13307 21316 13373 21317
rect 13307 21252 13308 21316
rect 13372 21252 13373 21316
rect 13307 21251 13373 21252
rect 12939 13020 13005 13021
rect 12939 12956 12940 13020
rect 13004 12956 13005 13020
rect 12939 12955 13005 12956
rect 12939 12340 13005 12341
rect 12939 12276 12940 12340
rect 13004 12276 13005 12340
rect 12939 12275 13005 12276
rect 12942 11389 13002 12275
rect 13310 11389 13370 21251
rect 14411 21180 14477 21181
rect 14411 21116 14412 21180
rect 14476 21116 14477 21180
rect 14411 21115 14477 21116
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13491 13836 13557 13837
rect 13491 13772 13492 13836
rect 13556 13772 13557 13836
rect 13491 13771 13557 13772
rect 12939 11388 13005 11389
rect 12939 11324 12940 11388
rect 13004 11324 13005 11388
rect 12939 11323 13005 11324
rect 13307 11388 13373 11389
rect 13307 11324 13308 11388
rect 13372 11324 13373 11388
rect 13307 11323 13373 11324
rect 12755 11116 12821 11117
rect 12755 11052 12756 11116
rect 12820 11052 12821 11116
rect 12755 11051 12821 11052
rect 12571 9892 12637 9893
rect 12571 9828 12572 9892
rect 12636 9828 12637 9892
rect 12571 9827 12637 9828
rect 12571 9756 12637 9757
rect 12571 9692 12572 9756
rect 12636 9692 12637 9756
rect 12571 9691 12637 9692
rect 12574 4045 12634 9691
rect 12571 4044 12637 4045
rect 12571 3980 12572 4044
rect 12636 3980 12637 4044
rect 12571 3979 12637 3980
rect 12203 2412 12269 2413
rect 12203 2348 12204 2412
rect 12268 2348 12269 2412
rect 12203 2347 12269 2348
rect 5395 1324 5461 1325
rect 5395 1260 5396 1324
rect 5460 1260 5461 1324
rect 5395 1259 5461 1260
rect 12019 1324 12085 1325
rect 12019 1260 12020 1324
rect 12084 1260 12085 1324
rect 12019 1259 12085 1260
rect 4107 1052 4173 1053
rect 4107 988 4108 1052
rect 4172 988 4173 1052
rect 4107 987 4173 988
rect 3003 644 3069 645
rect 3003 580 3004 644
rect 3068 580 3069 644
rect 3003 579 3069 580
rect 12758 101 12818 11051
rect 12942 4725 13002 11323
rect 12939 4724 13005 4725
rect 12939 4660 12940 4724
rect 13004 4660 13005 4724
rect 12939 4659 13005 4660
rect 13494 4589 13554 13771
rect 13939 13632 14259 14656
rect 14414 14245 14474 21115
rect 14411 14244 14477 14245
rect 14411 14180 14412 14244
rect 14476 14180 14477 14244
rect 14411 14179 14477 14180
rect 14411 14108 14477 14109
rect 14411 14044 14412 14108
rect 14476 14044 14477 14108
rect 14411 14043 14477 14044
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13675 12884 13741 12885
rect 13675 12820 13676 12884
rect 13740 12820 13741 12884
rect 13675 12819 13741 12820
rect 13491 4588 13557 4589
rect 13491 4524 13492 4588
rect 13556 4524 13557 4588
rect 13491 4523 13557 4524
rect 13678 1189 13738 12819
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 14414 12069 14474 14043
rect 14411 12068 14477 12069
rect 14411 12004 14412 12068
rect 14476 12004 14477 12068
rect 14411 12003 14477 12004
rect 14411 11932 14477 11933
rect 14411 11868 14412 11932
rect 14476 11868 14477 11932
rect 14411 11867 14477 11868
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 14414 4181 14474 11867
rect 14598 11661 14658 22475
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 19563 19412 19629 19413
rect 19563 19348 19564 19412
rect 19628 19348 19629 19412
rect 19563 19347 19629 19348
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 17171 17916 17237 17917
rect 17171 17852 17172 17916
rect 17236 17852 17237 17916
rect 17171 17851 17237 17852
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 15699 16556 15765 16557
rect 15699 16492 15700 16556
rect 15764 16492 15765 16556
rect 15699 16491 15765 16492
rect 14963 13836 15029 13837
rect 14963 13772 14964 13836
rect 15028 13772 15029 13836
rect 14963 13771 15029 13772
rect 14779 12068 14845 12069
rect 14779 12004 14780 12068
rect 14844 12004 14845 12068
rect 14779 12003 14845 12004
rect 14595 11660 14661 11661
rect 14595 11596 14596 11660
rect 14660 11596 14661 11660
rect 14595 11595 14661 11596
rect 14595 10844 14661 10845
rect 14595 10780 14596 10844
rect 14660 10780 14661 10844
rect 14595 10779 14661 10780
rect 14411 4180 14477 4181
rect 14411 4116 14412 4180
rect 14476 4116 14477 4180
rect 14411 4115 14477 4116
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 14598 2957 14658 10779
rect 14782 9349 14842 12003
rect 14779 9348 14845 9349
rect 14779 9284 14780 9348
rect 14844 9284 14845 9348
rect 14779 9283 14845 9284
rect 14966 6221 15026 13771
rect 15331 11932 15397 11933
rect 15331 11868 15332 11932
rect 15396 11868 15397 11932
rect 15331 11867 15397 11868
rect 15334 11525 15394 11867
rect 15331 11524 15397 11525
rect 15331 11460 15332 11524
rect 15396 11460 15397 11524
rect 15331 11459 15397 11460
rect 15147 11252 15213 11253
rect 15147 11188 15148 11252
rect 15212 11188 15213 11252
rect 15147 11187 15213 11188
rect 14963 6220 15029 6221
rect 14963 6156 14964 6220
rect 15028 6156 15029 6220
rect 14963 6155 15029 6156
rect 15150 5405 15210 11187
rect 15334 7989 15394 11459
rect 15331 7988 15397 7989
rect 15331 7924 15332 7988
rect 15396 7924 15397 7988
rect 15331 7923 15397 7924
rect 15702 5949 15762 16491
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16067 13292 16133 13293
rect 16067 13228 16068 13292
rect 16132 13228 16133 13292
rect 16067 13227 16133 13228
rect 15883 12340 15949 12341
rect 15883 12276 15884 12340
rect 15948 12276 15949 12340
rect 15883 12275 15949 12276
rect 15886 6901 15946 12275
rect 15883 6900 15949 6901
rect 15883 6836 15884 6900
rect 15948 6836 15949 6900
rect 15883 6835 15949 6836
rect 15699 5948 15765 5949
rect 15699 5884 15700 5948
rect 15764 5884 15765 5948
rect 15699 5883 15765 5884
rect 15147 5404 15213 5405
rect 15147 5340 15148 5404
rect 15212 5340 15213 5404
rect 15147 5339 15213 5340
rect 15702 3365 15762 5883
rect 16070 5813 16130 13227
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16987 12884 17053 12885
rect 16987 12820 16988 12884
rect 17052 12820 17053 12884
rect 16987 12819 17053 12820
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16990 9077 17050 12819
rect 17174 11661 17234 17851
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 17539 16012 17605 16013
rect 17539 15948 17540 16012
rect 17604 15948 17605 16012
rect 17539 15947 17605 15948
rect 17171 11660 17237 11661
rect 17171 11596 17172 11660
rect 17236 11596 17237 11660
rect 17171 11595 17237 11596
rect 17171 11524 17237 11525
rect 17171 11460 17172 11524
rect 17236 11460 17237 11524
rect 17171 11459 17237 11460
rect 16987 9076 17053 9077
rect 16987 9012 16988 9076
rect 17052 9012 17053 9076
rect 16987 9011 17053 9012
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 17174 7173 17234 11459
rect 17542 10573 17602 15947
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19566 15469 19626 19347
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 20483 18052 20549 18053
rect 20483 17988 20484 18052
rect 20548 17988 20549 18052
rect 20483 17987 20549 17988
rect 19747 16692 19813 16693
rect 19747 16628 19748 16692
rect 19812 16628 19813 16692
rect 19747 16627 19813 16628
rect 20299 16692 20365 16693
rect 20299 16628 20300 16692
rect 20364 16628 20365 16692
rect 20299 16627 20365 16628
rect 19563 15468 19629 15469
rect 19563 15404 19564 15468
rect 19628 15404 19629 15468
rect 19563 15403 19629 15404
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19563 14108 19629 14109
rect 19563 14044 19564 14108
rect 19628 14044 19629 14108
rect 19563 14043 19629 14044
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 17723 12612 17789 12613
rect 17723 12548 17724 12612
rect 17788 12548 17789 12612
rect 17723 12547 17789 12548
rect 17539 10572 17605 10573
rect 17539 10508 17540 10572
rect 17604 10508 17605 10572
rect 17539 10507 17605 10508
rect 17539 10436 17605 10437
rect 17539 10372 17540 10436
rect 17604 10372 17605 10436
rect 17539 10371 17605 10372
rect 17355 9348 17421 9349
rect 17355 9284 17356 9348
rect 17420 9284 17421 9348
rect 17355 9283 17421 9284
rect 17171 7172 17237 7173
rect 17171 7108 17172 7172
rect 17236 7108 17237 7172
rect 17171 7107 17237 7108
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16067 5812 16133 5813
rect 16067 5748 16068 5812
rect 16132 5748 16133 5812
rect 16067 5747 16133 5748
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 15699 3364 15765 3365
rect 15699 3300 15700 3364
rect 15764 3300 15765 3364
rect 15699 3299 15765 3300
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 14595 2956 14661 2957
rect 14595 2892 14596 2956
rect 14660 2892 14661 2956
rect 14595 2891 14661 2892
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 17358 2005 17418 9283
rect 17542 7445 17602 10371
rect 17539 7444 17605 7445
rect 17539 7380 17540 7444
rect 17604 7380 17605 7444
rect 17539 7379 17605 7380
rect 17542 4453 17602 7379
rect 17539 4452 17605 4453
rect 17539 4388 17540 4452
rect 17604 4388 17605 4452
rect 17539 4387 17605 4388
rect 17355 2004 17421 2005
rect 17355 1940 17356 2004
rect 17420 1940 17421 2004
rect 17355 1939 17421 1940
rect 17726 1325 17786 12547
rect 19137 12544 19457 13568
rect 19566 13293 19626 14043
rect 19563 13292 19629 13293
rect 19563 13228 19564 13292
rect 19628 13228 19629 13292
rect 19563 13227 19629 13228
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 18643 11660 18709 11661
rect 18643 11596 18644 11660
rect 18708 11596 18709 11660
rect 18643 11595 18709 11596
rect 17907 8396 17973 8397
rect 17907 8332 17908 8396
rect 17972 8332 17973 8396
rect 17907 8331 17973 8332
rect 17910 3093 17970 8331
rect 18646 6901 18706 11595
rect 19137 11456 19457 12480
rect 19750 11522 19810 16627
rect 19931 13836 19997 13837
rect 19931 13772 19932 13836
rect 19996 13772 19997 13836
rect 19931 13771 19997 13772
rect 19934 12450 19994 13771
rect 19934 12390 20178 12450
rect 19750 11462 19994 11522
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19747 11252 19813 11253
rect 19747 11188 19748 11252
rect 19812 11188 19813 11252
rect 19747 11187 19813 11188
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 18827 10300 18893 10301
rect 18827 10236 18828 10300
rect 18892 10236 18893 10300
rect 18827 10235 18893 10236
rect 18643 6900 18709 6901
rect 18643 6836 18644 6900
rect 18708 6836 18709 6900
rect 18643 6835 18709 6836
rect 18830 3909 18890 10235
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 18827 3908 18893 3909
rect 18827 3844 18828 3908
rect 18892 3844 18893 3908
rect 18827 3843 18893 3844
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 17907 3092 17973 3093
rect 17907 3028 17908 3092
rect 17972 3028 17973 3092
rect 17907 3027 17973 3028
rect 19137 2752 19457 3776
rect 19750 3773 19810 11187
rect 19934 11117 19994 11462
rect 19931 11116 19997 11117
rect 19931 11052 19932 11116
rect 19996 11052 19997 11116
rect 19931 11051 19997 11052
rect 19934 8261 19994 11051
rect 20118 10165 20178 12390
rect 20115 10164 20181 10165
rect 20115 10100 20116 10164
rect 20180 10100 20181 10164
rect 20115 10099 20181 10100
rect 19931 8260 19997 8261
rect 19931 8196 19932 8260
rect 19996 8196 19997 8260
rect 19931 8195 19997 8196
rect 20302 4045 20362 16627
rect 20299 4044 20365 4045
rect 20299 3980 20300 4044
rect 20364 3980 20365 4044
rect 20299 3979 20365 3980
rect 20486 3909 20546 17987
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21035 13564 21101 13565
rect 21035 13500 21036 13564
rect 21100 13500 21101 13564
rect 21035 13499 21101 13500
rect 21038 10845 21098 13499
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21035 10844 21101 10845
rect 21035 10780 21036 10844
rect 21100 10780 21101 10844
rect 21035 10779 21101 10780
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 20483 3908 20549 3909
rect 20483 3844 20484 3908
rect 20548 3844 20549 3908
rect 20483 3843 20549 3844
rect 19747 3772 19813 3773
rect 19747 3708 19748 3772
rect 19812 3708 19813 3772
rect 19747 3707 19813 3708
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
rect 17723 1324 17789 1325
rect 17723 1260 17724 1324
rect 17788 1260 17789 1324
rect 17723 1259 17789 1260
rect 13675 1188 13741 1189
rect 13675 1124 13676 1188
rect 13740 1124 13741 1188
rect 13675 1123 13741 1124
rect 12755 100 12821 101
rect 12755 36 12756 100
rect 12820 36 12821 100
rect 12755 35 12821 36
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1649977179
transform 1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1649977179
transform -1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1649977179
transform 1 0 5796 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1649977179
transform 1 0 3864 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1649977179
transform 1 0 4232 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1649977179
transform 1 0 4048 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1649977179
transform 1 0 9016 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1649977179
transform 1 0 9200 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1649977179
transform 1 0 5980 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1649977179
transform 1 0 20332 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1649977179
transform -1 0 21252 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1649977179
transform -1 0 21252 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1649977179
transform -1 0 20516 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1649977179
transform -1 0 21252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1649977179
transform 1 0 20056 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1649977179
transform -1 0 20608 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1649977179
transform -1 0 21252 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1649977179
transform 1 0 19688 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1649977179
transform -1 0 20056 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1649977179
transform 1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1649977179
transform 1 0 17020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1649977179
transform 1 0 13248 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform -1 0 19780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1649977179
transform 1 0 15732 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1649977179
transform 1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform 1 0 12696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform 1 0 14352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1649977179
transform -1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1649977179
transform -1 0 12328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1649977179
transform -1 0 11868 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1649977179
transform 1 0 13248 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1649977179
transform 1 0 14720 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1649977179
transform -1 0 15088 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1649977179
transform 1 0 15088 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1649977179
transform -1 0 16284 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1649977179
transform 1 0 16100 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1649977179
transform -1 0 16468 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1649977179
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1649977179
transform -1 0 19136 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 13524 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 13340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 10856 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 12512 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 10304 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 11040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 8004 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 13892 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 10580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 10488 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 1564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 8372 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 4140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 7636 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 6716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 13892 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 12696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 10120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 13708 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 9936 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 20700 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 20424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 15732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 20240 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 16468 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 21620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 20516 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 21252 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 20516 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 19596 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 21252 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 20332 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 20884 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 16836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 16284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 11040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 11684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 8556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 5428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 10948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 12512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 14996 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 16652 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 13340 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 9108 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 12052 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 11132 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 11316 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 13984 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 4876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 15640 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 15456 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 8832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform -1 0 6716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 4232 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 9016 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 13800 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 11684 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 13616 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform -1 0 10304 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform -1 0 9108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 2668 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 6900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform -1 0 15824 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform -1 0 13616 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 13892 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1649977179
transform -1 0 7820 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1649977179
transform -1 0 13432 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1649977179
transform -1 0 6532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1649977179
transform -1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1649977179
transform -1 0 19688 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1649977179
transform -1 0 18676 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1649977179
transform -1 0 4600 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1649977179
transform -1 0 13708 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1649977179
transform -1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1649977179
transform -1 0 12972 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1649977179
transform -1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1649977179
transform -1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1649977179
transform 1 0 4048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1649977179
transform -1 0 10396 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1649977179
transform -1 0 18492 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1649977179
transform -1 0 18860 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1649977179
transform -1 0 17480 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1649977179
transform -1 0 17296 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1649977179
transform -1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1649977179
transform -1 0 20148 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1649977179
transform -1 0 13984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1649977179
transform -1 0 16560 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1649977179
transform -1 0 20148 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1649977179
transform -1 0 19780 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1649977179
transform -1 0 14352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1649977179
transform -1 0 3680 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1649977179
transform 1 0 2760 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1649977179
transform -1 0 3956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1649977179
transform -1 0 5796 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1649977179
transform -1 0 6348 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1649977179
transform -1 0 2852 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1649977179
transform -1 0 2852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1649977179
transform -1 0 7084 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 17204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 19504 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13708 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 11960 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16652 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12972 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11776 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13156 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 10948 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 10672 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 10304 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 11224 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A0
timestamp 1649977179
transform -1 0 1564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1
timestamp 1649977179
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 10580 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 10764 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11224 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 12788 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15824 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 9568 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10488 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 14628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16100 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 9568 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8004 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1649977179
transform -1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 6716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 5704 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6992 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5612 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7268 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6808 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6624 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 8188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 7728 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10948 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 2668 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 6532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15180 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14352 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 20148 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 18584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 19688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A1
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A0
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 16192 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A1
timestamp 1649977179
transform -1 0 21620 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 14720 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 16192 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 17204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14720 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16008 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 15824 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 18768 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 18400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 19044 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 21252 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 17296 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 20792 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14352 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 18584 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5704 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 6532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 5612 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A1
timestamp 1649977179
transform -1 0 6348 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 3680 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4416 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8096 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 6808 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 7636 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 6624 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 7452 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5244 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1649977179
transform -1 0 11040 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A0
timestamp 1649977179
transform 1 0 9292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A1
timestamp 1649977179
transform -1 0 10856 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A0
timestamp 1649977179
transform 1 0 7820 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A1
timestamp 1649977179
transform 1 0 11040 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A0
timestamp 1649977179
transform 1 0 8004 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 7820 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12328 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10948 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14444 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13064 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11684 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 11132 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 18216 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 18400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 15456 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14904 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 13248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output218_A
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_E_FTB01_A
timestamp 1649977179
transform -1 0 19044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_N_FTB01_A
timestamp 1649977179
transform -1 0 17940 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_S_FTB01_A
timestamp 1649977179
transform -1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_W_FTB01_A
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_122
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1649977179
transform 1 0 18032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_192
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_56
timestamp 1649977179
transform 1 0 6256 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_95
timestamp 1649977179
transform 1 0 9844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_120
timestamp 1649977179
transform 1 0 12144 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_173
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_208
timestamp 1649977179
transform 1 0 20240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_119
timestamp 1649977179
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_126
timestamp 1649977179
transform 1 0 12696 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_202
timestamp 1649977179
transform 1 0 19688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_59
timestamp 1649977179
transform 1 0 6532 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_106
timestamp 1649977179
transform 1 0 10856 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_119
timestamp 1649977179
transform 1 0 12052 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_154
timestamp 1649977179
transform 1 0 15272 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_102
timestamp 1649977179
transform 1 0 10488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_212
timestamp 1649977179
transform 1 0 20608 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_32
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_106
timestamp 1649977179
transform 1 0 10856 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_124
timestamp 1649977179
transform 1 0 12512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_222
timestamp 1649977179
transform 1 0 21528 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_84
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_165
timestamp 1649977179
transform 1 0 16284 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_47
timestamp 1649977179
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_119
timestamp 1649977179
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_162
timestamp 1649977179
transform 1 0 16008 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1649977179
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_73
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_115
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_131
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_156
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_119
timestamp 1649977179
transform 1 0 12052 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_143
timestamp 1649977179
transform 1 0 14260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_148
timestamp 1649977179
transform 1 0 14720 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_192
timestamp 1649977179
transform 1 0 18768 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1649977179
transform 1 0 21528 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_66
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_133
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_196
timestamp 1649977179
transform 1 0 19136 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_218
timestamp 1649977179
transform 1 0 21160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_48
timestamp 1649977179
transform 1 0 5520 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_63
timestamp 1649977179
transform 1 0 6900 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_103
timestamp 1649977179
transform 1 0 10580 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_115
timestamp 1649977179
transform 1 0 11684 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_166
timestamp 1649977179
transform 1 0 16376 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_24
timestamp 1649977179
transform 1 0 3312 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_59
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_109
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_180
timestamp 1649977179
transform 1 0 17664 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp 1649977179
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_55
timestamp 1649977179
transform 1 0 6164 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_58
timestamp 1649977179
transform 1 0 6440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 1649977179
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_134
timestamp 1649977179
transform 1 0 13432 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_179
timestamp 1649977179
transform 1 0 17572 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_222
timestamp 1649977179
transform 1 0 21528 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_22
timestamp 1649977179
transform 1 0 3128 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_162
timestamp 1649977179
transform 1 0 16008 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_187
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_81
timestamp 1649977179
transform 1 0 8556 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_214
timestamp 1649977179
transform 1 0 20792 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_49
timestamp 1649977179
transform 1 0 5612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_163
timestamp 1649977179
transform 1 0 16100 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_175
timestamp 1649977179
transform 1 0 17204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp 1649977179
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_74
timestamp 1649977179
transform 1 0 7912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_118
timestamp 1649977179
transform 1 0 11960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_173
timestamp 1649977179
transform 1 0 17020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_11
timestamp 1649977179
transform 1 0 2116 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_145
timestamp 1649977179
transform 1 0 14444 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_169 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_177
timestamp 1649977179
transform 1 0 17388 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_208
timestamp 1649977179
transform 1 0 20240 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_31
timestamp 1649977179
transform 1 0 3956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_182
timestamp 1649977179
transform 1 0 17848 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_190
timestamp 1649977179
transform 1 0 18584 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_17
timestamp 1649977179
transform 1 0 2668 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_72
timestamp 1649977179
transform 1 0 7728 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_124
timestamp 1649977179
transform 1 0 12512 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_146 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14536 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_150
timestamp 1649977179
transform 1 0 14904 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_154
timestamp 1649977179
transform 1 0 15272 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_191
timestamp 1649977179
transform 1 0 18676 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1649977179
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_201
timestamp 1649977179
transform 1 0 19596 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1649977179
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_118
timestamp 1649977179
transform 1 0 11960 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_131
timestamp 1649977179
transform 1 0 13156 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_134 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_149
timestamp 1649977179
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_152
timestamp 1649977179
transform 1 0 15088 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_14
timestamp 1649977179
transform 1 0 2392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_64
timestamp 1649977179
transform 1 0 6992 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_78
timestamp 1649977179
transform 1 0 8280 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1649977179
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_164
timestamp 1649977179
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_196
timestamp 1649977179
transform 1 0 19136 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1649977179
transform 1 0 19872 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_32
timestamp 1649977179
transform 1 0 4048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_88
timestamp 1649977179
transform 1 0 9200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_120
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1649977179
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_200
timestamp 1649977179
transform 1 0 19504 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_208
timestamp 1649977179
transform 1 0 20240 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_61
timestamp 1649977179
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_133
timestamp 1649977179
transform 1 0 13340 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1649977179
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_201
timestamp 1649977179
transform 1 0 19596 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_206
timestamp 1649977179
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_11
timestamp 1649977179
transform 1 0 2116 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_167
timestamp 1649977179
transform 1 0 16468 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_179
timestamp 1649977179
transform 1 0 17572 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_191
timestamp 1649977179
transform 1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1649977179
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_212
timestamp 1649977179
transform 1 0 20608 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_129
timestamp 1649977179
transform 1 0 12972 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_149 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_155
timestamp 1649977179
transform 1 0 15364 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_158
timestamp 1649977179
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_208
timestamp 1649977179
transform 1 0 20240 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_150
timestamp 1649977179
transform 1 0 14904 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_162
timestamp 1649977179
transform 1 0 16008 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_174
timestamp 1649977179
transform 1 0 17112 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_186
timestamp 1649977179
transform 1 0 18216 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_211
timestamp 1649977179
transform 1 0 20516 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_218
timestamp 1649977179
transform 1 0 21160 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_138
timestamp 1649977179
transform 1 0 13800 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_141
timestamp 1649977179
transform 1 0 14076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_160
timestamp 1649977179
transform 1 0 15824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_176
timestamp 1649977179
transform 1 0 17296 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_180
timestamp 1649977179
transform 1 0 17664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_204
timestamp 1649977179
transform 1 0 19872 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_144
timestamp 1649977179
transform 1 0 14352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_208
timestamp 1649977179
transform 1 0 20240 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_97
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_139
timestamp 1649977179
transform 1 0 13892 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_N_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18768 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1649977179
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1649977179
transform 1 0 3036 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1649977179
transform 1 0 2944 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1649977179
transform 1 0 1840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1649977179
transform 1 0 1840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1649977179
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1649977179
transform 1 0 2668 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1649977179
transform 1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1649977179
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1649977179
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 1840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 2392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 2392 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform -1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform -1 0 19136 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform -1 0 19504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform -1 0 20792 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform -1 0 21068 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform -1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform -1 0 21068 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform -1 0 20792 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform -1 0 21068 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform -1 0 20792 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 20792 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 21068 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 20516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform -1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform -1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform -1 0 20792 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform -1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 21252 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 20608 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform -1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform -1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 12052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform 1 0 14720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 12420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform -1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 13984 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 15548 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform -1 0 16468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 16560 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform -1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1649977179
transform -1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform -1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1649977179
transform -1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform -1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1649977179
transform -1 0 19136 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1649977179
transform 1 0 10120 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1649977179
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1649977179
transform -1 0 9200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1649977179
transform -1 0 12144 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1649977179
transform -1 0 11316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1649977179
transform -1 0 13156 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1649977179
transform -1 0 12880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1649977179
transform -1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1649977179
transform -1 0 13432 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1649977179
transform -1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1649977179
transform -1 0 14720 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1649977179
transform -1 0 14996 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1649977179
transform -1 0 15272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1649977179
transform -1 0 15548 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1649977179
transform -1 0 16100 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1649977179
transform -1 0 16560 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1649977179
transform -1 0 15824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1649977179
transform -1 0 16744 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1649977179
transform -1 0 17296 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1649977179
transform -1 0 18308 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_E_FTB01
timestamp 1649977179
transform -1 0 19136 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_W_FTB01
timestamp 1649977179
transform 1 0 17756 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_E_FTB01
timestamp 1649977179
transform -1 0 18768 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_N_FTB01
timestamp 1649977179
transform -1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_S_FTB01
timestamp 1649977179
transform -1 0 20240 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_W_FTB01
timestamp 1649977179
transform 1 0 16744 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_E_FTB01
timestamp 1649977179
transform -1 0 19136 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_N_FTB01
timestamp 1649977179
transform -1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_S_FTB01
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_W_FTB01
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3220 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 4416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 4784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 6164 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform -1 0 2300 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1649977179
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 19228 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1649977179
transform -1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform -1 0 21620 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1649977179
transform -1 0 19136 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1649977179
transform 1 0 20700 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 21620 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1649977179
transform -1 0 21620 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform -1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1649977179
transform -1 0 21620 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform -1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform -1 0 21620 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1649977179
transform -1 0 21620 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1649977179
transform -1 0 19136 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform -1 0 18952 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1649977179
transform 1 0 20700 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform -1 0 20608 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1649977179
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1649977179
transform -1 0 10212 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1649977179
transform -1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1649977179
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1649977179
transform -1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1649977179
transform -1 0 12144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1649977179
transform -1 0 11408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1649977179
transform -1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform -1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform -1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform -1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1649977179
transform 1 0 6532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform -1 0 7636 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1649977179
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1649977179
transform 1 0 8372 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1649977179
transform -1 0 4692 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1649977179
transform -1 0 3680 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1649977179
transform -1 0 4968 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1649977179
transform 1 0 4968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1649977179
transform -1 0 7912 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1649977179
transform -1 0 8832 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1649977179
transform -1 0 10028 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1649977179
transform -1 0 10120 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1649977179
transform -1 0 9568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1649977179
transform 1 0 10488 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1649977179
transform -1 0 4600 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1649977179
transform 1 0 2944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1649977179
transform -1 0 2944 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1649977179
transform 1 0 2576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1649977179
transform -1 0 6256 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1649977179
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1649977179
transform -1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1649977179
transform 1 0 2944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1649977179
transform 1 0 4232 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1649977179
transform 1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1649977179
transform -1 0 19596 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1649977179
transform -1 0 19872 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1649977179
transform 1 0 6900 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input95
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1649977179
transform 1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1649977179
transform -1 0 4416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1649977179
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1649977179
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1649977179
transform 1 0 20240 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1649977179
transform -1 0 19688 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1649977179
transform -1 0 16560 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input105
timestamp 1649977179
transform 1 0 20700 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input106
timestamp 1649977179
transform -1 0 20700 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input107
timestamp 1649977179
transform 1 0 20700 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1649977179
transform -1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input109
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1649977179
transform -1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1649977179
transform -1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1649977179
transform -1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1649977179
transform -1 0 3220 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1649977179
transform -1 0 3496 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1649977179
transform -1 0 2944 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1649977179
transform 1 0 4968 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1649977179
transform -1 0 2392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1649977179
transform -1 0 2760 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1649977179
transform -1 0 4968 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1649977179
transform -1 0 2392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17388 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14444 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12512 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13892 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10304 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10948 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8648 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8004 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7820 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6900 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 8188 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12880 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11776 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11040 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8832 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8096 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9752 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11040 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 13432 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13800 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 4692 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 3404 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4416 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3036 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3312 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4784 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 4140 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 3312 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 3036 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4232 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4508 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7912 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4232 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10396 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3680 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 2944 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2208 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4232 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5244 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15364 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16836 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17112 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19320 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17296 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17296 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17664 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 18952 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14720 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15548 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14352 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 18492 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17204 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17664 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17572 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14812 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4232 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3496 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 2208 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3220 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4140 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4692 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4140 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4232 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5704 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6440 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7268 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 8740 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11040 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7360 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9384 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10488 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9844 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12052 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 13064 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14168 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13984 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13432 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12236 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15088 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15272 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12604 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1649977179
transform -1 0 12972 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1649977179
transform 1 0 12972 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14444 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12972 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13616 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l2_in_3__293 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13892 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13616 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12512 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 12420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11776 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 11408 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8004 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8740 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 10580 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l2_in_3__296
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 9752 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 9752 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9476 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8004 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1649977179
transform -1 0 8004 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1649977179
transform 1 0 10488 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l2_in_7__298
timestamp 1649977179
transform -1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8004 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1649977179
transform -1 0 7176 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1649977179
transform -1 0 9568 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12144 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11776 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11776 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 10304 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 11408 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_3__299
timestamp 1649977179
transform 1 0 11776 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10672 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1649977179
transform -1 0 10580 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8740 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1649977179
transform -1 0 8096 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8004 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8832 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l2_in_3__294
timestamp 1649977179
transform 1 0 10580 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9936 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1649977179
transform -1 0 10212 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13248 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13524 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12512 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12512 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_3__295
timestamp 1649977179
transform 1 0 12052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1649977179
transform -1 0 12420 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12604 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1649977179
transform -1 0 12696 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13616 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16192 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14996 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1649977179
transform -1 0 15732 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13432 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_33.mux_l1_in_3__297
timestamp 1649977179
transform 1 0 14996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1649977179
transform 1 0 14168 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15824 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14904 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16100 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5336 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform -1 0 4784 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1649977179
transform -1 0 3864 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5336 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5244 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 7176 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l2_in_3__300
timestamp 1649977179
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10212 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2024 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7176 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5520 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5336 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 2852 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l2_in_3__303
timestamp 1649977179
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2392 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4324 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3220 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3680 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6532 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5704 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5152 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5428 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1649977179
transform 1 0 2208 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1649977179
transform 1 0 1932 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1649977179
transform 1 0 1840 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l2_in_7__277
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1649977179
transform -1 0 2484 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4600 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1649977179
transform -1 0 2208 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1649977179
transform -1 0 2484 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3404 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1649977179
transform -1 0 2484 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7268 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6992 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6440 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6716 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5796 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l2_in_3__278
timestamp 1649977179
transform -1 0 4508 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4692 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5428 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6256 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6900 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7912 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7820 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6532 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6900 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4968 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l2_in_3__301
timestamp 1649977179
transform 1 0 5704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4876 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2392 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9476 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9016 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l2_in_3__302
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3220 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3036 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2208 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5244 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l1_in_3__276
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1649977179
transform -1 0 3312 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4324 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3496 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16560 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 19044 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1649977179
transform -1 0 18216 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1649977179
transform -1 0 15272 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16560 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18308 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 18216 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_3__279
timestamp 1649977179
transform 1 0 19044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 18216 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 18584 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1649977179
transform -1 0 17664 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1649977179
transform 1 0 20700 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1649977179
transform -1 0 16560 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19780 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 19044 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l2_in_3__281
timestamp 1649977179
transform -1 0 17112 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 18952 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19412 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 19412 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19136 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13156 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13340 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20700 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1649977179
transform -1 0 21436 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1649977179
transform -1 0 21436 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1649977179
transform 1 0 20424 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1649977179
transform -1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1649977179
transform -1 0 17296 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l2_in_7__284
timestamp 1649977179
transform -1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1649977179
transform 1 0 20056 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20332 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1649977179
transform 1 0 19504 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 20240 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1649977179
transform -1 0 20240 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1649977179
transform -1 0 20332 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20424 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15732 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14720 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l2_in_3__285
timestamp 1649977179
transform -1 0 16376 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16376 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15180 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 16100 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20792 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15732 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16192 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16376 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16468 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1649977179
transform -1 0 16560 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1649977179
transform 1 0 18308 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l2_in_3__280
timestamp 1649977179
transform -1 0 18768 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17848 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1649977179
transform -1 0 18032 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18032 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18584 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1649977179
transform 1 0 18584 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18032 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform -1 0 18308 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l2_in_3__282
timestamp 1649977179
transform -1 0 20240 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1649977179
transform 1 0 19780 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1649977179
transform -1 0 19964 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1649977179
transform 1 0 20056 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19964 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15732 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1649977179
transform 1 0 19780 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1649977179
transform -1 0 14996 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1649977179
transform 1 0 17756 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l1_in_3__283
timestamp 1649977179
transform -1 0 17756 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16560 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 16560 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19504 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3220 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3220 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1649977179
transform 1 0 4600 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1649977179
transform 1 0 6072 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_3__286
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3680 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3220 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3772 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 4324 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4692 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7084 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6808 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1649977179
transform 1 0 6624 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5796 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6164 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_2.mux_l2_in_3__288
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1649977179
transform -1 0 6256 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10580 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7912 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1649977179
transform 1 0 9016 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1649977179
transform 1 0 9108 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1649977179
transform 1 0 8188 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l2_in_7__291
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1649977179
transform -1 0 8832 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7268 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8280 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1649977179
transform -1 0 9108 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1649977179
transform -1 0 8832 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1649977179
transform -1 0 11040 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10396 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7452 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9936 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9016 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9844 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l2_in_3__292
timestamp 1649977179
transform 1 0 10672 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9844 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10304 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9936 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10304 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10580 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13432 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12236 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12696 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_16.mux_l2_in_3__287
timestamp 1649977179
transform 1 0 12696 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11684 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12880 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11408 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12604 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16376 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15640 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16284 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15916 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1649977179
transform -1 0 15088 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l2_in_3__289
timestamp 1649977179
transform -1 0 16192 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1649977179
transform -1 0 14628 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14444 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12512 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13432 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13432 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1649977179
transform 1 0 13432 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_32.mux_l1_in_3__290
timestamp 1649977179
transform -1 0 13984 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13156 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 13432 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13524 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14720 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform -1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform -1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform -1 0 2116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform -1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1649977179
transform -1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform -1 0 1748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform -1 0 2116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform -1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1649977179
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1649977179
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1649977179
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1649977179
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1649977179
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1649977179
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1649977179
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1649977179
transform 1 0 20884 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1649977179
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1649977179
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1649977179
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1649977179
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1649977179
transform 1 0 20884 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1649977179
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1649977179
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1649977179
transform 1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1649977179
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1649977179
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1649977179
transform -1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1649977179
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1649977179
transform 1 0 10120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1649977179
transform 1 0 17388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1649977179
transform 1 0 18492 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1649977179
transform -1 0 11684 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1649977179
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1649977179
transform 1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1649977179
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1649977179
transform -1 0 13156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1649977179
transform 1 0 13156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1649977179
transform -1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1649977179
transform 1 0 14444 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1649977179
transform -1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1649977179
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1649977179
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1649977179
transform -1 0 2116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1649977179
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1649977179
transform -1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1649977179
transform -1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1649977179
transform -1 0 19780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1649977179
transform -1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output215
timestamp 1649977179
transform -1 0 20332 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output216
timestamp 1649977179
transform -1 0 19688 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output217
timestamp 1649977179
transform -1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output218
timestamp 1649977179
transform 1 0 4600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1649977179
transform -1 0 20700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1649977179
transform -1 0 2116 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_0_FTB00
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_E_FTB01
timestamp 1649977179
transform 1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_W_FTB01
timestamp 1649977179
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1649977179
transform 1 0 20700 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1649977179
transform 1 0 20608 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1649977179
transform -1 0 20240 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_E_FTB01
timestamp 1649977179
transform -1 0 18216 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_N_FTB01
timestamp 1649977179
transform -1 0 19964 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_S_FTB01
timestamp 1649977179
transform 1 0 20700 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_W_FTB01
timestamp 1649977179
transform 1 0 17480 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater223
timestamp 1649977179
transform -1 0 10304 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater224
timestamp 1649977179
transform 1 0 3864 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater225
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater226
timestamp 1649977179
transform -1 0 6164 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater227
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater228
timestamp 1649977179
transform -1 0 19136 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater229
timestamp 1649977179
transform -1 0 21620 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater230
timestamp 1649977179
transform 1 0 15364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater231
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater232
timestamp 1649977179
transform 1 0 6624 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater233
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater234
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater235
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater236
timestamp 1649977179
transform -1 0 8004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater237
timestamp 1649977179
transform -1 0 12328 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater238
timestamp 1649977179
transform -1 0 16468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater239
timestamp 1649977179
transform -1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater240
timestamp 1649977179
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater241
timestamp 1649977179
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater242
timestamp 1649977179
transform 1 0 7636 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater243
timestamp 1649977179
transform -1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater244
timestamp 1649977179
transform -1 0 9200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater245
timestamp 1649977179
transform 1 0 8004 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater246
timestamp 1649977179
transform -1 0 9384 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater247
timestamp 1649977179
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater248
timestamp 1649977179
transform 1 0 4968 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater249
timestamp 1649977179
transform 1 0 4048 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater250
timestamp 1649977179
transform 1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater251
timestamp 1649977179
transform 1 0 5888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater252
timestamp 1649977179
transform 1 0 6440 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater253
timestamp 1649977179
transform 1 0 8372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater254
timestamp 1649977179
transform 1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater255
timestamp 1649977179
transform 1 0 3864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater256
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater257
timestamp 1649977179
transform 1 0 12972 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater258
timestamp 1649977179
transform 1 0 14536 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater259
timestamp 1649977179
transform 1 0 13524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater260
timestamp 1649977179
transform -1 0 14536 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater261
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater262
timestamp 1649977179
transform 1 0 13432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater263
timestamp 1649977179
transform -1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater264
timestamp 1649977179
transform 1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater265
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater266
timestamp 1649977179
transform 1 0 13524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater267
timestamp 1649977179
transform -1 0 15272 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater268
timestamp 1649977179
transform 1 0 15272 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater269
timestamp 1649977179
transform 1 0 17020 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater270
timestamp 1649977179
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater271
timestamp 1649977179
transform 1 0 18676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater272
timestamp 1649977179
transform -1 0 18676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater273
timestamp 1649977179
transform -1 0 17572 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater274
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater275
timestamp 1649977179
transform 1 0 16928 0 -1 15232
box -38 -48 314 592
<< labels >>
flabel metal2 s 18234 22200 18290 23000 0 FreeSans 224 90 0 0 Test_en_N_out
port 0 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 Test_en_S_in
port 1 nsew signal input
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_42_
port 4 nsew signal input
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_43_
port 5 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_44_
port 6 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_45_
port 7 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_46_
port 8 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_47_
port 9 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_48_
port 10 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_49_
port 11 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 ccff_head
port 12 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 ccff_tail
port 13 nsew signal tristate
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 14 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 15 nsew signal input
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 16 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 17 nsew signal input
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 18 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 19 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 20 nsew signal input
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 21 nsew signal input
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 22 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 23 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 24 nsew signal input
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 25 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 26 nsew signal input
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 27 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 28 nsew signal input
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 29 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 30 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 31 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 32 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 33 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 34 nsew signal tristate
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 35 nsew signal tristate
flabel metal3 s 0 16464 800 16584 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 36 nsew signal tristate
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 37 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 38 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 39 nsew signal tristate
flabel metal3 s 0 18096 800 18216 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 40 nsew signal tristate
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 41 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 42 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 43 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 44 nsew signal tristate
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 45 nsew signal tristate
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 46 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 47 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 48 nsew signal tristate
flabel metal3 s 0 14016 800 14136 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 49 nsew signal tristate
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 50 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 51 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 52 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 53 nsew signal tristate
flabel metal3 s 22200 3816 23000 3936 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 54 nsew signal input
flabel metal3 s 22200 7896 23000 8016 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 55 nsew signal input
flabel metal3 s 22200 8304 23000 8424 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 56 nsew signal input
flabel metal3 s 22200 8712 23000 8832 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 57 nsew signal input
flabel metal3 s 22200 9120 23000 9240 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 58 nsew signal input
flabel metal3 s 22200 9528 23000 9648 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 59 nsew signal input
flabel metal3 s 22200 9936 23000 10056 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 60 nsew signal input
flabel metal3 s 22200 10344 23000 10464 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 61 nsew signal input
flabel metal3 s 22200 10752 23000 10872 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 62 nsew signal input
flabel metal3 s 22200 11160 23000 11280 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 63 nsew signal input
flabel metal3 s 22200 11568 23000 11688 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 64 nsew signal input
flabel metal3 s 22200 4224 23000 4344 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 65 nsew signal input
flabel metal3 s 22200 4632 23000 4752 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 66 nsew signal input
flabel metal3 s 22200 5040 23000 5160 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 67 nsew signal input
flabel metal3 s 22200 5448 23000 5568 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 68 nsew signal input
flabel metal3 s 22200 5856 23000 5976 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 69 nsew signal input
flabel metal3 s 22200 6264 23000 6384 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 70 nsew signal input
flabel metal3 s 22200 6672 23000 6792 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 71 nsew signal input
flabel metal3 s 22200 7080 23000 7200 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 72 nsew signal input
flabel metal3 s 22200 7488 23000 7608 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 73 nsew signal input
flabel metal3 s 22200 11976 23000 12096 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 74 nsew signal tristate
flabel metal3 s 22200 16056 23000 16176 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 75 nsew signal tristate
flabel metal3 s 22200 16464 23000 16584 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 76 nsew signal tristate
flabel metal3 s 22200 16872 23000 16992 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 77 nsew signal tristate
flabel metal3 s 22200 17280 23000 17400 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 78 nsew signal tristate
flabel metal3 s 22200 17688 23000 17808 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 79 nsew signal tristate
flabel metal3 s 22200 18096 23000 18216 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 80 nsew signal tristate
flabel metal3 s 22200 18504 23000 18624 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 81 nsew signal tristate
flabel metal3 s 22200 18912 23000 19032 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 82 nsew signal tristate
flabel metal3 s 22200 19320 23000 19440 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 83 nsew signal tristate
flabel metal3 s 22200 19728 23000 19848 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 84 nsew signal tristate
flabel metal3 s 22200 12384 23000 12504 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 85 nsew signal tristate
flabel metal3 s 22200 12792 23000 12912 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 86 nsew signal tristate
flabel metal3 s 22200 13200 23000 13320 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 87 nsew signal tristate
flabel metal3 s 22200 13608 23000 13728 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 88 nsew signal tristate
flabel metal3 s 22200 14016 23000 14136 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 89 nsew signal tristate
flabel metal3 s 22200 14424 23000 14544 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 90 nsew signal tristate
flabel metal3 s 22200 14832 23000 14952 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 91 nsew signal tristate
flabel metal3 s 22200 15240 23000 15360 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 92 nsew signal tristate
flabel metal3 s 22200 15648 23000 15768 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 93 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 94 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 95 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 96 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 97 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 98 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 99 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 100 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 101 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 102 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 103 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 104 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 105 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 106 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 107 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 108 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 109 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 110 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 111 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 112 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 113 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 114 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 115 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 116 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 117 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 118 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 119 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 120 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 121 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 122 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 123 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 124 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 125 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 126 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 127 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 128 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 129 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 130 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 131 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 132 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 133 nsew signal tristate
flabel metal2 s 3514 22200 3570 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 134 nsew signal input
flabel metal2 s 7194 22200 7250 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 135 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 136 nsew signal input
flabel metal2 s 7930 22200 7986 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 137 nsew signal input
flabel metal2 s 8298 22200 8354 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 138 nsew signal input
flabel metal2 s 8666 22200 8722 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 139 nsew signal input
flabel metal2 s 9034 22200 9090 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 140 nsew signal input
flabel metal2 s 9402 22200 9458 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 141 nsew signal input
flabel metal2 s 9770 22200 9826 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 142 nsew signal input
flabel metal2 s 10138 22200 10194 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 143 nsew signal input
flabel metal2 s 10506 22200 10562 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 144 nsew signal input
flabel metal2 s 3882 22200 3938 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 145 nsew signal input
flabel metal2 s 4250 22200 4306 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 146 nsew signal input
flabel metal2 s 4618 22200 4674 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 147 nsew signal input
flabel metal2 s 4986 22200 5042 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 148 nsew signal input
flabel metal2 s 5354 22200 5410 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 149 nsew signal input
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 150 nsew signal input
flabel metal2 s 6090 22200 6146 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 151 nsew signal input
flabel metal2 s 6458 22200 6514 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 152 nsew signal input
flabel metal2 s 6826 22200 6882 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 153 nsew signal input
flabel metal2 s 10874 22200 10930 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 154 nsew signal tristate
flabel metal2 s 14554 22200 14610 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 155 nsew signal tristate
flabel metal2 s 14922 22200 14978 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 156 nsew signal tristate
flabel metal2 s 15290 22200 15346 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 157 nsew signal tristate
flabel metal2 s 15658 22200 15714 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 158 nsew signal tristate
flabel metal2 s 16026 22200 16082 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 159 nsew signal tristate
flabel metal2 s 16394 22200 16450 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 160 nsew signal tristate
flabel metal2 s 16762 22200 16818 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 161 nsew signal tristate
flabel metal2 s 17130 22200 17186 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 162 nsew signal tristate
flabel metal2 s 17498 22200 17554 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 163 nsew signal tristate
flabel metal2 s 17866 22200 17922 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 164 nsew signal tristate
flabel metal2 s 11242 22200 11298 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 165 nsew signal tristate
flabel metal2 s 11610 22200 11666 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 166 nsew signal tristate
flabel metal2 s 11978 22200 12034 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 167 nsew signal tristate
flabel metal2 s 12346 22200 12402 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 168 nsew signal tristate
flabel metal2 s 12714 22200 12770 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 169 nsew signal tristate
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 170 nsew signal tristate
flabel metal2 s 13450 22200 13506 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 171 nsew signal tristate
flabel metal2 s 13818 22200 13874 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 172 nsew signal tristate
flabel metal2 s 14186 22200 14242 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 173 nsew signal tristate
flabel metal3 s 22200 20136 23000 20256 0 FreeSans 480 0 0 0 clk_1_E_out
port 174 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 clk_1_N_in
port 175 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 clk_1_W_out
port 176 nsew signal tristate
flabel metal3 s 22200 20544 23000 20664 0 FreeSans 480 0 0 0 clk_2_E_out
port 177 nsew signal tristate
flabel metal2 s 18970 22200 19026 23000 0 FreeSans 224 90 0 0 clk_2_N_in
port 178 nsew signal input
flabel metal2 s 21178 22200 21234 23000 0 FreeSans 224 90 0 0 clk_2_N_out
port 179 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 clk_2_S_out
port 180 nsew signal tristate
flabel metal3 s 0 20544 800 20664 0 FreeSans 480 0 0 0 clk_2_W_out
port 181 nsew signal tristate
flabel metal3 s 22200 20952 23000 21072 0 FreeSans 480 0 0 0 clk_3_E_out
port 182 nsew signal tristate
flabel metal2 s 19338 22200 19394 23000 0 FreeSans 224 90 0 0 clk_3_N_in
port 183 nsew signal input
flabel metal2 s 21546 22200 21602 23000 0 FreeSans 224 90 0 0 clk_3_N_out
port 184 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 clk_3_S_out
port 185 nsew signal tristate
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 clk_3_W_out
port 186 nsew signal tristate
flabel metal3 s 0 552 800 672 0 FreeSans 480 0 0 0 left_bottom_grid_pin_34_
port 187 nsew signal input
flabel metal3 s 0 960 800 1080 0 FreeSans 480 0 0 0 left_bottom_grid_pin_35_
port 188 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 left_bottom_grid_pin_36_
port 189 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 left_bottom_grid_pin_37_
port 190 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 left_bottom_grid_pin_38_
port 191 nsew signal input
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 left_bottom_grid_pin_39_
port 192 nsew signal input
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 left_bottom_grid_pin_40_
port 193 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 left_bottom_grid_pin_41_
port 194 nsew signal input
flabel metal2 s 19706 22200 19762 23000 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 195 nsew signal input
flabel metal3 s 22200 21360 23000 21480 0 FreeSans 480 0 0 0 prog_clk_1_E_out
port 196 nsew signal tristate
flabel metal2 s 20074 22200 20130 23000 0 FreeSans 224 90 0 0 prog_clk_1_N_in
port 197 nsew signal input
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 prog_clk_1_W_out
port 198 nsew signal tristate
flabel metal3 s 22200 21768 23000 21888 0 FreeSans 480 0 0 0 prog_clk_2_E_out
port 199 nsew signal tristate
flabel metal2 s 20442 22200 20498 23000 0 FreeSans 224 90 0 0 prog_clk_2_N_in
port 200 nsew signal input
flabel metal2 s 21914 22200 21970 23000 0 FreeSans 224 90 0 0 prog_clk_2_N_out
port 201 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 prog_clk_2_S_out
port 202 nsew signal tristate
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 prog_clk_2_W_out
port 203 nsew signal tristate
flabel metal3 s 22200 22176 23000 22296 0 FreeSans 480 0 0 0 prog_clk_3_E_out
port 204 nsew signal tristate
flabel metal2 s 20810 22200 20866 23000 0 FreeSans 224 90 0 0 prog_clk_3_N_in
port 205 nsew signal input
flabel metal2 s 22282 22200 22338 23000 0 FreeSans 224 90 0 0 prog_clk_3_N_out
port 206 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 prog_clk_3_S_out
port 207 nsew signal tristate
flabel metal3 s 0 22176 800 22296 0 FreeSans 480 0 0 0 prog_clk_3_W_out
port 208 nsew signal tristate
flabel metal3 s 22200 552 23000 672 0 FreeSans 480 0 0 0 right_bottom_grid_pin_34_
port 209 nsew signal input
flabel metal3 s 22200 960 23000 1080 0 FreeSans 480 0 0 0 right_bottom_grid_pin_35_
port 210 nsew signal input
flabel metal3 s 22200 1368 23000 1488 0 FreeSans 480 0 0 0 right_bottom_grid_pin_36_
port 211 nsew signal input
flabel metal3 s 22200 1776 23000 1896 0 FreeSans 480 0 0 0 right_bottom_grid_pin_37_
port 212 nsew signal input
flabel metal3 s 22200 2184 23000 2304 0 FreeSans 480 0 0 0 right_bottom_grid_pin_38_
port 213 nsew signal input
flabel metal3 s 22200 2592 23000 2712 0 FreeSans 480 0 0 0 right_bottom_grid_pin_39_
port 214 nsew signal input
flabel metal3 s 22200 3000 23000 3120 0 FreeSans 480 0 0 0 right_bottom_grid_pin_40_
port 215 nsew signal input
flabel metal3 s 22200 3408 23000 3528 0 FreeSans 480 0 0 0 right_bottom_grid_pin_41_
port 216 nsew signal input
flabel metal2 s 570 22200 626 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_42_
port 217 nsew signal input
flabel metal2 s 938 22200 994 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_43_
port 218 nsew signal input
flabel metal2 s 1306 22200 1362 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_44_
port 219 nsew signal input
flabel metal2 s 1674 22200 1730 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_45_
port 220 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_46_
port 221 nsew signal input
flabel metal2 s 2410 22200 2466 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_47_
port 222 nsew signal input
flabel metal2 s 2778 22200 2834 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_48_
port 223 nsew signal input
flabel metal2 s 3146 22200 3202 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_49_
port 224 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
