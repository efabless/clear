* NGSPICE file created from sb_0__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

.subckt sb_0__1_ VGND VPWR bottom_left_grid_pin_1_ ccff_head ccff_tail chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] prog_clk_0_E_in right_bottom_grid_pin_34_ right_bottom_grid_pin_35_
+ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_ right_bottom_grid_pin_39_
+ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ top_left_grid_pin_1_
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_20.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_2
XFILLER_9_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_3.mux_l1_in_1_ input5/X input17/X mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__124__A _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_36.sky130_fd_sc_hd__buf_4_0_ mux_right_track_36.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _084_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input55_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_0.mux_l2_in_1__162 VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/A0
+ mux_right_track_0.mux_l2_in_1__162/LO sky130_fd_sc_hd__conb_1
XANTENNA__119__A _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_114_ _114_/A VGND VGND VPWR VPWR _114_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l1_in_0_ _104_/A _095_/A mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input18_A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput75 _077_/X VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _087_/A sky130_fd_sc_hd__clkbuf_1
Xoutput97 _099_/X VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
Xoutput86 _069_/X VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_34.mux_l2_in_0__143 VGND VGND VPWR VPWR mux_right_track_34.mux_l2_in_0_/A0
+ mux_right_track_34.mux_l2_in_0__143/LO sky130_fd_sc_hd__conb_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_3.mux_l1_in_0_ _100_/A _091_/A mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l1_in_1__133 VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/A0
+ mux_right_track_16.mux_l1_in_1__133/LO sky130_fd_sc_hd__conb_1
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_10.mux_l2_in_0__A0 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_26.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input48_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_6.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_113_ _113_/A VGND VGND VPWR VPWR _113_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput76 _078_/X VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
Xoutput98 _100_/X VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xoutput87 _070_/X VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_6.mux_l1_in_1__A0 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_0.mux_l2_in_1__148 VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/A0
+ mux_top_track_0.mux_l2_in_1__148/LO sky130_fd_sc_hd__conb_1
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_10.mux_l3_in_0_ mux_right_track_10.mux_l2_in_1_/X mux_right_track_10.mux_l2_in_0_/X
+ mux_right_track_10.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_10.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_24.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_26.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_112_ _112_/A VGND VGND VPWR VPWR _112_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input60_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_10.mux_l2_in_1_ mux_right_track_10.mux_l2_in_1_/A0 _116_/A mux_right_track_10.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_17.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_20.mux_l1_in_1__136 VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_1_/A0
+ mux_right_track_20.mux_l1_in_1__136/LO sky130_fd_sc_hd__conb_1
XFILLER_25_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput77 _079_/X VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xoutput88 _071_/X VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
Xoutput99 _101_/X VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
XANTENNA_input23_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l1_in_1__A1 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_3__A1 _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xprog_clk_0_FTB00 prog_clk_0_E_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_2_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_111_ _111_/A VGND VGND VPWR VPWR _111_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input53_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_10.mux_l2_in_0_ input64/X mux_right_track_10.mux_l1_in_0_/X mux_right_track_10.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_25_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_12.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xoutput78 _080_/X VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
Xoutput89 _072_/X VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
XANTENNA_input16_A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l2_in_1_ mux_right_track_8.mux_l2_in_1_/A0 _115_/A mux_right_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ mux_top_track_0.mux_l2_in_1_/A0 mux_top_track_0.mux_l1_in_2_/X
+ mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_1.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input8_A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_22.mux_l1_in_0__A0 _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_2_ _119_/A _109_/A mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _114_/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_12.mux_l2_in_1__164 VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_1_/A0
+ mux_right_track_12.mux_l2_in_1__164/LO sky130_fd_sc_hd__conb_1
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_14.mux_l1_in_0__A1 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_5 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_110_ _110_/A VGND VGND VPWR VPWR _110_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input46_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_24.mux_l2_in_1__S mux_top_track_24.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_8.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _106_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_12.mux_l2_in_1__A1 _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_10.mux_l1_in_0_ input45/X _096_/A mux_right_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xoutput79 _081_/X VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
XFILLER_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_8.mux_l2_in_0_ input63/X mux_right_track_8.mux_l1_in_0_/X mux_right_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_22.mux_l2_in_0_ mux_right_track_22.mux_l1_in_1_/X mux_right_track_22.mux_l1_in_0_/X
+ mux_right_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_22.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__D mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l2_in_1__154 VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/A0
+ mux_top_track_8.mux_l2_in_1__154/LO sky130_fd_sc_hd__conb_1
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_17 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_22.mux_l1_in_0__A1 _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_0.mux_l1_in_1_ input9/X input21/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_22.mux_l1_in_1_ mux_right_track_22.mux_l1_in_1_/A0 _124_/A mux_right_track_22.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__091__A _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_5.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_14_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_17.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input39_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_10.sky130_fd_sc_hd__buf_4_0_ mux_right_track_10.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _071_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A0 _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_10.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_30.mux_l1_in_0__A1 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_33.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _102_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input21_A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l1_in_0_ _095_/A input60/X mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_28.mux_l2_in_0__140 VGND VGND VPWR VPWR mux_right_track_28.mux_l2_in_0_/A0
+ mux_right_track_28.mux_l2_in_0__140/LO sky130_fd_sc_hd__conb_1
XANTENNA__089__A _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_0_ input14/X input71/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input69_A right_bottom_grid_pin_40_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_22.mux_l1_in_0_ _085_/A _104_/A mux_right_track_22.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_34.mux_l2_in_0_ mux_right_track_34.mux_l2_in_0_/A0 mux_right_track_34.mux_l1_in_0_/X
+ mux_right_track_34.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_34.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _070_/A sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_25.mux_l2_in_1_ mux_bottom_track_25.mux_l2_in_1_/A0 input8/X mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_099_ _099_/A VGND VGND VPWR VPWR _099_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__097__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input51_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_1_ mux_bottom_track_9.mux_l2_in_1_/A0 mux_bottom_track_9.mux_l1_in_2_/X
+ mux_bottom_track_9.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _082_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_32.mux_l2_in_0__142 VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/A0
+ mux_right_track_32.mux_l2_in_0__142/LO sky130_fd_sc_hd__conb_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_9.mux_l1_in_2_ input1/X input10/X mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input14_A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_26.sky130_fd_sc_hd__buf_4_0_ mux_right_track_26.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input6_A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_9.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_30.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_30.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_34.mux_l1_in_0_ input34/X input68/X mux_right_track_34.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_34.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_098_ _098_/A VGND VGND VPWR VPWR _098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l1_in_1_ input20/X input3/X mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input44_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_0_ mux_bottom_track_9.mux_l1_in_1_/X mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_6.mux_l1_in_3__146 VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_3_/A0
+ mux_right_track_6.mux_l1_in_3__146/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l1_in_1_ input22/X input15/X mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_28.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_30.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_097_ _097_/A VGND VGND VPWR VPWR _097_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l2_in_1_ mux_top_track_16.mux_l2_in_1_/A0 _124_/A mux_top_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l1_in_0_ _105_/A _096_/A mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input37_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_36.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_36.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_9.mux_l1_in_0_ _103_/A _093_/A mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _090_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input67_A right_bottom_grid_pin_38_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__100__A _100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_096_ _096_/A VGND VGND VPWR VPWR _096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_079_ _079_/A VGND VGND VPWR VPWR _079_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_3_ mux_right_track_4.mux_l1_in_3_/A0 _112_/A mux_right_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_16.mux_l1_in_1_ _115_/A input13/X mux_top_track_16.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_34.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_36.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__103__A _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input12_A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_28.mux_l1_in_0__A1 input65/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_10.mux_l2_in_1__163 VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_1_/A0
+ mux_right_track_10.mux_l2_in_1__163/LO sky130_fd_sc_hd__conb_1
XANTENNA_input4_A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_1_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_095_ _095_/A VGND VGND VPWR VPWR _095_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__111__A _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_078_ _078_/A VGND VGND VPWR VPWR _078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_2_ input69/X input67/X mux_right_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input42_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l1_in_0_ input6/X input18/X mux_top_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__109__A _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_094_ _094_/A VGND VGND VPWR VPWR _094_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ _077_/A VGND VGND VPWR VPWR _077_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_16.mux_l1_in_1_ mux_right_track_16.mux_l1_in_1_/A0 _120_/A mux_right_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_4.mux_l1_in_1_ input65/X input63/X mux_right_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input35_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 _100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_1__S mux_bottom_track_3.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.mux_l1_in_1__159 VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/A0
+ mux_bottom_track_33.mux_l1_in_1__159/LO sky130_fd_sc_hd__conb_1
XANTENNA__117__A _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_22.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_2
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input65_A right_bottom_grid_pin_36_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_093_ _093_/A VGND VGND VPWR VPWR _093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput1 bottom_left_grid_pin_1_ VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_3.mux_l2_in_1__158 VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/A0
+ mux_bottom_track_3.mux_l2_in_1__158/LO sky130_fd_sc_hd__conb_1
XFILLER_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_076_ _076_/A VGND VGND VPWR VPWR _076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_0_ input67/X _100_/A mux_right_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_0_ _092_/A input54/X mux_right_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_28.mux_l2_in_0_ mux_right_track_28.mux_l2_in_0_/A0 mux_right_track_28.mux_l1_in_0_/X
+ mux_right_track_28.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_28.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _068_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input28_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_30.mux_l2_in_0__141 VGND VGND VPWR VPWR mux_right_track_30.mux_l2_in_0_/A0
+ mux_right_track_30.mux_l2_in_0__141/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_10.mux_l1_in_0__A1 _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_30.mux_l2_in_0_ mux_right_track_30.mux_l2_in_0_/A0 mux_right_track_30.mux_l1_in_0_/X
+ mux_right_track_30.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_30.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2__S mux_right_track_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0__A0 _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput70 right_bottom_grid_pin_41_ VGND VGND VPWR VPWR _085_/A sky130_fd_sc_hd__clkbuf_2
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _094_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_32_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_20.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l2_in_1_/A0 mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input10_A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input2_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input58_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_092_ _092_/A VGND VGND VPWR VPWR _092_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_22.sky130_fd_sc_hd__buf_4_0_ mux_right_track_22.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__clkbuf_1
Xinput2 ccff_head VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l1_in_2_ input1/X input11/X mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_075_ _075_/A VGND VGND VPWR VPWR _075_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_28.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_28.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _074_/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_4.mux_l1_in_3__145 VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_3_/A0
+ mux_right_track_4.mux_l1_in_3__145/LO sky130_fd_sc_hd__conb_1
XFILLER_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput71 top_left_grid_pin_1_ VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput60 chany_top_in[7] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input40_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_28.mux_l1_in_0_ input25/X input65/X mux_right_track_28.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_28.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 input67/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_30.mux_l1_in_0_ input40/X input66/X mux_right_track_30.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_30.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_091_ _091_/A VGND VGND VPWR VPWR _091_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 chanx_right_in[0] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_5.mux_l1_in_1_ input4/X input16/X mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input70_A right_bottom_grid_pin_41_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_074_ _074_/A VGND VGND VPWR VPWR _074_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_26.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_28.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_12.mux_l2_in_0__A0 input65/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput61 chany_top_in[8] VGND VGND VPWR VPWR _095_/A sky130_fd_sc_hd__clkbuf_2
Xinput50 chany_top_in[16] VGND VGND VPWR VPWR _103_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_E_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input33_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_109_ _109_/A VGND VGND VPWR VPWR _109_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_0.mux_l1_in_2__A1 _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l2_in_1__147 VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/A0
+ mux_right_track_8.mux_l2_in_1__147/LO sky130_fd_sc_hd__conb_1
XFILLER_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ output72/A VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_090_ _090_/A VGND VGND VPWR VPWR _090_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _088_/A sky130_fd_sc_hd__clkbuf_1
Xinput4 chanx_right_in[10] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l1_in_0_ _101_/A _092_/A mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l1_in_1_ mux_bottom_track_33.mux_l1_in_1_/A0 input7/X mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input63_A right_bottom_grid_pin_34_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_073_ _073_/A VGND VGND VPWR VPWR _073_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_125_ _125_/A VGND VGND VPWR VPWR _125_/X sky130_fd_sc_hd__clkbuf_1
Xinput51 chany_top_in[17] VGND VGND VPWR VPWR _104_/A sky130_fd_sc_hd__clkbuf_2
Xinput62 chany_top_in[9] VGND VGND VPWR VPWR _096_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput40 chany_bottom_in[7] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input26_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_108_ _108_/A VGND VGND VPWR VPWR _108_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_14.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_20.mux_l1_in_1__A1 _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_3.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.mux_l2_in_1__157 VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/A0
+ mux_bottom_track_25.mux_l2_in_1__157/LO sky130_fd_sc_hd__conb_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput5 chanx_right_in[11] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_24.mux_l2_in_1_ mux_top_track_24.mux_l2_in_1_/A0 _125_/A mux_top_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_1__155 VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/A0
+ mux_bottom_track_1.mux_l2_in_1__155/LO sky130_fd_sc_hd__conb_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.mux_l1_in_0_ input19/X _097_/A mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input56_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_072_ _072_/A VGND VGND VPWR VPWR _072_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A mux_right_track_10.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_6.mux_l1_in_3__A1 _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_124_ _124_/A VGND VGND VPWR VPWR _124_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_12.mux_l3_in_0_ mux_right_track_12.mux_l2_in_1_/X mux_right_track_12.mux_l2_in_0_/X
+ mux_right_track_12.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_12.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xinput52 chany_top_in[18] VGND VGND VPWR VPWR _105_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput63 right_bottom_grid_pin_34_ VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__clkbuf_2
Xinput41 chany_bottom_in[8] VGND VGND VPWR VPWR _115_/A sky130_fd_sc_hd__clkbuf_2
Xinput30 chany_bottom_in[16] VGND VGND VPWR VPWR _123_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 input67/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input19_A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_107_ _107_/A VGND VGND VPWR VPWR _107_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_12.mux_l2_in_1_ mux_right_track_12.mux_l2_in_1_/A0 _117_/A mux_right_track_12.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_0.mux_l2_in_1_ mux_right_track_0.mux_l2_in_1_/A0 mux_right_track_0.mux_l1_in_2_/X
+ mux_right_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l1_in_2_ _109_/A input69/X mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__092__A _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 chanx_right_in[12] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_24.mux_l2_in_0_ _116_/A mux_top_track_24.mux_l1_in_0_/X mux_top_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_071_ _071_/A VGND VGND VPWR VPWR _071_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input49_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_123_ _123_/A VGND VGND VPWR VPWR _123_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_4.mux_l2_in_1__153 VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/A0
+ mux_top_track_4.mux_l2_in_1__153/LO sky130_fd_sc_hd__conb_1
Xinput31 chany_bottom_in[17] VGND VGND VPWR VPWR _124_/A sky130_fd_sc_hd__clkbuf_2
Xinput20 chanx_right_in[7] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_1
Xinput53 chany_top_in[19] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_1
Xinput64 right_bottom_grid_pin_35_ VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_2
Xinput42 chany_bottom_in[9] VGND VGND VPWR VPWR _116_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l2_in_1__138 VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/A0
+ mux_right_track_24.mux_l2_in_1__138/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 _100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_106_ _106_/A VGND VGND VPWR VPWR _106_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__095__A _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_12.mux_l2_in_0_ input65/X mux_right_track_12.mux_l1_in_0_/X mux_right_track_12.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input31_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_12.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_14.mux_l2_in_1__A1 _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_1_ input67/X input65/X mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_2.mux_l2_in_1_ mux_top_track_2.mux_l2_in_1_/A0 _120_/A mux_top_track_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_1_ mux_right_track_24.mux_l2_in_1_/A0 input33/X mux_right_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 chanx_right_in[13] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_070_ _070_/A VGND VGND VPWR VPWR _070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _118_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput130 _113_/X VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
XFILLER_15_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input61_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_122_ _122_/A VGND VGND VPWR VPWR _122_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_24.mux_l1_in_0_ input7/X input19/X mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput54 chany_top_in[1] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_1
Xinput43 chany_top_in[0] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
Xinput32 chany_bottom_in[18] VGND VGND VPWR VPWR _125_/A sky130_fd_sc_hd__clkbuf_2
Xinput21 chanx_right_in[8] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_1
Xinput10 chanx_right_in[16] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput65 right_bottom_grid_pin_36_ VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_105_ _105_/A VGND VGND VPWR VPWR _105_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input24_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _066_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_12.mux_l1_in_0_ input49/X _097_/A mux_right_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_0_ input63/X _089_/A mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _107_/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_24.mux_l2_in_0_ _125_/A mux_right_track_24.mux_l1_in_0_/X mux_right_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 input67/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput8 chanx_right_in[14] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_9.mux_l2_in_1__161 VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/A0
+ mux_bottom_track_9.mux_l2_in_1__161/LO sky130_fd_sc_hd__conb_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l1_in_1_ _111_/A input10/X mux_top_track_2.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput131 _114_/X VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
Xoutput120 _122_/X VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
X_121_ _121_/A VGND VGND VPWR VPWR _121_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input54_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xinput44 chany_top_in[10] VGND VGND VPWR VPWR _097_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput55 chany_top_in[2] VGND VGND VPWR VPWR _089_/A sky130_fd_sc_hd__clkbuf_2
Xinput66 right_bottom_grid_pin_37_ VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput33 chany_bottom_in[19] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
Xinput22 chanx_right_in[9] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput11 chanx_right_in[17] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_104_ _104_/A VGND VGND VPWR VPWR _104_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_1.mux_l2_in_1_ mux_bottom_track_1.mux_l2_in_1_/A0 mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input17_A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_12.sky130_fd_sc_hd__buf_4_0_ mux_right_track_12.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _072_/A sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l1_in_2_ input1/X input13/X mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input9_A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 chanx_right_in[15] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_18.mux_l1_in_1__A1 _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_2.mux_l1_in_0_ input22/X input15/X mux_top_track_2.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_0_ input63/X _105_/A mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput132 _115_/X VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
Xoutput121 _123_/X VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
Xoutput110 _093_/X VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_120_ _120_/A VGND VGND VPWR VPWR _120_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_36.mux_l2_in_0_ mux_right_track_36.mux_l2_in_0_/A0 mux_right_track_36.mux_l1_in_0_/X
+ mux_right_track_36.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_36.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input47_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_30.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xinput56 chany_top_in[3] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__clkbuf_1
Xinput45 chany_top_in[11] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_1
Xinput67 right_bottom_grid_pin_38_ VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 chany_bottom_in[0] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_1
Xinput34 chany_bottom_in[1] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_1
Xinput12 chanx_right_in[18] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_32.mux_l2_in_1__152 VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/A0
+ mux_top_track_32.mux_l2_in_1__152/LO sky130_fd_sc_hd__conb_1
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_103_ _103_/A VGND VGND VPWR VPWR _103_/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_1.mux_l1_in_1_ input6/X input18/X mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_34.sky130_fd_sc_hd__buf_4_0_ mux_right_track_34.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _083_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__101__A _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X input2/X VGND VGND
+ VPWR VPWR mux_top_track_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_28.sky130_fd_sc_hd__buf_4_0_ mux_right_track_28.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _080_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput122 _124_/X VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
Xoutput100 _102_/X VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
Xoutput111 _094_/X VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
Xmux_right_track_2.mux_l1_in_3__135 VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_3_/A0
+ mux_right_track_2.mux_l1_in_3__135/LO sky130_fd_sc_hd__conb_1
XFILLER_23_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 chanx_right_in[19] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
Xinput46 chany_top_in[12] VGND VGND VPWR VPWR _099_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput57 chany_top_in[4] VGND VGND VPWR VPWR _091_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput68 right_bottom_grid_pin_39_ VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput35 chany_bottom_in[2] VGND VGND VPWR VPWR _109_/A sky130_fd_sc_hd__clkbuf_2
Xinput24 chany_bottom_in[10] VGND VGND VPWR VPWR _117_/A sky130_fd_sc_hd__clkbuf_2
Xmux_top_track_2.mux_l2_in_1__150 VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/A0
+ mux_top_track_2.mux_l2_in_1__150/LO sky130_fd_sc_hd__conb_1
XFILLER_20_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _086_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_102_ _102_/A VGND VGND VPWR VPWR _102_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_36.mux_l1_in_0_ input23/X input69/X mux_right_track_36.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_36.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__104__A _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l1_in_0_ _099_/A _089_/A mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__112__A _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput123 _125_/X VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
Xoutput101 _103_/X VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xoutput112 _095_/X VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_6.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput14 chanx_right_in[1] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_1
Xinput36 chany_bottom_in[3] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__clkbuf_1
Xinput25 chany_bottom_in[11] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
Xinput58 chany_top_in[5] VGND VGND VPWR VPWR _092_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput47 chany_top_in[13] VGND VGND VPWR VPWR _100_/A sky130_fd_sc_hd__clkbuf_2
Xinput69 right_bottom_grid_pin_40_ VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_101_ _101_/A VGND VGND VPWR VPWR _101_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input52_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_26.mux_l2_in_0__139 VGND VGND VPWR VPWR mux_right_track_26.mux_l2_in_0_/A0
+ mux_right_track_26.mux_l2_in_0__139/LO sky130_fd_sc_hd__conb_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__120__A _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input15_A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__115__A _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_32.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_2
Xmux_top_track_16.mux_l2_in_1__149 VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/A0
+ mux_top_track_16.mux_l2_in_1__149/LO sky130_fd_sc_hd__conb_1
XANTENNA_input7_A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput124 _107_/X VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
Xoutput113 _106_/X VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
Xoutput102 _104_/X VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput59 chany_top_in[6] VGND VGND VPWR VPWR _093_/A sky130_fd_sc_hd__clkbuf_2
Xinput48 chany_top_in[14] VGND VGND VPWR VPWR _101_/A sky130_fd_sc_hd__clkbuf_2
Xinput37 chany_bottom_in[4] VGND VGND VPWR VPWR _111_/A sky130_fd_sc_hd__clkbuf_2
Xinput26 chany_bottom_in[12] VGND VGND VPWR VPWR _119_/A sky130_fd_sc_hd__clkbuf_2
Xinput15 chanx_right_in[2] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__123__A _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_100_ _100_/A VGND VGND VPWR VPWR _100_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input45_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 input65/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_6.mux_l1_in_3_ mux_right_track_6.mux_l1_in_3_/A0 _113_/A mux_right_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_32.mux_l2_in_1_ mux_top_track_32.mux_l2_in_1_/A0 _117_/A mux_top_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput114 _116_/X VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
Xoutput125 _108_/X VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
Xoutput103 _105_/X VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_2
XFILLER_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_6.mux_l3_in_0_ mux_right_track_6.mux_l2_in_1_/X mux_right_track_6.mux_l2_in_0_/X
+ mux_right_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput49 chany_top_in[15] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_1
Xinput38 chany_bottom_in[5] VGND VGND VPWR VPWR _112_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput27 chany_bottom_in[13] VGND VGND VPWR VPWR _120_/A sky130_fd_sc_hd__clkbuf_2
Xinput16 chanx_right_in[3] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input38_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_6.mux_l2_in_1_ mux_right_track_6.mux_l1_in_3_/X mux_right_track_6.mux_l1_in_2_/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l1_in_3__A1 _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_6.mux_l1_in_2_ _085_/A input68/X mux_right_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input20_A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l2_in_0_ input8/X mux_top_track_32.mux_l1_in_0_/X mux_top_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input68_A right_bottom_grid_pin_39_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_14 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput126 _109_/X VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
Xoutput115 _117_/X VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_22.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xoutput104 _087_/X VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
XFILLER_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput39 chany_bottom_in[6] VGND VGND VPWR VPWR _113_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput28 chany_bottom_in[14] VGND VGND VPWR VPWR _121_/A sky130_fd_sc_hd__clkbuf_2
Xinput17 chanx_right_in[4] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_089_ _089_/A VGND VGND VPWR VPWR _089_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_18.mux_l2_in_0_ mux_right_track_18.mux_l1_in_1_/X mux_right_track_18.mux_l1_in_0_/X
+ mux_right_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_18.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_0_ mux_right_track_6.mux_l1_in_1_/X mux_right_track_6.mux_l1_in_0_/X
+ mux_right_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_20.mux_l2_in_0_ mux_right_track_20.mux_l1_in_1_/X mux_right_track_20.mux_l1_in_0_/X
+ mux_right_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_20.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input50_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_18.mux_l1_in_1_ mux_right_track_18.mux_l1_in_1_/A0 _121_/A mux_right_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_6.mux_l1_in_1_ input66/X input64/X mux_right_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_8.mux_l2_in_1_ mux_top_track_8.mux_l2_in_1_/A0 mux_top_track_8.mux_l1_in_2_/X
+ mux_top_track_8.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_20.mux_l1_in_1_ mux_right_track_20.mux_l1_in_1_/A0 _123_/A mux_right_track_20.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_12.mux_l1_in_0__A1 _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input13_A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input5_A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_8.mux_l1_in_2_ _123_/A _113_/A mux_top_track_8.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput116 _118_/X VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
Xoutput127 _110_/X VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
Xoutput105 _088_/X VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l1_in_2__A0 _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 chanx_right_in[5] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 chany_bottom_in[15] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l1_in_0_ input20/X input3/X mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_10.mux_l2_in_1__A1 _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_088_ _088_/A VGND VGND VPWR VPWR _088_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input43_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_10.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_20.mux_l1_in_0__A1 _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_11 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_18.mux_l1_in_0_ input68/X _101_/A mux_right_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_36.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_6.mux_l1_in_0_ _093_/A input56/X mux_right_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _098_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_20.mux_l1_in_0_ input69/X _103_/A mux_right_track_20.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_20.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_6.sky130_fd_sc_hd__buf_4_0_ mux_right_track_6.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _069_/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l2_in_0_/A0 mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_1_ input12/X input5/X mux_top_track_8.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _110_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput128 _111_/X VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
Xoutput117 _119_/X VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
Xoutput106 _089_/X VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput19 chanx_right_in[6] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_30.sky130_fd_sc_hd__buf_4_0_ mux_right_track_30.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_087_ _087_/A VGND VGND VPWR VPWR _087_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input36_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_24.mux_l2_in_0__S mux_top_track_24.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_right_track_14.mux_l2_in_0__A0 input66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_18.sky130_fd_sc_hd__buf_4_0_ mux_right_track_18.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _075_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_8.mux_l1_in_0_ input17/X input71/X mux_top_track_8.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput107 _090_/X VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
Xoutput129 _112_/X VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
Xoutput118 _120_/X VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
Xmux_right_track_32.mux_l1_in_0_ input36/X input67/X mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input66_A right_bottom_grid_pin_37_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ _086_/A VGND VGND VPWR VPWR _086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__085__A _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input29_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_8.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_10.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_069_ _069_/A VGND VGND VPWR VPWR _069_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__093__A _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input11_A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput119 _121_/X VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
Xoutput108 _091_/X VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xoutput90 _073_/X VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input3_A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input59_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_22.mux_l1_in_1__A1 _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_085_ _085_/A VGND VGND VPWR VPWR _085_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_068_ _068_/A VGND VGND VPWR VPWR _068_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__096__A _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input41_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l2_in_1__156 VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/A0
+ mux_bottom_track_17.mux_l2_in_1__156/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_14.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput109 _092_/X VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
Xoutput80 _082_/X VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
XANTENNA_output72_A output72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput91 _074_/X VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
Xmux_right_track_36.mux_l2_in_0__144 VGND VGND VPWR VPWR mux_right_track_36.mux_l2_in_0_/A0
+ mux_right_track_36.mux_l2_in_0__144/LO sky130_fd_sc_hd__conb_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_24.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_18.mux_l1_in_1__134 VGND VGND VPWR VPWR mux_right_track_18.mux_l1_in_1_/A0
+ mux_right_track_18.mux_l1_in_1__134/LO sky130_fd_sc_hd__conb_1
XFILLER_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__099__A _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input71_A top_left_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_084_ _084_/A VGND VGND VPWR VPWR _084_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l1_in_3_ mux_right_track_2.mux_l1_in_3_/A0 _111_/A mux_right_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_067_ _067_/A VGND VGND VPWR VPWR _067_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input34_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_119_ _119_/A VGND VGND VPWR VPWR _119_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_14.mux_l3_in_0_ mux_right_track_14.mux_l2_in_1_/X mux_right_track_14.mux_l2_in_0_/X
+ mux_right_track_14.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_14.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_18.mux_l1_in_0__A1 _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput92 _075_/X VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
Xmux_right_track_14.mux_l2_in_1_ mux_right_track_14.mux_l2_in_1_/A0 _119_/A mux_right_track_14.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xoutput81 _083_/X VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ mux_right_track_2.mux_l1_in_3_/X mux_right_track_2.mux_l1_in_2_/X
+ mux_right_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_083_ _083_/A VGND VGND VPWR VPWR _083_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input64_A right_bottom_grid_pin_35_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_2.mux_l1_in_2_ _085_/A input68/X mux_right_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_066_ _066_/A VGND VGND VPWR VPWR _066_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_34.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_34.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input27_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_118_ _118_/A VGND VGND VPWR VPWR _118_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_26.mux_l1_in_0__A1 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_1__160 VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/A0
+ mux_bottom_track_5.mux_l2_in_1__160/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR output72/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_22.mux_l1_in_1__137 VGND VGND VPWR VPWR mux_right_track_22.mux_l1_in_1_/A0
+ mux_right_track_22.mux_l1_in_1__137/LO sky130_fd_sc_hd__conb_1
XFILLER_17_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 input67/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput82 _084_/X VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
Xoutput93 _086_/X VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
Xmux_right_track_14.mux_l2_in_0_ input66/X mux_right_track_14.mux_l1_in_0_/X mux_right_track_14.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_8.mux_l1_in_2__A0 _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input1_A bottom_left_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l2_in_1__A1 _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_082_ _082_/A VGND VGND VPWR VPWR _082_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input57_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l1_in_1_ input66/X input64/X mux_right_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l2_in_1_/A0 mux_top_track_4.mux_l1_in_2_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _122_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A mux_right_track_36.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_34.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l1_in_2_ _121_/A _112_/A mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_117_ _117_/A VGND VGND VPWR VPWR _117_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 input65/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput83 _085_/X VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
Xoutput72 output72/A VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_2
Xoutput94 _096_/X VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_8.mux_l1_in_2__A1 _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _067_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_14.mux_l1_in_0_ input53/X _099_/A mux_right_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_081_ _081_/A VGND VGND VPWR VPWR _081_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_2.mux_l1_in_0_ _091_/A input43/X mux_right_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_26.mux_l2_in_0_ mux_right_track_26.mux_l2_in_0_/A0 mux_right_track_26.mux_l1_in_0_/X
+ mux_right_track_26.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_26.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _108_/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_14.mux_l2_in_1__165 VGND VGND VPWR VPWR mux_right_track_14.mux_l2_in_1_/A0
+ mux_right_track_14.mux_l2_in_1__165/LO sky130_fd_sc_hd__conb_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_17.mux_l2_in_1_ mux_bottom_track_17.mux_l2_in_1_/A0 input9/X mux_bottom_track_17.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l1_in_1_ input11/X input4/X mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_116_ _116_/A VGND VGND VPWR VPWR _116_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__105__A _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input32_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_32.mux_l2_in_1__A1 _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l2_in_1_ mux_bottom_track_3.mux_l2_in_1_/A0 input12/X mux_bottom_track_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_20.sky130_fd_sc_hd__buf_4_0_ mux_right_track_20.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _076_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput95 _097_/X VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xoutput73 _066_/X VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
Xoutput84 _067_/X VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__113__A _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_14.sky130_fd_sc_hd__buf_4_0_ mux_right_track_14.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_080_ _080_/A VGND VGND VPWR VPWR _080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l2_in_1__151 VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/A0
+ mux_top_track_24.mux_l2_in_1__151/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input62_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l1_in_2__A0 _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_0_ input16/X input71/X mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_26.mux_l1_in_0_ input29/X input64/X mux_right_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_26.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_115_ _115_/A VGND VGND VPWR VPWR _115_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__121__A _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_1_ input21/X input14/X mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input25_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__S mux_bottom_track_3.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__116__A _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_33.mux_l2_in_0__S output72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_16.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput74 _076_/X VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
Xoutput96 _098_/X VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
Xoutput85 _068_/X VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

