magic
tech sky130A
magscale 1 2
timestamp 1625784544
<< locali >>
rect 3709 18615 3743 18717
rect 22017 16643 22051 17697
rect 9321 13243 9355 13481
rect 2697 12155 2731 12393
rect 22017 11339 22051 12257
rect 8953 10999 8987 11237
rect 6285 9503 6319 9605
rect 18613 8823 18647 9061
rect 9689 6647 9723 6885
rect 22017 5831 22051 6409
rect 6745 5151 6779 5321
rect 11989 4471 12023 4709
rect 22017 2839 22051 3961
rect 6687 1853 6837 1887
<< viali >>
rect 1869 20553 1903 20587
rect 2237 20553 2271 20587
rect 2605 20553 2639 20587
rect 7297 20553 7331 20587
rect 19073 20553 19107 20587
rect 19625 20553 19659 20587
rect 2881 20485 2915 20519
rect 4537 20485 4571 20519
rect 10885 20485 10919 20519
rect 11253 20485 11287 20519
rect 11897 20485 11931 20519
rect 12265 20485 12299 20519
rect 12633 20485 12667 20519
rect 13001 20485 13035 20519
rect 13369 20485 13403 20519
rect 13737 20485 13771 20519
rect 14105 20485 14139 20519
rect 14749 20485 14783 20519
rect 15117 20485 15151 20519
rect 15485 20485 15519 20519
rect 15853 20485 15887 20519
rect 16313 20485 16347 20519
rect 16681 20485 16715 20519
rect 17233 20485 17267 20519
rect 17601 20485 17635 20519
rect 17969 20485 18003 20519
rect 18613 20485 18647 20519
rect 20453 20485 20487 20519
rect 20821 20485 20855 20519
rect 3525 20417 3559 20451
rect 5917 20417 5951 20451
rect 6653 20417 6687 20451
rect 21189 20417 21223 20451
rect 3065 20349 3099 20383
rect 3341 20349 3375 20383
rect 3617 20349 3651 20383
rect 3985 20349 4019 20383
rect 4629 20349 4663 20383
rect 4905 20349 4939 20383
rect 5365 20349 5399 20383
rect 5549 20349 5583 20383
rect 5733 20349 5767 20383
rect 6193 20349 6227 20383
rect 6377 20349 6411 20383
rect 7573 20349 7607 20383
rect 8033 20349 8067 20383
rect 8217 20349 8251 20383
rect 8401 20349 8435 20383
rect 8769 20349 8803 20383
rect 9229 20349 9263 20383
rect 9597 20349 9631 20383
rect 9965 20349 9999 20383
rect 10333 20349 10367 20383
rect 10701 20349 10735 20383
rect 18337 20349 18371 20383
rect 19165 20349 19199 20383
rect 19901 20349 19935 20383
rect 20269 20349 20303 20383
rect 20620 20349 20654 20383
rect 21005 20349 21039 20383
rect 1593 20281 1627 20315
rect 1961 20281 1995 20315
rect 2329 20281 2363 20315
rect 2697 20281 2731 20315
rect 4353 20281 4387 20315
rect 5089 20281 5123 20315
rect 6929 20281 6963 20315
rect 8953 20281 8987 20315
rect 11069 20281 11103 20315
rect 11437 20281 11471 20315
rect 12081 20281 12115 20315
rect 12449 20281 12483 20315
rect 12817 20281 12851 20315
rect 13185 20281 13219 20315
rect 13553 20281 13587 20315
rect 13921 20281 13955 20315
rect 14289 20281 14323 20315
rect 14933 20281 14967 20315
rect 15301 20281 15335 20315
rect 15669 20281 15703 20315
rect 16037 20281 16071 20315
rect 16497 20281 16531 20315
rect 16865 20281 16899 20315
rect 17417 20281 17451 20315
rect 17785 20281 17819 20315
rect 18153 20281 18187 20315
rect 18797 20281 18831 20315
rect 19533 20281 19567 20315
rect 21373 20281 21407 20315
rect 21557 20281 21591 20315
rect 1501 20213 1535 20247
rect 4077 20213 4111 20247
rect 5273 20213 5307 20247
rect 6837 20213 6871 20247
rect 7481 20213 7515 20247
rect 7941 20213 7975 20247
rect 8677 20213 8711 20247
rect 9505 20213 9539 20247
rect 9873 20213 9907 20247
rect 10241 20213 10275 20247
rect 10517 20213 10551 20247
rect 18521 20213 18555 20247
rect 20085 20213 20119 20247
rect 1869 20009 1903 20043
rect 5641 20009 5675 20043
rect 8125 20009 8159 20043
rect 9321 20009 9355 20043
rect 9781 20009 9815 20043
rect 10517 20009 10551 20043
rect 11621 20009 11655 20043
rect 16773 20009 16807 20043
rect 16957 20009 16991 20043
rect 17233 20009 17267 20043
rect 18337 20009 18371 20043
rect 1593 19941 1627 19975
rect 7389 19941 7423 19975
rect 9137 19941 9171 19975
rect 11345 19941 11379 19975
rect 14381 19941 14415 19975
rect 20085 19941 20119 19975
rect 20453 19941 20487 19975
rect 20637 19941 20671 19975
rect 20913 19941 20947 19975
rect 1961 19873 1995 19907
rect 2145 19873 2179 19907
rect 2421 19873 2455 19907
rect 2697 19873 2731 19907
rect 2965 19873 2999 19907
rect 3249 19873 3283 19907
rect 3525 19873 3559 19907
rect 5109 19873 5143 19907
rect 5457 19873 5491 19907
rect 6092 19873 6126 19907
rect 8033 19873 8067 19907
rect 8677 19873 8711 19907
rect 8769 19873 8803 19907
rect 10149 19873 10183 19907
rect 10333 19873 10367 19907
rect 10793 19873 10827 19907
rect 11437 19873 11471 19907
rect 12173 19873 12207 19907
rect 14565 19873 14599 19907
rect 17049 19873 17083 19907
rect 17325 19873 17359 19907
rect 17601 19873 17635 19907
rect 17877 19873 17911 19907
rect 18153 19873 18187 19907
rect 18613 19873 18647 19907
rect 19165 19873 19199 19907
rect 19257 19873 19291 19907
rect 19717 19873 19751 19907
rect 21189 19873 21223 19907
rect 21373 19873 21407 19907
rect 5365 19805 5399 19839
rect 5825 19805 5859 19839
rect 8217 19805 8251 19839
rect 18889 19805 18923 19839
rect 19901 19805 19935 19839
rect 20269 19805 20303 19839
rect 2329 19737 2363 19771
rect 2605 19737 2639 19771
rect 11069 19737 11103 19771
rect 17509 19737 17543 19771
rect 18429 19737 18463 19771
rect 19441 19737 19475 19771
rect 1501 19669 1535 19703
rect 2881 19669 2915 19703
rect 3157 19669 3191 19703
rect 3433 19669 3467 19703
rect 3709 19669 3743 19703
rect 3985 19669 4019 19703
rect 7205 19669 7239 19703
rect 7481 19669 7515 19703
rect 7665 19669 7699 19703
rect 8493 19669 8527 19703
rect 10609 19669 10643 19703
rect 10885 19669 10919 19703
rect 11805 19669 11839 19703
rect 12357 19669 12391 19703
rect 17785 19669 17819 19703
rect 18061 19669 18095 19703
rect 21465 19669 21499 19703
rect 1777 19465 1811 19499
rect 3157 19465 3191 19499
rect 3709 19465 3743 19499
rect 3985 19465 4019 19499
rect 6837 19465 6871 19499
rect 10149 19465 10183 19499
rect 11437 19465 11471 19499
rect 12541 19465 12575 19499
rect 13001 19465 13035 19499
rect 13277 19465 13311 19499
rect 13829 19465 13863 19499
rect 14565 19465 14599 19499
rect 15761 19465 15795 19499
rect 16681 19465 16715 19499
rect 17417 19465 17451 19499
rect 18061 19465 18095 19499
rect 21373 19465 21407 19499
rect 6469 19397 6503 19431
rect 15301 19397 15335 19431
rect 18245 19397 18279 19431
rect 9045 19329 9079 19363
rect 10977 19329 11011 19363
rect 11897 19329 11931 19363
rect 21005 19329 21039 19363
rect 1409 19261 1443 19295
rect 1961 19261 1995 19295
rect 2053 19261 2087 19295
rect 2329 19261 2363 19295
rect 2789 19261 2823 19295
rect 2881 19261 2915 19295
rect 3341 19261 3375 19295
rect 3801 19261 3835 19295
rect 5282 19261 5316 19295
rect 5549 19261 5583 19295
rect 5917 19261 5951 19295
rect 6653 19261 6687 19295
rect 8401 19261 8435 19295
rect 9321 19261 9355 19295
rect 9689 19261 9723 19295
rect 9965 19261 9999 19295
rect 11253 19261 11287 19295
rect 12725 19261 12759 19295
rect 12817 19261 12851 19295
rect 13093 19261 13127 19295
rect 13369 19261 13403 19295
rect 13645 19261 13679 19295
rect 14289 19261 14323 19295
rect 14381 19261 14415 19295
rect 14841 19261 14875 19295
rect 15117 19261 15151 19295
rect 15393 19261 15427 19295
rect 15577 19261 15611 19295
rect 16129 19261 16163 19295
rect 16497 19261 16531 19295
rect 17233 19261 17267 19295
rect 17601 19261 17635 19295
rect 17877 19261 17911 19295
rect 18521 19261 18555 19295
rect 18889 19261 18923 19295
rect 20821 19261 20855 19295
rect 21557 19261 21591 19295
rect 1593 19193 1627 19227
rect 5641 19193 5675 19227
rect 6193 19193 6227 19227
rect 8134 19193 8168 19227
rect 8861 19193 8895 19227
rect 10793 19193 10827 19227
rect 16221 19193 16255 19227
rect 18337 19193 18371 19227
rect 18981 19193 19015 19227
rect 2237 19125 2271 19159
rect 2513 19125 2547 19159
rect 2605 19125 2639 19159
rect 3065 19125 3099 19159
rect 4169 19125 4203 19159
rect 6101 19125 6135 19159
rect 7021 19125 7055 19159
rect 8493 19125 8527 19159
rect 8953 19125 8987 19159
rect 9505 19125 9539 19159
rect 9873 19125 9907 19159
rect 10425 19125 10459 19159
rect 10885 19125 10919 19159
rect 11989 19125 12023 19159
rect 12081 19125 12115 19159
rect 12449 19125 12483 19159
rect 13553 19125 13587 19159
rect 14013 19125 14047 19159
rect 14749 19125 14783 19159
rect 15025 19125 15059 19159
rect 15945 19125 15979 19159
rect 17049 19125 17083 19159
rect 17785 19125 17819 19159
rect 18705 19125 18739 19159
rect 20269 19125 20303 19159
rect 1777 18921 1811 18955
rect 2053 18921 2087 18955
rect 2329 18921 2363 18955
rect 2973 18921 3007 18955
rect 3525 18921 3559 18955
rect 4813 18921 4847 18955
rect 5365 18921 5399 18955
rect 7113 18921 7147 18955
rect 7665 18921 7699 18955
rect 8033 18921 8067 18955
rect 8585 18921 8619 18955
rect 10149 18921 10183 18955
rect 10517 18921 10551 18955
rect 11989 18921 12023 18955
rect 12725 18921 12759 18955
rect 14381 18921 14415 18955
rect 18153 18921 18187 18955
rect 18429 18921 18463 18955
rect 19257 18921 19291 18955
rect 19717 18921 19751 18955
rect 20177 18921 20211 18955
rect 20729 18921 20763 18955
rect 1409 18853 1443 18887
rect 1593 18853 1627 18887
rect 2605 18853 2639 18887
rect 3341 18853 3375 18887
rect 4905 18853 4939 18887
rect 21189 18853 21223 18887
rect 1961 18785 1995 18819
rect 2237 18785 2271 18819
rect 2513 18785 2547 18819
rect 3157 18785 3191 18819
rect 4353 18785 4387 18819
rect 6478 18785 6512 18819
rect 8493 18785 8527 18819
rect 10876 18785 10910 18819
rect 12357 18785 12391 18819
rect 14565 18785 14599 18819
rect 14657 18785 14691 18819
rect 18889 18785 18923 18819
rect 19165 18785 19199 18819
rect 19441 18785 19475 18819
rect 19901 18785 19935 18819
rect 19993 18785 20027 18819
rect 20453 18785 20487 18819
rect 20637 18785 20671 18819
rect 21005 18785 21039 18819
rect 21373 18785 21407 18819
rect 21557 18785 21591 18819
rect 3709 18717 3743 18751
rect 5089 18717 5123 18751
rect 6745 18717 6779 18751
rect 6837 18717 6871 18751
rect 7389 18717 7423 18751
rect 7573 18717 7607 18751
rect 8677 18717 8711 18751
rect 9873 18717 9907 18751
rect 10057 18717 10091 18751
rect 10609 18717 10643 18751
rect 17509 18717 17543 18751
rect 2789 18649 2823 18683
rect 3985 18649 4019 18683
rect 4445 18649 4479 18683
rect 8125 18649 8159 18683
rect 17693 18649 17727 18683
rect 18705 18649 18739 18683
rect 18981 18649 19015 18683
rect 20269 18649 20303 18683
rect 3709 18581 3743 18615
rect 4169 18581 4203 18615
rect 12909 18581 12943 18615
rect 17049 18581 17083 18615
rect 17969 18581 18003 18615
rect 1869 18377 1903 18411
rect 2697 18377 2731 18411
rect 5457 18377 5491 18411
rect 8217 18377 8251 18411
rect 14657 18377 14691 18411
rect 16589 18377 16623 18411
rect 19349 18377 19383 18411
rect 19625 18377 19659 18411
rect 19901 18377 19935 18411
rect 20269 18377 20303 18411
rect 2145 18309 2179 18343
rect 10885 18309 10919 18343
rect 16037 18309 16071 18343
rect 19073 18309 19107 18343
rect 20545 18309 20579 18343
rect 21189 18309 21223 18343
rect 3617 18241 3651 18275
rect 3801 18241 3835 18275
rect 4445 18241 4479 18275
rect 4537 18241 4571 18275
rect 5733 18241 5767 18275
rect 7021 18241 7055 18275
rect 7573 18241 7607 18275
rect 8493 18241 8527 18275
rect 1593 18173 1627 18207
rect 2329 18173 2363 18207
rect 2605 18173 2639 18207
rect 2881 18173 2915 18207
rect 5917 18173 5951 18207
rect 6837 18173 6871 18207
rect 7849 18173 7883 18207
rect 8677 18173 8711 18207
rect 9505 18173 9539 18207
rect 11713 18173 11747 18207
rect 14473 18173 14507 18207
rect 15853 18173 15887 18207
rect 16405 18173 16439 18207
rect 18797 18173 18831 18207
rect 18889 18173 18923 18207
rect 19717 18173 19751 18207
rect 20085 18173 20119 18207
rect 20361 18173 20395 18207
rect 20637 18173 20671 18207
rect 21373 18173 21407 18207
rect 1961 18105 1995 18139
rect 9772 18105 9806 18139
rect 11958 18105 11992 18139
rect 21005 18105 21039 18139
rect 21557 18105 21591 18139
rect 1501 18037 1535 18071
rect 2421 18037 2455 18071
rect 2973 18037 3007 18071
rect 3157 18037 3191 18071
rect 3525 18037 3559 18071
rect 3985 18037 4019 18071
rect 4353 18037 4387 18071
rect 5825 18037 5859 18071
rect 6285 18037 6319 18071
rect 6469 18037 6503 18071
rect 6929 18037 6963 18071
rect 7757 18037 7791 18071
rect 8585 18037 8619 18071
rect 9045 18037 9079 18071
rect 10977 18037 11011 18071
rect 13093 18037 13127 18071
rect 20821 18037 20855 18071
rect 2605 17833 2639 17867
rect 3341 17833 3375 17867
rect 4077 17833 4111 17867
rect 4445 17833 4479 17867
rect 4537 17833 4571 17867
rect 4905 17833 4939 17867
rect 5273 17833 5307 17867
rect 6377 17833 6411 17867
rect 6837 17833 6871 17867
rect 7021 17833 7055 17867
rect 7389 17833 7423 17867
rect 7849 17833 7883 17867
rect 8217 17833 8251 17867
rect 9137 17833 9171 17867
rect 9965 17833 9999 17867
rect 10425 17833 10459 17867
rect 10793 17833 10827 17867
rect 12357 17833 12391 17867
rect 13829 17833 13863 17867
rect 15117 17833 15151 17867
rect 15485 17833 15519 17867
rect 15945 17833 15979 17867
rect 16497 17833 16531 17867
rect 19441 17833 19475 17867
rect 20361 17833 20395 17867
rect 20637 17833 20671 17867
rect 1593 17765 1627 17799
rect 3433 17765 3467 17799
rect 11161 17765 11195 17799
rect 14749 17765 14783 17799
rect 19809 17765 19843 17799
rect 1961 17697 1995 17731
rect 2513 17697 2547 17731
rect 6469 17697 6503 17731
rect 7481 17697 7515 17731
rect 9873 17697 9907 17731
rect 10333 17697 10367 17731
rect 11989 17697 12023 17731
rect 13185 17697 13219 17731
rect 13645 17697 13679 17731
rect 15577 17697 15611 17731
rect 16405 17697 16439 17731
rect 19901 17697 19935 17731
rect 20177 17697 20211 17731
rect 20453 17697 20487 17731
rect 21189 17697 21223 17731
rect 21373 17697 21407 17731
rect 22017 17697 22051 17731
rect 2697 17629 2731 17663
rect 3525 17629 3559 17663
rect 3985 17629 4019 17663
rect 4721 17629 4755 17663
rect 5365 17629 5399 17663
rect 5457 17629 5491 17663
rect 6193 17629 6227 17663
rect 7573 17629 7607 17663
rect 8309 17629 8343 17663
rect 8401 17629 8435 17663
rect 8953 17629 8987 17663
rect 10609 17629 10643 17663
rect 11253 17629 11287 17663
rect 11345 17629 11379 17663
rect 11713 17629 11747 17663
rect 11897 17629 11931 17663
rect 12909 17629 12943 17663
rect 13093 17629 13127 17663
rect 14565 17629 14599 17663
rect 14657 17629 14691 17663
rect 15393 17629 15427 17663
rect 16681 17629 16715 17663
rect 21005 17629 21039 17663
rect 1777 17561 1811 17595
rect 12449 17561 12483 17595
rect 13553 17561 13587 17595
rect 16037 17561 16071 17595
rect 21557 17561 21591 17595
rect 1501 17493 1535 17527
rect 2145 17493 2179 17527
rect 2973 17493 3007 17527
rect 6009 17493 6043 17527
rect 8677 17493 8711 17527
rect 20085 17493 20119 17527
rect 4077 17289 4111 17323
rect 7941 17289 7975 17323
rect 11253 17289 11287 17323
rect 13829 17289 13863 17323
rect 16773 17289 16807 17323
rect 21005 17289 21039 17323
rect 2605 17221 2639 17255
rect 4169 17221 4203 17255
rect 7849 17221 7883 17255
rect 10149 17221 10183 17255
rect 20729 17221 20763 17255
rect 2053 17153 2087 17187
rect 2145 17153 2179 17187
rect 4629 17153 4663 17187
rect 4813 17153 4847 17187
rect 5457 17153 5491 17187
rect 6469 17153 6503 17187
rect 8493 17153 8527 17187
rect 8769 17153 8803 17187
rect 10609 17153 10643 17187
rect 12449 17153 12483 17187
rect 21097 17153 21131 17187
rect 21557 17153 21591 17187
rect 1593 17085 1627 17119
rect 2237 17085 2271 17119
rect 2697 17085 2731 17119
rect 5549 17085 5583 17119
rect 8309 17085 8343 17119
rect 9025 17085 9059 17119
rect 10885 17085 10919 17119
rect 13921 17085 13955 17119
rect 14177 17085 14211 17119
rect 15393 17085 15427 17119
rect 20545 17085 20579 17119
rect 20821 17085 20855 17119
rect 2942 17017 2976 17051
rect 4537 17017 4571 17051
rect 4997 17017 5031 17051
rect 6736 17017 6770 17051
rect 12716 17017 12750 17051
rect 15660 17017 15694 17051
rect 21373 17017 21407 17051
rect 1501 16949 1535 16983
rect 5641 16949 5675 16983
rect 6009 16949 6043 16983
rect 8401 16949 8435 16983
rect 10425 16949 10459 16983
rect 10793 16949 10827 16983
rect 11713 16949 11747 16983
rect 15301 16949 15335 16983
rect 19993 16949 20027 16983
rect 20361 16949 20395 16983
rect 1777 16745 1811 16779
rect 3525 16745 3559 16779
rect 3985 16745 4019 16779
rect 7389 16745 7423 16779
rect 9137 16745 9171 16779
rect 9781 16745 9815 16779
rect 10241 16745 10275 16779
rect 10609 16745 10643 16779
rect 11161 16745 11195 16779
rect 11805 16745 11839 16779
rect 12265 16745 12299 16779
rect 12633 16745 12667 16779
rect 13093 16745 13127 16779
rect 13645 16745 13679 16779
rect 15761 16745 15795 16779
rect 16037 16745 16071 16779
rect 20177 16745 20211 16779
rect 21005 16745 21039 16779
rect 1593 16677 1627 16711
rect 4344 16677 4378 16711
rect 8502 16677 8536 16711
rect 11069 16677 11103 16711
rect 14648 16677 14682 16711
rect 17150 16677 17184 16711
rect 20361 16677 20395 16711
rect 21373 16677 21407 16711
rect 21557 16677 21591 16711
rect 2890 16609 2924 16643
rect 3433 16609 3467 16643
rect 3709 16609 3743 16643
rect 5549 16609 5583 16643
rect 5805 16609 5839 16643
rect 11897 16609 11931 16643
rect 12725 16609 12759 16643
rect 13553 16609 13587 16643
rect 14381 16609 14415 16643
rect 17417 16609 17451 16643
rect 19993 16609 20027 16643
rect 20545 16609 20579 16643
rect 20821 16609 20855 16643
rect 22017 16609 22051 16643
rect 3157 16541 3191 16575
rect 4077 16541 4111 16575
rect 8769 16541 8803 16575
rect 10057 16541 10091 16575
rect 10149 16541 10183 16575
rect 11253 16541 11287 16575
rect 11713 16541 11747 16575
rect 12449 16541 12483 16575
rect 13737 16541 13771 16575
rect 3249 16473 3283 16507
rect 8953 16473 8987 16507
rect 10701 16473 10735 16507
rect 13185 16473 13219 16507
rect 20729 16473 20763 16507
rect 1501 16405 1535 16439
rect 5457 16405 5491 16439
rect 6929 16405 6963 16439
rect 14013 16405 14047 16439
rect 21097 16405 21131 16439
rect 2329 16201 2363 16235
rect 3249 16201 3283 16235
rect 3525 16201 3559 16235
rect 4721 16201 4755 16235
rect 8953 16201 8987 16235
rect 9689 16201 9723 16235
rect 13277 16201 13311 16235
rect 14197 16201 14231 16235
rect 15301 16201 15335 16235
rect 20821 16201 20855 16235
rect 3801 16133 3835 16167
rect 7297 16133 7331 16167
rect 21557 16133 21591 16167
rect 1777 16065 1811 16099
rect 1869 16065 1903 16099
rect 3065 16065 3099 16099
rect 4353 16065 4387 16099
rect 5365 16065 5399 16099
rect 5549 16065 5583 16099
rect 6745 16065 6779 16099
rect 7481 16065 7515 16099
rect 8401 16065 8435 16099
rect 8493 16065 8527 16099
rect 11897 16065 11931 16099
rect 13461 16065 13495 16099
rect 14749 16065 14783 16099
rect 15853 16065 15887 16099
rect 3433 15997 3467 16031
rect 3709 15997 3743 16031
rect 11069 15997 11103 16031
rect 12164 15997 12198 16031
rect 13645 15997 13679 16031
rect 20637 15997 20671 16031
rect 1961 15929 1995 15963
rect 2881 15929 2915 15963
rect 4169 15929 4203 15963
rect 5641 15929 5675 15963
rect 6193 15929 6227 15963
rect 7665 15929 7699 15963
rect 8585 15929 8619 15963
rect 10802 15929 10836 15963
rect 14565 15929 14599 15963
rect 15669 15929 15703 15963
rect 21005 15929 21039 15963
rect 21189 15929 21223 15963
rect 21373 15929 21407 15963
rect 2421 15861 2455 15895
rect 2789 15861 2823 15895
rect 4261 15861 4295 15895
rect 5181 15861 5215 15895
rect 6009 15861 6043 15895
rect 6837 15861 6871 15895
rect 6929 15861 6963 15895
rect 7757 15861 7791 15895
rect 8125 15861 8159 15895
rect 11713 15861 11747 15895
rect 13737 15861 13771 15895
rect 14105 15861 14139 15895
rect 14657 15861 14691 15895
rect 15761 15861 15795 15895
rect 16129 15861 16163 15895
rect 16405 15861 16439 15895
rect 1869 15657 1903 15691
rect 2329 15657 2363 15691
rect 3893 15657 3927 15691
rect 4445 15657 4479 15691
rect 5641 15657 5675 15691
rect 6469 15657 6503 15691
rect 7665 15657 7699 15691
rect 11345 15657 11379 15691
rect 12633 15657 12667 15691
rect 13001 15657 13035 15691
rect 13921 15657 13955 15691
rect 14933 15657 14967 15691
rect 15761 15657 15795 15691
rect 20177 15657 20211 15691
rect 20453 15657 20487 15691
rect 20729 15657 20763 15691
rect 21005 15657 21039 15691
rect 4905 15589 4939 15623
rect 5549 15589 5583 15623
rect 6377 15589 6411 15623
rect 9404 15589 9438 15623
rect 19809 15589 19843 15623
rect 21373 15589 21407 15623
rect 1593 15521 1627 15555
rect 1961 15521 1995 15555
rect 3442 15521 3476 15555
rect 4077 15521 4111 15555
rect 4813 15521 4847 15555
rect 7297 15521 7331 15555
rect 7757 15521 7791 15555
rect 9137 15521 9171 15555
rect 10977 15521 11011 15555
rect 12541 15521 12575 15555
rect 13461 15521 13495 15555
rect 15669 15521 15703 15555
rect 18245 15521 18279 15555
rect 19993 15521 20027 15555
rect 20269 15521 20303 15555
rect 20545 15521 20579 15555
rect 20821 15521 20855 15555
rect 3709 15453 3743 15487
rect 4997 15453 5031 15487
rect 5457 15453 5491 15487
rect 6193 15453 6227 15487
rect 7021 15453 7055 15487
rect 7205 15453 7239 15487
rect 10793 15453 10827 15487
rect 10885 15453 10919 15487
rect 11989 15453 12023 15487
rect 12449 15453 12483 15487
rect 13185 15453 13219 15487
rect 13369 15453 13403 15487
rect 14749 15453 14783 15487
rect 14841 15453 14875 15487
rect 15485 15453 15519 15487
rect 17969 15453 18003 15487
rect 18153 15453 18187 15487
rect 19717 15453 19751 15487
rect 1409 15385 1443 15419
rect 4261 15385 4295 15419
rect 6009 15385 6043 15419
rect 10517 15385 10551 15419
rect 13829 15385 13863 15419
rect 21557 15385 21591 15419
rect 2145 15317 2179 15351
rect 6837 15317 6871 15351
rect 11805 15317 11839 15351
rect 12081 15317 12115 15351
rect 14473 15317 14507 15351
rect 15301 15317 15335 15351
rect 16129 15317 16163 15351
rect 18613 15317 18647 15351
rect 21097 15317 21131 15351
rect 2329 15113 2363 15147
rect 2697 15113 2731 15147
rect 4077 15113 4111 15147
rect 6285 15113 6319 15147
rect 6837 15113 6871 15147
rect 9413 15113 9447 15147
rect 11253 15113 11287 15147
rect 13921 15113 13955 15147
rect 16405 15113 16439 15147
rect 20177 15113 20211 15147
rect 20453 15113 20487 15147
rect 2053 15045 2087 15079
rect 10333 15045 10367 15079
rect 14841 15045 14875 15079
rect 1409 14977 1443 15011
rect 3249 14977 3283 15011
rect 4629 14977 4663 15011
rect 7849 14977 7883 15011
rect 8861 14977 8895 15011
rect 9965 14977 9999 15011
rect 10149 14977 10183 15011
rect 10977 14977 11011 15011
rect 13277 14977 13311 15011
rect 13461 14977 13495 15011
rect 15485 14977 15519 15011
rect 15761 14977 15795 15011
rect 15945 14977 15979 15011
rect 17509 14977 17543 15011
rect 21557 14977 21591 15011
rect 1961 14909 1995 14943
rect 2237 14909 2271 14943
rect 2513 14909 2547 14943
rect 3065 14909 3099 14943
rect 4905 14909 4939 14943
rect 5172 14909 5206 14943
rect 8401 14909 8435 14943
rect 9045 14909 9079 14943
rect 10701 14909 10735 14943
rect 11713 14909 11747 14943
rect 11980 14909 12014 14943
rect 14565 14909 14599 14943
rect 16037 14909 16071 14943
rect 19993 14909 20027 14943
rect 20269 14909 20303 14943
rect 20821 14909 20855 14943
rect 1593 14841 1627 14875
rect 3157 14841 3191 14875
rect 7205 14841 7239 14875
rect 7665 14841 7699 14875
rect 11437 14841 11471 14875
rect 13553 14841 13587 14875
rect 15209 14841 15243 14875
rect 17754 14841 17788 14875
rect 21373 14841 21407 14875
rect 1777 14773 1811 14807
rect 3525 14773 3559 14807
rect 3801 14773 3835 14807
rect 4445 14773 4479 14807
rect 4537 14773 4571 14807
rect 7297 14773 7331 14807
rect 7757 14773 7791 14807
rect 8125 14773 8159 14807
rect 8585 14773 8619 14807
rect 8953 14773 8987 14807
rect 9505 14773 9539 14807
rect 9873 14773 9907 14807
rect 10793 14773 10827 14807
rect 13093 14773 13127 14807
rect 14013 14773 14047 14807
rect 14197 14773 14231 14807
rect 14381 14773 14415 14807
rect 15301 14773 15335 14807
rect 18889 14773 18923 14807
rect 20729 14773 20763 14807
rect 21005 14773 21039 14807
rect 1869 14569 1903 14603
rect 2145 14569 2179 14603
rect 2605 14569 2639 14603
rect 2973 14569 3007 14603
rect 6469 14569 6503 14603
rect 6745 14569 6779 14603
rect 7113 14569 7147 14603
rect 10977 14569 11011 14603
rect 12909 14569 12943 14603
rect 19625 14569 19659 14603
rect 20821 14569 20855 14603
rect 1961 14501 1995 14535
rect 3065 14501 3099 14535
rect 3433 14501 3467 14535
rect 5825 14501 5859 14535
rect 6377 14501 6411 14535
rect 7818 14501 7852 14535
rect 10272 14501 10306 14535
rect 12357 14501 12391 14535
rect 15494 14501 15528 14535
rect 17264 14501 17298 14535
rect 21005 14501 21039 14535
rect 21189 14501 21223 14535
rect 1593 14433 1627 14467
rect 2329 14433 2363 14467
rect 4261 14433 4295 14467
rect 5917 14433 5951 14467
rect 6653 14433 6687 14467
rect 11805 14433 11839 14467
rect 11897 14433 11931 14467
rect 13553 14433 13587 14467
rect 15761 14433 15795 14467
rect 17509 14433 17543 14467
rect 17601 14433 17635 14467
rect 17868 14433 17902 14467
rect 19993 14433 20027 14467
rect 20637 14433 20671 14467
rect 21373 14433 21407 14467
rect 3249 14365 3283 14399
rect 3709 14365 3743 14399
rect 4353 14365 4387 14399
rect 4537 14365 4571 14399
rect 6101 14365 6135 14399
rect 7205 14365 7239 14399
rect 7297 14365 7331 14399
rect 7573 14365 7607 14399
rect 10517 14365 10551 14399
rect 11069 14365 11103 14399
rect 11161 14365 11195 14399
rect 12081 14365 12115 14399
rect 12633 14365 12667 14399
rect 12817 14365 12851 14399
rect 19073 14365 19107 14399
rect 20085 14365 20119 14399
rect 20177 14365 20211 14399
rect 3893 14297 3927 14331
rect 5457 14297 5491 14331
rect 8953 14297 8987 14331
rect 10609 14297 10643 14331
rect 13277 14297 13311 14331
rect 21557 14297 21591 14331
rect 1501 14229 1535 14263
rect 2513 14229 2547 14263
rect 4997 14229 5031 14263
rect 5181 14229 5215 14263
rect 9137 14229 9171 14263
rect 11437 14229 11471 14263
rect 13369 14229 13403 14263
rect 14381 14229 14415 14263
rect 16129 14229 16163 14263
rect 18981 14229 19015 14263
rect 20545 14229 20579 14263
rect 2697 14025 2731 14059
rect 8033 14025 8067 14059
rect 10241 14025 10275 14059
rect 12541 14025 12575 14059
rect 16497 14025 16531 14059
rect 16957 14025 16991 14059
rect 18705 14025 18739 14059
rect 19533 14025 19567 14059
rect 21005 14025 21039 14059
rect 2145 13957 2179 13991
rect 2421 13957 2455 13991
rect 3249 13957 3283 13991
rect 5549 13957 5583 13991
rect 6469 13957 6503 13991
rect 11345 13957 11379 13991
rect 13553 13957 13587 13991
rect 20729 13957 20763 13991
rect 6009 13889 6043 13923
rect 6193 13889 6227 13923
rect 7021 13889 7055 13923
rect 7481 13889 7515 13923
rect 9597 13889 9631 13923
rect 10793 13889 10827 13923
rect 11897 13889 11931 13923
rect 12817 13889 12851 13923
rect 15117 13889 15151 13923
rect 17509 13889 17543 13923
rect 18153 13889 18187 13923
rect 18889 13889 18923 13923
rect 1409 13821 1443 13855
rect 1777 13821 1811 13855
rect 1961 13821 1995 13855
rect 2329 13821 2363 13855
rect 2605 13821 2639 13855
rect 2881 13821 2915 13855
rect 4905 13821 4939 13855
rect 5457 13821 5491 13855
rect 6929 13821 6963 13855
rect 7573 13821 7607 13855
rect 11161 13821 11195 13855
rect 14933 13821 14967 13855
rect 17417 13821 17451 13855
rect 17785 13821 17819 13855
rect 18245 13821 18279 13855
rect 19165 13821 19199 13855
rect 20821 13821 20855 13855
rect 21557 13821 21591 13855
rect 1593 13753 1627 13787
rect 4660 13753 4694 13787
rect 9781 13753 9815 13787
rect 10609 13753 10643 13787
rect 13093 13753 13127 13787
rect 14688 13753 14722 13787
rect 15362 13753 15396 13787
rect 16773 13753 16807 13787
rect 17325 13753 17359 13787
rect 18337 13753 18371 13787
rect 21373 13753 21407 13787
rect 2973 13685 3007 13719
rect 3525 13685 3559 13719
rect 5917 13685 5951 13719
rect 6837 13685 6871 13719
rect 7665 13685 7699 13719
rect 8217 13685 8251 13719
rect 9321 13685 9355 13719
rect 9689 13685 9723 13719
rect 10149 13685 10183 13719
rect 10701 13685 10735 13719
rect 11437 13685 11471 13719
rect 11989 13685 12023 13719
rect 12081 13685 12115 13719
rect 12449 13685 12483 13719
rect 13001 13685 13035 13719
rect 13461 13685 13495 13719
rect 19073 13685 19107 13719
rect 2145 13481 2179 13515
rect 2697 13481 2731 13515
rect 3341 13481 3375 13515
rect 3709 13481 3743 13515
rect 5273 13481 5307 13515
rect 5917 13481 5951 13515
rect 6377 13481 6411 13515
rect 8217 13481 8251 13515
rect 8585 13481 8619 13515
rect 9321 13481 9355 13515
rect 9689 13481 9723 13515
rect 10425 13481 10459 13515
rect 11989 13481 12023 13515
rect 12081 13481 12115 13515
rect 12541 13481 12575 13515
rect 12909 13481 12943 13515
rect 13461 13481 13495 13515
rect 13829 13481 13863 13515
rect 14565 13481 14599 13515
rect 15301 13481 15335 13515
rect 15761 13481 15795 13515
rect 15853 13481 15887 13515
rect 16221 13481 16255 13515
rect 16865 13481 16899 13515
rect 17325 13481 17359 13515
rect 17877 13481 17911 13515
rect 18889 13481 18923 13515
rect 20361 13481 20395 13515
rect 21005 13481 21039 13515
rect 1593 13413 1627 13447
rect 3249 13413 3283 13447
rect 5365 13413 5399 13447
rect 6990 13413 7024 13447
rect 1961 13345 1995 13379
rect 2329 13345 2363 13379
rect 2605 13345 2639 13379
rect 2881 13345 2915 13379
rect 3893 13345 3927 13379
rect 4160 13345 4194 13379
rect 6285 13345 6319 13379
rect 6745 13345 6779 13379
rect 9229 13345 9263 13379
rect 3157 13277 3191 13311
rect 5733 13277 5767 13311
rect 6469 13277 6503 13311
rect 8677 13277 8711 13311
rect 8769 13277 8803 13311
rect 9781 13413 9815 13447
rect 15393 13413 15427 13447
rect 18797 13413 18831 13447
rect 21373 13413 21407 13447
rect 10609 13345 10643 13379
rect 10876 13345 10910 13379
rect 12449 13345 12483 13379
rect 14381 13345 14415 13379
rect 16313 13345 16347 13379
rect 16681 13345 16715 13379
rect 17417 13345 17451 13379
rect 18245 13345 18279 13379
rect 19073 13345 19107 13379
rect 20545 13345 20579 13379
rect 20821 13345 20855 13379
rect 21557 13345 21591 13379
rect 9505 13277 9539 13311
rect 12633 13277 12667 13311
rect 13921 13277 13955 13311
rect 14105 13277 14139 13311
rect 14749 13277 14783 13311
rect 15209 13277 15243 13311
rect 16497 13277 16531 13311
rect 17233 13277 17267 13311
rect 18337 13277 18371 13311
rect 18521 13277 18555 13311
rect 2421 13209 2455 13243
rect 9321 13209 9355 13243
rect 10149 13209 10183 13243
rect 13277 13209 13311 13243
rect 19257 13209 19291 13243
rect 1501 13141 1535 13175
rect 1869 13141 1903 13175
rect 8125 13141 8159 13175
rect 14933 13141 14967 13175
rect 17785 13141 17819 13175
rect 20729 13141 20763 13175
rect 1961 12937 1995 12971
rect 3433 12937 3467 12971
rect 5825 12937 5859 12971
rect 6469 12937 6503 12971
rect 7757 12937 7791 12971
rect 9505 12937 9539 12971
rect 11529 12937 11563 12971
rect 13829 12937 13863 12971
rect 14105 12937 14139 12971
rect 15761 12937 15795 12971
rect 17785 12937 17819 12971
rect 19349 12937 19383 12971
rect 21005 12937 21039 12971
rect 19257 12869 19291 12903
rect 3801 12801 3835 12835
rect 6009 12801 6043 12835
rect 7021 12801 7055 12835
rect 7573 12801 7607 12835
rect 10609 12801 10643 12835
rect 10885 12801 10919 12835
rect 11713 12801 11747 12835
rect 13185 12801 13219 12835
rect 14749 12801 14783 12835
rect 15577 12801 15611 12835
rect 16221 12801 16255 12835
rect 16405 12801 16439 12835
rect 17233 12801 17267 12835
rect 19901 12801 19935 12835
rect 21557 12801 21591 12835
rect 1777 12733 1811 12767
rect 2053 12733 2087 12767
rect 3893 12733 3927 12767
rect 4445 12733 4479 12767
rect 6101 12733 6135 12767
rect 7941 12733 7975 12767
rect 9146 12733 9180 12767
rect 9413 12733 9447 12767
rect 10333 12733 10367 12767
rect 10517 12733 10551 12767
rect 11069 12733 11103 12767
rect 11161 12733 11195 12767
rect 17417 12733 17451 12767
rect 17877 12733 17911 12767
rect 18133 12733 18167 12767
rect 20821 12733 20855 12767
rect 1593 12665 1627 12699
rect 2298 12665 2332 12699
rect 4712 12665 4746 12699
rect 6837 12665 6871 12699
rect 9873 12665 9907 12699
rect 10149 12665 10183 12699
rect 11958 12665 11992 12699
rect 15301 12665 15335 12699
rect 15393 12665 15427 12699
rect 16129 12665 16163 12699
rect 19809 12665 19843 12699
rect 21373 12665 21407 12699
rect 1501 12597 1535 12631
rect 3985 12597 4019 12631
rect 4353 12597 4387 12631
rect 6929 12597 6963 12631
rect 7297 12597 7331 12631
rect 8033 12597 8067 12631
rect 9689 12597 9723 12631
rect 13093 12597 13127 12631
rect 13921 12597 13955 12631
rect 14473 12597 14507 12631
rect 14565 12597 14599 12631
rect 14933 12597 14967 12631
rect 16773 12597 16807 12631
rect 17325 12597 17359 12631
rect 19717 12597 19751 12631
rect 2605 12393 2639 12427
rect 2697 12393 2731 12427
rect 3617 12393 3651 12427
rect 3985 12393 4019 12427
rect 4353 12393 4387 12427
rect 7665 12393 7699 12427
rect 8217 12393 8251 12427
rect 8677 12393 8711 12427
rect 9137 12393 9171 12427
rect 9597 12393 9631 12427
rect 10057 12393 10091 12427
rect 10333 12393 10367 12427
rect 12633 12393 12667 12427
rect 16221 12393 16255 12427
rect 16589 12393 16623 12427
rect 19257 12393 19291 12427
rect 20177 12393 20211 12427
rect 1685 12325 1719 12359
rect 1501 12257 1535 12291
rect 2237 12257 2271 12291
rect 1961 12189 1995 12223
rect 2145 12189 2179 12223
rect 6684 12325 6718 12359
rect 8585 12325 8619 12359
rect 9505 12325 9539 12359
rect 11446 12325 11480 12359
rect 13062 12325 13096 12359
rect 14381 12325 14415 12359
rect 14565 12325 14599 12359
rect 14994 12325 15028 12359
rect 21189 12325 21223 12359
rect 3157 12257 3191 12291
rect 4813 12257 4847 12291
rect 6929 12257 6963 12291
rect 7113 12257 7147 12291
rect 7573 12257 7607 12291
rect 11713 12257 11747 12291
rect 12173 12257 12207 12291
rect 12817 12257 12851 12291
rect 17049 12257 17083 12291
rect 17509 12257 17543 12291
rect 17776 12257 17810 12291
rect 19993 12257 20027 12291
rect 21005 12257 21039 12291
rect 21373 12257 21407 12291
rect 22017 12257 22051 12291
rect 3249 12189 3283 12223
rect 3341 12189 3375 12223
rect 4629 12189 4663 12223
rect 4721 12189 4755 12223
rect 7849 12189 7883 12223
rect 8769 12189 8803 12223
rect 9689 12189 9723 12223
rect 10149 12189 10183 12223
rect 11989 12189 12023 12223
rect 12081 12189 12115 12223
rect 14749 12189 14783 12223
rect 16681 12189 16715 12223
rect 16773 12189 16807 12223
rect 2697 12121 2731 12155
rect 2789 12121 2823 12155
rect 5365 12121 5399 12155
rect 21557 12121 21591 12155
rect 5181 12053 5215 12087
rect 5549 12053 5583 12087
rect 7205 12053 7239 12087
rect 8033 12053 8067 12087
rect 12541 12053 12575 12087
rect 14197 12053 14231 12087
rect 16129 12053 16163 12087
rect 17325 12053 17359 12087
rect 18889 12053 18923 12087
rect 19073 12053 19107 12087
rect 20821 12053 20855 12087
rect 1501 11849 1535 11883
rect 2973 11849 3007 11883
rect 3249 11849 3283 11883
rect 3617 11849 3651 11883
rect 4445 11849 4479 11883
rect 5549 11849 5583 11883
rect 6469 11849 6503 11883
rect 8769 11849 8803 11883
rect 10701 11849 10735 11883
rect 13277 11849 13311 11883
rect 18429 11849 18463 11883
rect 19993 11849 20027 11883
rect 20269 11849 20303 11883
rect 20729 11849 20763 11883
rect 21005 11849 21039 11883
rect 11713 11781 11747 11815
rect 18337 11781 18371 11815
rect 21281 11781 21315 11815
rect 2881 11713 2915 11747
rect 4169 11713 4203 11747
rect 4997 11713 5031 11747
rect 6101 11713 6135 11747
rect 8125 11713 8159 11747
rect 9321 11713 9355 11747
rect 10149 11713 10183 11747
rect 10241 11713 10275 11747
rect 11345 11713 11379 11747
rect 12265 11713 12299 11747
rect 12725 11713 12759 11747
rect 12817 11713 12851 11747
rect 15117 11713 15151 11747
rect 16221 11713 16255 11747
rect 18889 11713 18923 11747
rect 19073 11713 19107 11747
rect 19441 11713 19475 11747
rect 21189 11713 21223 11747
rect 2614 11645 2648 11679
rect 3157 11645 3191 11679
rect 3433 11645 3467 11679
rect 4905 11645 4939 11679
rect 6009 11645 6043 11679
rect 7849 11645 7883 11679
rect 9229 11645 9263 11679
rect 9873 11645 9907 11679
rect 12173 11645 12207 11679
rect 14850 11645 14884 11679
rect 15393 11645 15427 11679
rect 15853 11645 15887 11679
rect 16957 11645 16991 11679
rect 18797 11645 18831 11679
rect 19625 11645 19659 11679
rect 20177 11645 20211 11679
rect 20453 11645 20487 11679
rect 20545 11645 20579 11679
rect 20821 11645 20855 11679
rect 3985 11577 4019 11611
rect 4813 11577 4847 11611
rect 7582 11577 7616 11611
rect 8217 11577 8251 11611
rect 10333 11577 10367 11611
rect 11253 11577 11287 11611
rect 12081 11577 12115 11611
rect 15577 11577 15611 11611
rect 17224 11577 17258 11611
rect 19533 11577 19567 11611
rect 21465 11577 21499 11611
rect 4077 11509 4111 11543
rect 5273 11509 5307 11543
rect 5917 11509 5951 11543
rect 8309 11509 8343 11543
rect 8677 11509 8711 11543
rect 9137 11509 9171 11543
rect 9597 11509 9631 11543
rect 10793 11509 10827 11543
rect 11161 11509 11195 11543
rect 12909 11509 12943 11543
rect 13553 11509 13587 11543
rect 13737 11509 13771 11543
rect 16313 11509 16347 11543
rect 16405 11509 16439 11543
rect 16773 11509 16807 11543
rect 1593 11305 1627 11339
rect 1777 11305 1811 11339
rect 3893 11305 3927 11339
rect 6101 11305 6135 11339
rect 8125 11305 8159 11339
rect 8585 11305 8619 11339
rect 9137 11305 9171 11339
rect 10609 11305 10643 11339
rect 14749 11305 14783 11339
rect 15117 11305 15151 11339
rect 15577 11305 15611 11339
rect 17601 11305 17635 11339
rect 17785 11305 17819 11339
rect 18613 11305 18647 11339
rect 19073 11305 19107 11339
rect 19625 11305 19659 11339
rect 21005 11305 21039 11339
rect 22017 11305 22051 11339
rect 3617 11237 3651 11271
rect 5273 11237 5307 11271
rect 5365 11237 5399 11271
rect 6193 11237 6227 11271
rect 6898 11237 6932 11271
rect 8953 11237 8987 11271
rect 10057 11237 10091 11271
rect 10149 11237 10183 11271
rect 11437 11237 11471 11271
rect 13185 11237 13219 11271
rect 13737 11237 13771 11271
rect 21281 11237 21315 11271
rect 1501 11169 1535 11203
rect 2890 11169 2924 11203
rect 3341 11169 3375 11203
rect 4261 11169 4295 11203
rect 4721 11169 4755 11203
rect 8493 11169 8527 11203
rect 3157 11101 3191 11135
rect 4353 11101 4387 11135
rect 4445 11101 4479 11135
rect 5181 11101 5215 11135
rect 5917 11101 5951 11135
rect 6653 11101 6687 11135
rect 8677 11101 8711 11135
rect 4905 11033 4939 11067
rect 9321 11169 9355 11203
rect 10977 11169 11011 11203
rect 11069 11169 11103 11203
rect 13645 11169 13679 11203
rect 14657 11169 14691 11203
rect 16037 11169 16071 11203
rect 16293 11169 16327 11203
rect 18521 11169 18555 11203
rect 19993 11169 20027 11203
rect 20821 11169 20855 11203
rect 21465 11169 21499 11203
rect 9689 11101 9723 11135
rect 9965 11101 9999 11135
rect 11253 11101 11287 11135
rect 13553 11101 13587 11135
rect 14473 11101 14507 11135
rect 15669 11101 15703 11135
rect 15761 11101 15795 11135
rect 18061 11101 18095 11135
rect 18429 11101 18463 11135
rect 20085 11101 20119 11135
rect 20177 11101 20211 11135
rect 20729 11101 20763 11135
rect 21189 11101 21223 11135
rect 9413 11033 9447 11067
rect 10517 11033 10551 11067
rect 14105 11033 14139 11067
rect 17417 11033 17451 11067
rect 3433 10965 3467 10999
rect 5733 10965 5767 10999
rect 6561 10965 6595 10999
rect 8033 10965 8067 10999
rect 8953 10965 8987 10999
rect 15209 10965 15243 10999
rect 18981 10965 19015 10999
rect 19441 10965 19475 10999
rect 20545 10965 20579 10999
rect 2237 10761 2271 10795
rect 4629 10761 4663 10795
rect 5549 10761 5583 10795
rect 6469 10761 6503 10795
rect 7389 10761 7423 10795
rect 11345 10761 11379 10795
rect 11529 10761 11563 10795
rect 13829 10761 13863 10795
rect 15025 10761 15059 10795
rect 16037 10761 16071 10795
rect 18521 10761 18555 10795
rect 19349 10761 19383 10795
rect 20453 10761 20487 10795
rect 20729 10761 20763 10795
rect 4721 10693 4755 10727
rect 7573 10693 7607 10727
rect 9229 10693 9263 10727
rect 11713 10693 11747 10727
rect 15945 10693 15979 10727
rect 20913 10693 20947 10727
rect 1685 10625 1719 10659
rect 2329 10625 2363 10659
rect 3985 10625 4019 10659
rect 5273 10625 5307 10659
rect 6101 10625 6135 10659
rect 6929 10625 6963 10659
rect 7021 10625 7055 10659
rect 8401 10625 8435 10659
rect 9137 10625 9171 10659
rect 13553 10625 13587 10659
rect 14657 10625 14691 10659
rect 15393 10625 15427 10659
rect 16681 10625 16715 10659
rect 17601 10625 17635 10659
rect 17969 10625 18003 10659
rect 18705 10625 18739 10659
rect 19625 10625 19659 10659
rect 5089 10557 5123 10591
rect 6837 10557 6871 10591
rect 8309 10557 8343 10591
rect 8769 10557 8803 10591
rect 9965 10557 9999 10591
rect 13286 10557 13320 10591
rect 13653 10557 13687 10591
rect 15577 10557 15611 10591
rect 16405 10557 16439 10591
rect 17325 10557 17359 10591
rect 18153 10557 18187 10591
rect 18981 10557 19015 10591
rect 20269 10557 20303 10591
rect 20545 10557 20579 10591
rect 2596 10489 2630 10523
rect 5181 10489 5215 10523
rect 8217 10489 8251 10523
rect 8953 10489 8987 10523
rect 10232 10489 10266 10523
rect 11989 10489 12023 10523
rect 14473 10489 14507 10523
rect 15485 10489 15519 10523
rect 18061 10489 18095 10523
rect 21097 10489 21131 10523
rect 21281 10489 21315 10523
rect 21465 10489 21499 10523
rect 1777 10421 1811 10455
rect 1869 10421 1903 10455
rect 3709 10421 3743 10455
rect 4169 10421 4203 10455
rect 4261 10421 4295 10455
rect 5917 10421 5951 10455
rect 6009 10421 6043 10455
rect 7665 10421 7699 10455
rect 7849 10421 7883 10455
rect 9413 10421 9447 10455
rect 9873 10421 9907 10455
rect 12173 10421 12207 10455
rect 13921 10421 13955 10455
rect 14105 10421 14139 10455
rect 14565 10421 14599 10455
rect 16497 10421 16531 10455
rect 16957 10421 16991 10455
rect 17417 10421 17451 10455
rect 18889 10421 18923 10455
rect 19717 10421 19751 10455
rect 19809 10421 19843 10455
rect 20177 10421 20211 10455
rect 1869 10217 1903 10251
rect 2329 10217 2363 10251
rect 3157 10217 3191 10251
rect 3617 10217 3651 10251
rect 3985 10217 4019 10251
rect 4445 10217 4479 10251
rect 5549 10217 5583 10251
rect 6561 10217 6595 10251
rect 7021 10217 7055 10251
rect 7573 10217 7607 10251
rect 7941 10217 7975 10251
rect 8401 10217 8435 10251
rect 10977 10217 11011 10251
rect 11529 10217 11563 10251
rect 11897 10217 11931 10251
rect 14473 10217 14507 10251
rect 15301 10217 15335 10251
rect 15669 10217 15703 10251
rect 16129 10217 16163 10251
rect 17233 10217 17267 10251
rect 17417 10217 17451 10251
rect 18981 10217 19015 10251
rect 19165 10217 19199 10251
rect 21005 10217 21039 10251
rect 4905 10149 4939 10183
rect 5273 10149 5307 10183
rect 6377 10149 6411 10183
rect 8033 10149 8067 10183
rect 10885 10149 10919 10183
rect 14013 10149 14047 10183
rect 16589 10149 16623 10183
rect 18552 10149 18586 10183
rect 2697 10081 2731 10115
rect 3341 10081 3375 10115
rect 4813 10081 4847 10115
rect 5917 10081 5951 10115
rect 7113 10081 7147 10115
rect 10250 10081 10284 10115
rect 11989 10081 12023 10115
rect 13562 10081 13596 10115
rect 13829 10081 13863 10115
rect 14105 10081 14139 10115
rect 14841 10081 14875 10115
rect 15761 10081 15795 10115
rect 16497 10081 16531 10115
rect 19892 10081 19926 10115
rect 21189 10081 21223 10115
rect 21557 10081 21591 10115
rect 1685 10013 1719 10047
rect 1777 10013 1811 10047
rect 2789 10013 2823 10047
rect 2881 10013 2915 10047
rect 5089 10013 5123 10047
rect 6009 10013 6043 10047
rect 6101 10013 6135 10047
rect 6929 10013 6963 10047
rect 8125 10013 8159 10047
rect 10517 10013 10551 10047
rect 10701 10013 10735 10047
rect 11805 10013 11839 10047
rect 14933 10013 14967 10047
rect 15025 10013 15059 10047
rect 15853 10013 15887 10047
rect 16773 10013 16807 10047
rect 18797 10013 18831 10047
rect 19625 10013 19659 10047
rect 2237 9945 2271 9979
rect 4353 9945 4387 9979
rect 8769 9945 8803 9979
rect 12357 9945 12391 9979
rect 21373 9945 21407 9979
rect 3433 9877 3467 9911
rect 4169 9877 4203 9911
rect 7481 9877 7515 9911
rect 8585 9877 8619 9911
rect 9137 9877 9171 9911
rect 11345 9877 11379 9911
rect 12449 9877 12483 9911
rect 16957 9877 16991 9911
rect 19441 9877 19475 9911
rect 1593 9673 1627 9707
rect 4721 9673 4755 9707
rect 10517 9673 10551 9707
rect 20545 9673 20579 9707
rect 6285 9605 6319 9639
rect 6469 9605 6503 9639
rect 8953 9605 8987 9639
rect 11437 9605 11471 9639
rect 15301 9605 15335 9639
rect 16405 9605 16439 9639
rect 16957 9605 16991 9639
rect 20453 9605 20487 9639
rect 2145 9537 2179 9571
rect 2973 9537 3007 9571
rect 4169 9537 4203 9571
rect 4261 9537 4295 9571
rect 8493 9537 8527 9571
rect 9137 9537 9171 9571
rect 10701 9537 10735 9571
rect 13093 9537 13127 9571
rect 14105 9537 14139 9571
rect 14933 9537 14967 9571
rect 15853 9537 15887 9571
rect 15945 9537 15979 9571
rect 17601 9537 17635 9571
rect 18429 9537 18463 9571
rect 21189 9537 21223 9571
rect 2789 9469 2823 9503
rect 3249 9469 3283 9503
rect 3801 9469 3835 9503
rect 4353 9469 4387 9503
rect 5937 9469 5971 9503
rect 6193 9469 6227 9503
rect 6285 9469 6319 9503
rect 6653 9469 6687 9503
rect 8769 9469 8803 9503
rect 10977 9469 11011 9503
rect 14749 9469 14783 9503
rect 15577 9469 15611 9503
rect 16037 9469 16071 9503
rect 16497 9469 16531 9503
rect 16773 9469 16807 9503
rect 17417 9469 17451 9503
rect 18153 9469 18187 9503
rect 19073 9469 19107 9503
rect 19340 9469 19374 9503
rect 21557 9469 21591 9503
rect 1961 9401 1995 9435
rect 8237 9401 8271 9435
rect 9382 9401 9416 9435
rect 12848 9401 12882 9435
rect 13921 9401 13955 9435
rect 14013 9401 14047 9435
rect 14841 9401 14875 9435
rect 17969 9401 18003 9435
rect 18613 9401 18647 9435
rect 1501 9333 1535 9367
rect 2053 9333 2087 9367
rect 2421 9333 2455 9367
rect 2881 9333 2915 9367
rect 3433 9333 3467 9367
rect 3617 9333 3651 9367
rect 4813 9333 4847 9367
rect 6745 9333 6779 9367
rect 7021 9333 7055 9367
rect 7113 9333 7147 9367
rect 8585 9333 8619 9367
rect 10885 9333 10919 9367
rect 11345 9333 11379 9367
rect 11713 9333 11747 9367
rect 13185 9333 13219 9367
rect 13369 9333 13403 9367
rect 13553 9333 13587 9367
rect 14381 9333 14415 9367
rect 17325 9333 17359 9367
rect 18521 9333 18555 9367
rect 18981 9333 19015 9367
rect 20913 9333 20947 9367
rect 21005 9333 21039 9367
rect 21373 9333 21407 9367
rect 2329 9129 2363 9163
rect 2789 9129 2823 9163
rect 3525 9129 3559 9163
rect 5457 9129 5491 9163
rect 7941 9129 7975 9163
rect 8309 9129 8343 9163
rect 10241 9129 10275 9163
rect 10701 9129 10735 9163
rect 11161 9129 11195 9163
rect 12725 9129 12759 9163
rect 12909 9129 12943 9163
rect 13093 9129 13127 9163
rect 13277 9129 13311 9163
rect 13737 9129 13771 9163
rect 14841 9129 14875 9163
rect 17509 9129 17543 9163
rect 17877 9129 17911 9163
rect 18705 9129 18739 9163
rect 21005 9129 21039 9163
rect 1869 9061 1903 9095
rect 7757 9061 7791 9095
rect 8401 9061 8435 9095
rect 9597 9061 9631 9095
rect 11621 9061 11655 9095
rect 12081 9061 12115 9095
rect 18613 9061 18647 9095
rect 1777 8993 1811 9027
rect 2697 8993 2731 9027
rect 3157 8993 3191 9027
rect 3893 8993 3927 9027
rect 4160 8993 4194 9027
rect 5917 8993 5951 9027
rect 6184 8993 6218 9027
rect 7481 8993 7515 9027
rect 9505 8993 9539 9027
rect 10333 8993 10367 9027
rect 12173 8993 12207 9027
rect 13645 8993 13679 9027
rect 14381 8993 14415 9027
rect 15393 8993 15427 9027
rect 16782 8993 16816 9027
rect 17049 8993 17083 9027
rect 18061 8993 18095 9027
rect 1685 8925 1719 8959
rect 2881 8925 2915 8959
rect 5825 8925 5859 8959
rect 8493 8925 8527 8959
rect 9781 8925 9815 8959
rect 10057 8925 10091 8959
rect 10885 8925 10919 8959
rect 11069 8925 11103 8959
rect 13829 8925 13863 8959
rect 15117 8925 15151 8959
rect 17233 8925 17267 8959
rect 17417 8925 17451 8959
rect 2237 8857 2271 8891
rect 3341 8857 3375 8891
rect 5273 8857 5307 8891
rect 7297 8857 7331 8891
rect 8861 8857 8895 8891
rect 11529 8857 11563 8891
rect 12449 8857 12483 8891
rect 12633 8857 12667 8891
rect 14197 8857 14231 8891
rect 15577 8857 15611 8891
rect 18245 8857 18279 8891
rect 19073 8993 19107 9027
rect 19165 8993 19199 9027
rect 19892 8993 19926 9027
rect 21189 8993 21223 9027
rect 21557 8993 21591 9027
rect 19349 8925 19383 8959
rect 19625 8925 19659 8959
rect 7665 8789 7699 8823
rect 9137 8789 9171 8823
rect 11805 8789 11839 8823
rect 14565 8789 14599 8823
rect 14749 8789 14783 8823
rect 15209 8789 15243 8823
rect 15669 8789 15703 8823
rect 18429 8789 18463 8823
rect 18613 8789 18647 8823
rect 21373 8789 21407 8823
rect 4353 8585 4387 8619
rect 4721 8585 4755 8619
rect 6469 8585 6503 8619
rect 8861 8585 8895 8619
rect 10701 8585 10735 8619
rect 11529 8585 11563 8619
rect 17785 8585 17819 8619
rect 20453 8585 20487 8619
rect 1685 8517 1719 8551
rect 1961 8517 1995 8551
rect 4445 8517 4479 8551
rect 6285 8517 6319 8551
rect 9781 8517 9815 8551
rect 11713 8517 11747 8551
rect 13001 8517 13035 8551
rect 16773 8517 16807 8551
rect 21373 8517 21407 8551
rect 2697 8449 2731 8483
rect 5365 8449 5399 8483
rect 5733 8449 5767 8483
rect 7113 8449 7147 8483
rect 7757 8449 7791 8483
rect 7849 8449 7883 8483
rect 8309 8449 8343 8483
rect 9505 8449 9539 8483
rect 10425 8449 10459 8483
rect 10977 8449 11011 8483
rect 11069 8449 11103 8483
rect 12265 8449 12299 8483
rect 13553 8449 13587 8483
rect 17049 8449 17083 8483
rect 18337 8449 18371 8483
rect 18797 8449 18831 8483
rect 19901 8449 19935 8483
rect 21097 8449 21131 8483
rect 1777 8381 1811 8415
rect 2513 8381 2547 8415
rect 2973 8381 3007 8415
rect 5089 8381 5123 8415
rect 5917 8381 5951 8415
rect 6837 8381 6871 8415
rect 6929 8381 6963 8415
rect 8493 8381 8527 8415
rect 9321 8381 9355 8415
rect 10241 8381 10275 8415
rect 12173 8381 12207 8415
rect 12725 8381 12759 8415
rect 15045 8381 15079 8415
rect 15301 8381 15335 8415
rect 15393 8381 15427 8415
rect 18889 8381 18923 8415
rect 19533 8381 19567 8415
rect 20913 8381 20947 8415
rect 21005 8381 21039 8415
rect 21557 8381 21591 8415
rect 1501 8313 1535 8347
rect 2605 8313 2639 8347
rect 3218 8313 3252 8347
rect 5181 8313 5215 8347
rect 7665 8313 7699 8347
rect 11161 8313 11195 8347
rect 12633 8313 12667 8347
rect 15660 8313 15694 8347
rect 17325 8313 17359 8347
rect 18245 8313 18279 8347
rect 18981 8313 19015 8347
rect 2145 8245 2179 8279
rect 5825 8245 5859 8279
rect 7297 8245 7331 8279
rect 8401 8245 8435 8279
rect 8953 8245 8987 8279
rect 9413 8245 9447 8279
rect 10149 8245 10183 8279
rect 12081 8245 12115 8279
rect 13369 8245 13403 8279
rect 13461 8245 13495 8279
rect 13921 8245 13955 8279
rect 17233 8245 17267 8279
rect 17693 8245 17727 8279
rect 18153 8245 18187 8279
rect 19349 8245 19383 8279
rect 19993 8245 20027 8279
rect 20085 8245 20119 8279
rect 20545 8245 20579 8279
rect 1593 8041 1627 8075
rect 3065 8041 3099 8075
rect 3341 8041 3375 8075
rect 4721 8041 4755 8075
rect 7113 8041 7147 8075
rect 7481 8041 7515 8075
rect 7573 8041 7607 8075
rect 8125 8041 8159 8075
rect 8217 8041 8251 8075
rect 8677 8041 8711 8075
rect 10977 8041 11011 8075
rect 12817 8041 12851 8075
rect 13461 8041 13495 8075
rect 14381 8041 14415 8075
rect 14841 8041 14875 8075
rect 15945 8041 15979 8075
rect 16589 8041 16623 8075
rect 17141 8041 17175 8075
rect 17509 8041 17543 8075
rect 20545 8041 20579 8075
rect 21557 8041 21591 8075
rect 6754 7973 6788 8007
rect 9404 7973 9438 8007
rect 10885 7973 10919 8007
rect 13921 7973 13955 8007
rect 15485 7973 15519 8007
rect 20913 7973 20947 8007
rect 1409 7905 1443 7939
rect 1952 7905 1986 7939
rect 3249 7905 3283 7939
rect 3525 7905 3559 7939
rect 4261 7905 4295 7939
rect 5089 7905 5123 7939
rect 7941 7905 7975 7939
rect 8585 7905 8619 7939
rect 9137 7905 9171 7939
rect 12101 7905 12135 7939
rect 12357 7905 12391 7939
rect 13369 7905 13403 7939
rect 13829 7905 13863 7939
rect 14749 7905 14783 7939
rect 15577 7905 15611 7939
rect 16497 7905 16531 7939
rect 18236 7905 18270 7939
rect 20085 7905 20119 7939
rect 1685 7837 1719 7871
rect 4353 7837 4387 7871
rect 4445 7837 4479 7871
rect 5181 7837 5215 7871
rect 5273 7837 5307 7871
rect 7021 7837 7055 7871
rect 7665 7837 7699 7871
rect 8861 7837 8895 7871
rect 12909 7837 12943 7871
rect 13001 7837 13035 7871
rect 14013 7837 14047 7871
rect 14933 7837 14967 7871
rect 15393 7837 15427 7871
rect 16037 7837 16071 7871
rect 16405 7837 16439 7871
rect 17601 7837 17635 7871
rect 17693 7837 17727 7871
rect 17969 7837 18003 7871
rect 19901 7837 19935 7871
rect 19993 7837 20027 7871
rect 21005 7837 21039 7871
rect 21097 7837 21131 7871
rect 3893 7769 3927 7803
rect 12449 7769 12483 7803
rect 16957 7769 16991 7803
rect 3709 7701 3743 7735
rect 5641 7701 5675 7735
rect 10517 7701 10551 7735
rect 10609 7701 10643 7735
rect 19349 7701 19383 7735
rect 20453 7701 20487 7735
rect 1869 7497 1903 7531
rect 3341 7497 3375 7531
rect 4169 7497 4203 7531
rect 4997 7497 5031 7531
rect 6469 7497 6503 7531
rect 9137 7497 9171 7531
rect 10885 7497 10919 7531
rect 17969 7497 18003 7531
rect 19349 7497 19383 7531
rect 19625 7497 19659 7531
rect 6193 7429 6227 7463
rect 9045 7429 9079 7463
rect 10057 7429 10091 7463
rect 13277 7429 13311 7463
rect 15301 7429 15335 7463
rect 18797 7429 18831 7463
rect 3985 7361 4019 7395
rect 4813 7361 4847 7395
rect 5549 7361 5583 7395
rect 6929 7361 6963 7395
rect 7021 7361 7055 7395
rect 7665 7361 7699 7395
rect 9597 7361 9631 7395
rect 9689 7361 9723 7395
rect 14013 7361 14047 7395
rect 14749 7361 14783 7395
rect 16037 7361 16071 7395
rect 17141 7361 17175 7395
rect 17417 7361 17451 7395
rect 18245 7361 18279 7395
rect 20269 7361 20303 7395
rect 21005 7361 21039 7395
rect 1501 7293 1535 7327
rect 3249 7293 3283 7327
rect 4629 7293 4663 7327
rect 9505 7293 9539 7327
rect 11713 7293 11747 7327
rect 13737 7293 13771 7327
rect 14657 7293 14691 7327
rect 16681 7293 16715 7327
rect 17509 7293 17543 7327
rect 17601 7293 17635 7327
rect 19165 7293 19199 7327
rect 19441 7293 19475 7327
rect 20821 7293 20855 7327
rect 21557 7293 21591 7327
rect 1685 7225 1719 7259
rect 2993 7225 3027 7259
rect 3801 7225 3835 7259
rect 5825 7225 5859 7259
rect 7910 7225 7944 7259
rect 10149 7225 10183 7259
rect 11958 7225 11992 7259
rect 13829 7225 13863 7259
rect 14565 7225 14599 7259
rect 15025 7225 15059 7259
rect 16221 7225 16255 7259
rect 20085 7225 20119 7259
rect 3709 7157 3743 7191
rect 4537 7157 4571 7191
rect 5365 7157 5399 7191
rect 5457 7157 5491 7191
rect 6009 7157 6043 7191
rect 6837 7157 6871 7191
rect 7297 7157 7331 7191
rect 7481 7157 7515 7191
rect 10333 7157 10367 7191
rect 10609 7157 10643 7191
rect 11069 7157 11103 7191
rect 11161 7157 11195 7191
rect 11437 7157 11471 7191
rect 13093 7157 13127 7191
rect 13369 7157 13403 7191
rect 14197 7157 14231 7191
rect 15485 7157 15519 7191
rect 15669 7157 15703 7191
rect 16129 7157 16163 7191
rect 16589 7157 16623 7191
rect 18337 7157 18371 7191
rect 18429 7157 18463 7191
rect 18889 7157 18923 7191
rect 19993 7157 20027 7191
rect 20453 7157 20487 7191
rect 20913 7157 20947 7191
rect 21373 7157 21407 7191
rect 2329 6953 2363 6987
rect 2697 6953 2731 6987
rect 3157 6953 3191 6987
rect 6101 6953 6135 6987
rect 6469 6953 6503 6987
rect 6929 6953 6963 6987
rect 7297 6953 7331 6987
rect 10333 6953 10367 6987
rect 11253 6953 11287 6987
rect 13737 6953 13771 6987
rect 14105 6953 14139 6987
rect 15853 6953 15887 6987
rect 16497 6953 16531 6987
rect 16957 6953 16991 6987
rect 18797 6953 18831 6987
rect 20177 6953 20211 6987
rect 21005 6953 21039 6987
rect 21557 6953 21591 6987
rect 1685 6885 1719 6919
rect 3617 6885 3651 6919
rect 7389 6885 7423 6919
rect 9689 6885 9723 6919
rect 11345 6885 11379 6919
rect 15025 6885 15059 6919
rect 15485 6885 15519 6919
rect 15945 6885 15979 6919
rect 17417 6885 17451 6919
rect 1501 6817 1535 6851
rect 5006 6817 5040 6851
rect 5273 6817 5307 6851
rect 5557 6817 5591 6851
rect 5825 6817 5859 6851
rect 8677 6817 8711 6851
rect 9229 6817 9263 6851
rect 2145 6749 2179 6783
rect 2237 6749 2271 6783
rect 3249 6749 3283 6783
rect 3341 6749 3375 6783
rect 5917 6749 5951 6783
rect 6561 6749 6595 6783
rect 6653 6749 6687 6783
rect 7481 6749 7515 6783
rect 8309 6749 8343 6783
rect 9505 6749 9539 6783
rect 2789 6681 2823 6715
rect 5365 6681 5399 6715
rect 8125 6681 8159 6715
rect 8493 6681 8527 6715
rect 10885 6817 10919 6851
rect 12918 6817 12952 6851
rect 13645 6817 13679 6851
rect 14565 6817 14599 6851
rect 17325 6817 17359 6851
rect 18337 6817 18371 6851
rect 18429 6817 18463 6851
rect 19073 6817 19107 6851
rect 19349 6817 19383 6851
rect 20085 6817 20119 6851
rect 21097 6817 21131 6851
rect 9781 6749 9815 6783
rect 10425 6749 10459 6783
rect 10517 6749 10551 6783
rect 11161 6749 11195 6783
rect 13185 6749 13219 6783
rect 13829 6749 13863 6783
rect 15301 6749 15335 6783
rect 15393 6749 15427 6783
rect 16589 6749 16623 6783
rect 16681 6749 16715 6783
rect 17509 6749 17543 6783
rect 17785 6749 17819 6783
rect 18153 6749 18187 6783
rect 19165 6749 19199 6783
rect 19901 6749 19935 6783
rect 21189 6749 21223 6783
rect 19717 6681 19751 6715
rect 20545 6681 20579 6715
rect 1777 6613 1811 6647
rect 3893 6613 3927 6647
rect 5641 6613 5675 6647
rect 7757 6613 7791 6647
rect 7941 6613 7975 6647
rect 8861 6613 8895 6647
rect 9413 6613 9447 6647
rect 9689 6613 9723 6647
rect 9965 6613 9999 6647
rect 11713 6613 11747 6647
rect 11805 6613 11839 6647
rect 13277 6613 13311 6647
rect 14381 6613 14415 6647
rect 14657 6613 14691 6647
rect 16129 6613 16163 6647
rect 20637 6613 20671 6647
rect 1961 6409 1995 6443
rect 2789 6409 2823 6443
rect 4629 6409 4663 6443
rect 5457 6409 5491 6443
rect 8033 6409 8067 6443
rect 10333 6409 10367 6443
rect 12265 6409 12299 6443
rect 13093 6409 13127 6443
rect 21373 6409 21407 6443
rect 22017 6409 22051 6443
rect 1593 6341 1627 6375
rect 4353 6341 4387 6375
rect 13921 6341 13955 6375
rect 15025 6341 15059 6375
rect 18521 6341 18555 6375
rect 20637 6341 20671 6375
rect 2237 6273 2271 6307
rect 3985 6273 4019 6307
rect 5089 6273 5123 6307
rect 5181 6273 5215 6307
rect 6009 6273 6043 6307
rect 6929 6273 6963 6307
rect 7113 6273 7147 6307
rect 7389 6273 7423 6307
rect 7573 6273 7607 6307
rect 8953 6273 8987 6307
rect 9781 6273 9815 6307
rect 10517 6273 10551 6307
rect 12725 6273 12759 6307
rect 12817 6273 12851 6307
rect 13553 6273 13587 6307
rect 13645 6273 13679 6307
rect 14289 6273 14323 6307
rect 14473 6273 14507 6307
rect 15853 6273 15887 6307
rect 16773 6273 16807 6307
rect 17509 6273 17543 6307
rect 17877 6273 17911 6307
rect 19257 6273 19291 6307
rect 1409 6205 1443 6239
rect 1777 6205 1811 6239
rect 4169 6205 4203 6239
rect 7665 6205 7699 6239
rect 9965 6205 9999 6239
rect 10701 6205 10735 6239
rect 13461 6205 13495 6239
rect 14565 6205 14599 6239
rect 15485 6205 15519 6239
rect 16037 6205 16071 6239
rect 2421 6137 2455 6171
rect 2881 6137 2915 6171
rect 4445 6137 4479 6171
rect 4997 6137 5031 6171
rect 8125 6137 8159 6171
rect 8861 6137 8895 6171
rect 9321 6137 9355 6171
rect 11345 6137 11379 6171
rect 12633 6137 12667 6171
rect 15945 6137 15979 6171
rect 19165 6137 19199 6171
rect 19524 6137 19558 6171
rect 20913 6137 20947 6171
rect 21097 6137 21131 6171
rect 21465 6137 21499 6171
rect 2329 6069 2363 6103
rect 3157 6069 3191 6103
rect 3341 6069 3375 6103
rect 3709 6069 3743 6103
rect 3801 6069 3835 6103
rect 5825 6069 5859 6103
rect 5917 6069 5951 6103
rect 6469 6069 6503 6103
rect 6837 6069 6871 6103
rect 8401 6069 8435 6103
rect 8769 6069 8803 6103
rect 9413 6069 9447 6103
rect 9873 6069 9907 6103
rect 10793 6069 10827 6103
rect 11161 6069 11195 6103
rect 11437 6069 11471 6103
rect 11713 6069 11747 6103
rect 11897 6069 11931 6103
rect 12173 6069 12207 6103
rect 14933 6069 14967 6103
rect 15301 6069 15335 6103
rect 16405 6069 16439 6103
rect 16957 6069 16991 6103
rect 17325 6069 17359 6103
rect 17417 6069 17451 6103
rect 18061 6069 18095 6103
rect 18153 6069 18187 6103
rect 18797 6069 18831 6103
rect 18981 6069 19015 6103
rect 1593 5865 1627 5899
rect 3157 5865 3191 5899
rect 3893 5865 3927 5899
rect 5549 5865 5583 5899
rect 6377 5865 6411 5899
rect 6745 5865 6779 5899
rect 6837 5865 6871 5899
rect 11713 5865 11747 5899
rect 12173 5865 12207 5899
rect 16221 5865 16255 5899
rect 16589 5865 16623 5899
rect 17417 5865 17451 5899
rect 18061 5865 18095 5899
rect 20177 5865 20211 5899
rect 20637 5865 20671 5899
rect 2022 5797 2056 5831
rect 7481 5797 7515 5831
rect 8125 5797 8159 5831
rect 8585 5797 8619 5831
rect 11253 5797 11287 5831
rect 12786 5797 12820 5831
rect 14105 5797 14139 5831
rect 14626 5797 14660 5831
rect 20913 5797 20947 5831
rect 21097 5797 21131 5831
rect 22017 5797 22051 5831
rect 1409 5729 1443 5763
rect 3341 5729 3375 5763
rect 4169 5729 4203 5763
rect 4436 5729 4470 5763
rect 5825 5729 5859 5763
rect 6101 5729 6135 5763
rect 7389 5729 7423 5763
rect 10526 5729 10560 5763
rect 12081 5729 12115 5763
rect 12541 5729 12575 5763
rect 16957 5729 16991 5763
rect 17049 5729 17083 5763
rect 19174 5729 19208 5763
rect 20453 5729 20487 5763
rect 21465 5729 21499 5763
rect 1777 5661 1811 5695
rect 3617 5661 3651 5695
rect 6929 5661 6963 5695
rect 8217 5661 8251 5695
rect 8401 5661 8435 5695
rect 10793 5661 10827 5695
rect 11345 5661 11379 5695
rect 11437 5661 11471 5695
rect 12265 5661 12299 5695
rect 14381 5661 14415 5695
rect 15945 5661 15979 5695
rect 16129 5661 16163 5695
rect 16773 5661 16807 5695
rect 19441 5661 19475 5695
rect 19901 5661 19935 5695
rect 21281 5661 21315 5695
rect 7205 5593 7239 5627
rect 8861 5593 8895 5627
rect 9413 5593 9447 5627
rect 10885 5593 10919 5627
rect 15761 5593 15795 5627
rect 17693 5593 17727 5627
rect 17969 5593 18003 5627
rect 19717 5593 19751 5627
rect 3525 5525 3559 5559
rect 5641 5525 5675 5559
rect 5917 5525 5951 5559
rect 6193 5525 6227 5559
rect 7757 5525 7791 5559
rect 9137 5525 9171 5559
rect 13921 5525 13955 5559
rect 20085 5525 20119 5559
rect 20821 5525 20855 5559
rect 1869 5321 1903 5355
rect 4077 5321 4111 5355
rect 6745 5321 6779 5355
rect 8861 5321 8895 5355
rect 14933 5321 14967 5355
rect 16405 5321 16439 5355
rect 17693 5321 17727 5355
rect 17969 5321 18003 5355
rect 19441 5321 19475 5355
rect 20269 5321 20303 5355
rect 20729 5321 20763 5355
rect 1593 5253 1627 5287
rect 2421 5185 2455 5219
rect 2697 5185 2731 5219
rect 4629 5185 4663 5219
rect 4813 5185 4847 5219
rect 6009 5185 6043 5219
rect 9045 5253 9079 5287
rect 20637 5253 20671 5287
rect 7021 5185 7055 5219
rect 8217 5185 8251 5219
rect 10793 5185 10827 5219
rect 10977 5185 11011 5219
rect 12173 5185 12207 5219
rect 12357 5185 12391 5219
rect 12725 5185 12759 5219
rect 12817 5185 12851 5219
rect 13921 5185 13955 5219
rect 14289 5185 14323 5219
rect 15025 5185 15059 5219
rect 17049 5185 17083 5219
rect 18061 5185 18095 5219
rect 19625 5185 19659 5219
rect 21281 5185 21315 5219
rect 1409 5117 1443 5151
rect 4537 5117 4571 5151
rect 5181 5117 5215 5151
rect 5825 5117 5859 5151
rect 6469 5117 6503 5151
rect 6745 5117 6779 5151
rect 8033 5117 8067 5151
rect 8585 5117 8619 5151
rect 10342 5117 10376 5151
rect 10609 5117 10643 5151
rect 11069 5117 11103 5151
rect 12081 5117 12115 5151
rect 12909 5117 12943 5151
rect 14565 5117 14599 5151
rect 15292 5117 15326 5151
rect 17325 5117 17359 5151
rect 20453 5117 20487 5151
rect 20913 5117 20947 5151
rect 21189 5117 21223 5151
rect 2942 5049 2976 5083
rect 16681 5049 16715 5083
rect 17233 5049 17267 5083
rect 18306 5049 18340 5083
rect 19901 5049 19935 5083
rect 21465 5049 21499 5083
rect 2237 4981 2271 5015
rect 2329 4981 2363 5015
rect 4169 4981 4203 5015
rect 4997 4981 5031 5015
rect 5273 4981 5307 5015
rect 5457 4981 5491 5015
rect 5917 4981 5951 5015
rect 6653 4981 6687 5015
rect 7113 4981 7147 5015
rect 7205 4981 7239 5015
rect 7573 4981 7607 5015
rect 7665 4981 7699 5015
rect 8125 4981 8159 5015
rect 8677 4981 8711 5015
rect 9229 4981 9263 5015
rect 11437 4981 11471 5015
rect 11713 4981 11747 5015
rect 13277 4981 13311 5015
rect 13369 4981 13403 5015
rect 13737 4981 13771 5015
rect 13829 4981 13863 5015
rect 14473 4981 14507 5015
rect 16589 4981 16623 5015
rect 19809 4981 19843 5015
rect 21005 4981 21039 5015
rect 1409 4777 1443 4811
rect 2973 4777 3007 4811
rect 3341 4777 3375 4811
rect 3893 4777 3927 4811
rect 4353 4777 4387 4811
rect 4721 4777 4755 4811
rect 5181 4777 5215 4811
rect 7297 4777 7331 4811
rect 7757 4777 7791 4811
rect 8585 4777 8619 4811
rect 10241 4777 10275 4811
rect 10701 4777 10735 4811
rect 11161 4777 11195 4811
rect 12265 4777 12299 4811
rect 14933 4777 14967 4811
rect 16957 4777 16991 4811
rect 17969 4777 18003 4811
rect 18797 4777 18831 4811
rect 19625 4777 19659 4811
rect 20085 4777 20119 4811
rect 20453 4777 20487 4811
rect 20729 4777 20763 4811
rect 21373 4777 21407 4811
rect 4261 4709 4295 4743
rect 6776 4709 6810 4743
rect 7849 4709 7883 4743
rect 10609 4709 10643 4743
rect 11989 4709 12023 4743
rect 14381 4709 14415 4743
rect 15844 4709 15878 4743
rect 17601 4709 17635 4743
rect 2533 4641 2567 4675
rect 5089 4641 5123 4675
rect 7113 4641 7147 4675
rect 9137 4641 9171 4675
rect 9873 4641 9907 4675
rect 11529 4641 11563 4675
rect 2789 4573 2823 4607
rect 3433 4573 3467 4607
rect 3525 4573 3559 4607
rect 4445 4573 4479 4607
rect 5273 4573 5307 4607
rect 7021 4573 7055 4607
rect 8033 4573 8067 4607
rect 8309 4573 8343 4607
rect 8493 4573 8527 4607
rect 9597 4573 9631 4607
rect 9781 4573 9815 4607
rect 10517 4573 10551 4607
rect 11621 4573 11655 4607
rect 11805 4573 11839 4607
rect 5641 4505 5675 4539
rect 12081 4641 12115 4675
rect 12541 4641 12575 4675
rect 13838 4641 13872 4675
rect 14105 4641 14139 4675
rect 15209 4641 15243 4675
rect 15577 4641 15611 4675
rect 18429 4641 18463 4675
rect 19165 4641 19199 4675
rect 19993 4641 20027 4675
rect 20637 4641 20671 4675
rect 20913 4641 20947 4675
rect 21189 4641 21223 4675
rect 21465 4641 21499 4675
rect 14657 4573 14691 4607
rect 17417 4573 17451 4607
rect 17509 4573 17543 4607
rect 18245 4573 18279 4607
rect 18337 4573 18371 4607
rect 20177 4573 20211 4607
rect 12725 4505 12759 4539
rect 7389 4437 7423 4471
rect 8953 4437 8987 4471
rect 9321 4437 9355 4471
rect 11069 4437 11103 4471
rect 11989 4437 12023 4471
rect 12357 4437 12391 4471
rect 14749 4437 14783 4471
rect 15393 4437 15427 4471
rect 17141 4437 17175 4471
rect 19073 4437 19107 4471
rect 19441 4437 19475 4471
rect 21005 4437 21039 4471
rect 2697 4233 2731 4267
rect 6285 4233 6319 4267
rect 8217 4233 8251 4267
rect 15761 4233 15795 4267
rect 17693 4233 17727 4267
rect 19165 4233 19199 4267
rect 8309 4165 8343 4199
rect 9505 4165 9539 4199
rect 20453 4165 20487 4199
rect 20821 4165 20855 4199
rect 1961 4097 1995 4131
rect 4077 4097 4111 4131
rect 5273 4097 5307 4131
rect 5733 4097 5767 4131
rect 6837 4097 6871 4131
rect 8769 4097 8803 4131
rect 8861 4097 8895 4131
rect 9137 4097 9171 4131
rect 10057 4097 10091 4131
rect 11069 4097 11103 4131
rect 12173 4097 12207 4131
rect 12265 4097 12299 4131
rect 13369 4097 13403 4131
rect 14105 4097 14139 4131
rect 15117 4097 15151 4131
rect 19073 4097 19107 4131
rect 19809 4097 19843 4131
rect 19993 4097 20027 4131
rect 1409 4029 1443 4063
rect 2145 4029 2179 4063
rect 4353 4029 4387 4063
rect 4629 4029 4663 4063
rect 6653 4029 6687 4063
rect 8677 4029 8711 4063
rect 10517 4029 10551 4063
rect 10793 4029 10827 4063
rect 11437 4029 11471 4063
rect 11713 4029 11747 4063
rect 13185 4029 13219 4063
rect 13645 4029 13679 4063
rect 14381 4029 14415 4063
rect 14657 4029 14691 4063
rect 15945 4029 15979 4063
rect 16313 4029 16347 4063
rect 16589 4029 16623 4063
rect 16957 4029 16991 4063
rect 17417 4029 17451 4063
rect 18806 4029 18840 4063
rect 20269 4029 20303 4063
rect 20729 4029 20763 4063
rect 21005 4029 21039 4063
rect 21281 4029 21315 4063
rect 21557 4029 21591 4063
rect 2237 3961 2271 3995
rect 3832 3961 3866 3995
rect 5917 3961 5951 3995
rect 7082 3961 7116 3995
rect 9321 3961 9355 3995
rect 9965 3961 9999 3995
rect 10885 3961 10919 3995
rect 11253 3961 11287 3995
rect 13921 3961 13955 3995
rect 15301 3961 15335 3995
rect 19625 3961 19659 3995
rect 22017 3961 22051 3995
rect 1593 3893 1627 3927
rect 1777 3893 1811 3927
rect 2605 3893 2639 3927
rect 4169 3893 4203 3927
rect 4445 3893 4479 3927
rect 4721 3893 4755 3927
rect 5089 3893 5123 3927
rect 5181 3893 5215 3927
rect 5825 3893 5859 3927
rect 6469 3893 6503 3927
rect 9873 3893 9907 3927
rect 10333 3893 10367 3927
rect 10609 3893 10643 3927
rect 11897 3893 11931 3927
rect 12357 3893 12391 3927
rect 12725 3893 12759 3927
rect 12817 3893 12851 3927
rect 13277 3893 13311 3927
rect 13829 3893 13863 3927
rect 14565 3893 14599 3927
rect 14841 3893 14875 3927
rect 15209 3893 15243 3927
rect 15669 3893 15703 3927
rect 16129 3893 16163 3927
rect 16497 3893 16531 3927
rect 16773 3893 16807 3927
rect 17141 3893 17175 3927
rect 17601 3893 17635 3927
rect 19533 3893 19567 3927
rect 20545 3893 20579 3927
rect 21097 3893 21131 3927
rect 21373 3893 21407 3927
rect 1593 3689 1627 3723
rect 2145 3689 2179 3723
rect 2973 3689 3007 3723
rect 4261 3689 4295 3723
rect 6285 3689 6319 3723
rect 8217 3689 8251 3723
rect 9321 3689 9355 3723
rect 12725 3689 12759 3723
rect 14933 3689 14967 3723
rect 15393 3689 15427 3723
rect 18705 3689 18739 3723
rect 20085 3689 20119 3723
rect 3341 3621 3375 3655
rect 5374 3621 5408 3655
rect 6193 3621 6227 3655
rect 9229 3621 9263 3655
rect 12817 3621 12851 3655
rect 13645 3621 13679 3655
rect 21373 3621 21407 3655
rect 1409 3553 1443 3587
rect 1685 3553 1719 3587
rect 2513 3553 2547 3587
rect 3433 3553 3467 3587
rect 5641 3553 5675 3587
rect 7858 3553 7892 3587
rect 8585 3553 8619 3587
rect 10629 3553 10663 3587
rect 12090 3553 12124 3587
rect 12357 3553 12391 3587
rect 13737 3553 13771 3587
rect 14381 3553 14415 3587
rect 15025 3553 15059 3587
rect 15485 3553 15519 3587
rect 15761 3553 15795 3587
rect 17242 3553 17276 3587
rect 17601 3553 17635 3587
rect 17877 3553 17911 3587
rect 19165 3553 19199 3587
rect 19993 3553 20027 3587
rect 20453 3553 20487 3587
rect 21005 3553 21039 3587
rect 2605 3485 2639 3519
rect 2697 3485 2731 3519
rect 3617 3485 3651 3519
rect 3893 3485 3927 3519
rect 6009 3485 6043 3519
rect 8125 3485 8159 3519
rect 8677 3485 8711 3519
rect 8769 3485 8803 3519
rect 10885 3485 10919 3519
rect 12633 3485 12667 3519
rect 13829 3485 13863 3519
rect 14841 3485 14875 3519
rect 17509 3485 17543 3519
rect 18429 3485 18463 3519
rect 18613 3485 18647 3519
rect 20177 3485 20211 3519
rect 20821 3485 20855 3519
rect 1869 3417 1903 3451
rect 6653 3417 6687 3451
rect 14105 3417 14139 3451
rect 16129 3417 16163 3451
rect 18061 3417 18095 3451
rect 19625 3417 19659 3451
rect 21557 3417 21591 3451
rect 1961 3349 1995 3383
rect 5733 3349 5767 3383
rect 6745 3349 6779 3383
rect 9505 3349 9539 3383
rect 10977 3349 11011 3383
rect 13185 3349 13219 3383
rect 13277 3349 13311 3383
rect 15669 3349 15703 3383
rect 15945 3349 15979 3383
rect 17785 3349 17819 3383
rect 18245 3349 18279 3383
rect 19073 3349 19107 3383
rect 19349 3349 19383 3383
rect 20637 3349 20671 3383
rect 21097 3349 21131 3383
rect 2053 3145 2087 3179
rect 3065 3145 3099 3179
rect 5273 3145 5307 3179
rect 6285 3145 6319 3179
rect 8493 3145 8527 3179
rect 10977 3145 11011 3179
rect 11713 3145 11747 3179
rect 18337 3145 18371 3179
rect 19165 3145 19199 3179
rect 1593 3077 1627 3111
rect 6469 3077 6503 3111
rect 6837 3077 6871 3111
rect 15577 3077 15611 3111
rect 19441 3077 19475 3111
rect 19717 3077 19751 3111
rect 3617 3009 3651 3043
rect 3893 3009 3927 3043
rect 5733 3009 5767 3043
rect 9045 3009 9079 3043
rect 13645 3009 13679 3043
rect 13737 3009 13771 3043
rect 16957 3009 16991 3043
rect 18521 3009 18555 3043
rect 1409 2941 1443 2975
rect 1869 2941 1903 2975
rect 2237 2941 2271 2975
rect 2697 2941 2731 2975
rect 3525 2941 3559 2975
rect 4160 2941 4194 2975
rect 5917 2941 5951 2975
rect 7961 2941 7995 2975
rect 8217 2941 8251 2975
rect 8861 2941 8895 2975
rect 10526 2941 10560 2975
rect 10793 2941 10827 2975
rect 11253 2941 11287 2975
rect 13093 2941 13127 2975
rect 13553 2941 13587 2975
rect 14197 2941 14231 2975
rect 14289 2941 14323 2975
rect 14565 2941 14599 2975
rect 14841 2941 14875 2975
rect 15117 2941 15151 2975
rect 15393 2941 15427 2975
rect 15853 2941 15887 2975
rect 16221 2941 16255 2975
rect 16681 2941 16715 2975
rect 19257 2941 19291 2975
rect 19533 2941 19567 2975
rect 19993 2941 20027 2975
rect 20821 2941 20855 2975
rect 21189 2941 21223 2975
rect 1685 2873 1719 2907
rect 6653 2873 6687 2907
rect 8953 2873 8987 2907
rect 11069 2873 11103 2907
rect 12848 2873 12882 2907
rect 15669 2873 15703 2907
rect 16037 2873 16071 2907
rect 17202 2873 17236 2907
rect 19809 2873 19843 2907
rect 20269 2873 20303 2907
rect 20453 2873 20487 2907
rect 20637 2873 20671 2907
rect 21373 2873 21407 2907
rect 2421 2805 2455 2839
rect 2513 2805 2547 2839
rect 2881 2805 2915 2839
rect 3433 2805 3467 2839
rect 5825 2805 5859 2839
rect 8309 2805 8343 2839
rect 9413 2805 9447 2839
rect 11437 2805 11471 2839
rect 13185 2805 13219 2839
rect 14013 2805 14047 2839
rect 14473 2805 14507 2839
rect 14749 2805 14783 2839
rect 15025 2805 15059 2839
rect 15301 2805 15335 2839
rect 16589 2805 16623 2839
rect 18705 2805 18739 2839
rect 18797 2805 18831 2839
rect 21005 2805 21039 2839
rect 21465 2805 21499 2839
rect 22017 2805 22051 2839
rect 2881 2601 2915 2635
rect 3341 2601 3375 2635
rect 4077 2601 4111 2635
rect 4445 2601 4479 2635
rect 5641 2601 5675 2635
rect 6745 2601 6779 2635
rect 7021 2601 7055 2635
rect 7297 2601 7331 2635
rect 7665 2601 7699 2635
rect 8585 2601 8619 2635
rect 10241 2601 10275 2635
rect 10517 2601 10551 2635
rect 11253 2601 11287 2635
rect 11897 2601 11931 2635
rect 12265 2601 12299 2635
rect 12357 2601 12391 2635
rect 12817 2601 12851 2635
rect 14381 2601 14415 2635
rect 17601 2601 17635 2635
rect 18061 2601 18095 2635
rect 18521 2601 18555 2635
rect 18613 2601 18647 2635
rect 19073 2601 19107 2635
rect 19993 2601 20027 2635
rect 21373 2601 21407 2635
rect 3249 2533 3283 2567
rect 4537 2533 4571 2567
rect 5181 2533 5215 2567
rect 7757 2533 7791 2567
rect 9597 2533 9631 2567
rect 10149 2533 10183 2567
rect 11345 2533 11379 2567
rect 14013 2533 14047 2567
rect 14749 2533 14783 2567
rect 15117 2533 15151 2567
rect 15485 2533 15519 2567
rect 16221 2533 16255 2567
rect 16589 2533 16623 2567
rect 16865 2533 16899 2567
rect 17417 2533 17451 2567
rect 18153 2533 18187 2567
rect 18981 2533 19015 2567
rect 20453 2533 20487 2567
rect 20821 2533 20855 2567
rect 21189 2533 21223 2567
rect 1409 2465 1443 2499
rect 1685 2465 1719 2499
rect 1961 2465 1995 2499
rect 2237 2465 2271 2499
rect 2605 2465 2639 2499
rect 3985 2465 4019 2499
rect 4905 2465 4939 2499
rect 5365 2465 5399 2499
rect 6009 2465 6043 2499
rect 6653 2465 6687 2499
rect 7205 2465 7239 2499
rect 8493 2465 8527 2499
rect 10609 2465 10643 2499
rect 12909 2465 12943 2499
rect 13093 2465 13127 2499
rect 13277 2465 13311 2499
rect 13645 2465 13679 2499
rect 14197 2465 14231 2499
rect 14565 2465 14599 2499
rect 15853 2465 15887 2499
rect 19625 2465 19659 2499
rect 20085 2465 20119 2499
rect 21557 2465 21591 2499
rect 3525 2397 3559 2431
rect 4721 2397 4755 2431
rect 6101 2397 6135 2431
rect 6193 2397 6227 2431
rect 7941 2397 7975 2431
rect 8769 2397 8803 2431
rect 9689 2397 9723 2431
rect 9781 2397 9815 2431
rect 11069 2397 11103 2431
rect 12449 2397 12483 2431
rect 14933 2397 14967 2431
rect 16405 2397 16439 2431
rect 17049 2397 17083 2431
rect 17969 2397 18003 2431
rect 19165 2397 19199 2431
rect 20637 2397 20671 2431
rect 2789 2329 2823 2363
rect 8125 2329 8159 2363
rect 9229 2329 9263 2363
rect 10793 2329 10827 2363
rect 11713 2329 11747 2363
rect 13829 2329 13863 2363
rect 16037 2329 16071 2363
rect 17233 2329 17267 2363
rect 19441 2329 19475 2363
rect 20269 2329 20303 2363
rect 1593 2261 1627 2295
rect 1869 2261 1903 2295
rect 2145 2261 2179 2295
rect 2421 2261 2455 2295
rect 5089 2261 5123 2295
rect 8953 2261 8987 2295
rect 13553 2261 13587 2295
rect 15393 2261 15427 2295
rect 15761 2261 15795 2295
rect 21097 2261 21131 2295
rect 6653 1853 6687 1887
rect 6837 1853 6871 1887
<< metal1 >>
rect 2866 21904 2872 21956
rect 2924 21944 2930 21956
rect 3142 21944 3148 21956
rect 2924 21916 3148 21944
rect 2924 21904 2930 21916
rect 3142 21904 3148 21916
rect 3200 21904 3206 21956
rect 7098 20748 7104 20800
rect 7156 20788 7162 20800
rect 8846 20788 8852 20800
rect 7156 20760 8852 20788
rect 7156 20748 7162 20760
rect 8846 20748 8852 20760
rect 8904 20748 8910 20800
rect 18046 20748 18052 20800
rect 18104 20788 18110 20800
rect 19334 20788 19340 20800
rect 18104 20760 19340 20788
rect 18104 20748 18110 20760
rect 19334 20748 19340 20760
rect 19392 20748 19398 20800
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 1854 20584 1860 20596
rect 1815 20556 1860 20584
rect 1854 20544 1860 20556
rect 1912 20544 1918 20596
rect 2222 20584 2228 20596
rect 2183 20556 2228 20584
rect 2222 20544 2228 20556
rect 2280 20544 2286 20596
rect 2593 20587 2651 20593
rect 2593 20553 2605 20587
rect 2639 20584 2651 20587
rect 2774 20584 2780 20596
rect 2639 20556 2780 20584
rect 2639 20553 2651 20556
rect 2593 20547 2651 20553
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 7285 20587 7343 20593
rect 3160 20556 6776 20584
rect 2866 20516 2872 20528
rect 2827 20488 2872 20516
rect 2866 20476 2872 20488
rect 2924 20476 2930 20528
rect 934 20408 940 20460
rect 992 20448 998 20460
rect 2682 20448 2688 20460
rect 992 20420 2688 20448
rect 992 20408 998 20420
rect 2682 20408 2688 20420
rect 2740 20408 2746 20460
rect 566 20340 572 20392
rect 624 20380 630 20392
rect 2406 20380 2412 20392
rect 624 20352 2412 20380
rect 624 20340 630 20352
rect 2406 20340 2412 20352
rect 2464 20340 2470 20392
rect 3053 20383 3111 20389
rect 3053 20349 3065 20383
rect 3099 20380 3111 20383
rect 3160 20380 3188 20556
rect 4525 20519 4583 20525
rect 4525 20485 4537 20519
rect 4571 20516 4583 20519
rect 5074 20516 5080 20528
rect 4571 20488 5080 20516
rect 4571 20485 4583 20488
rect 4525 20479 4583 20485
rect 5074 20476 5080 20488
rect 5132 20476 5138 20528
rect 5258 20476 5264 20528
rect 5316 20516 5322 20528
rect 6748 20516 6776 20556
rect 7285 20553 7297 20587
rect 7331 20584 7343 20587
rect 9858 20584 9864 20596
rect 7331 20556 9864 20584
rect 7331 20553 7343 20556
rect 7285 20547 7343 20553
rect 9858 20544 9864 20556
rect 9916 20544 9922 20596
rect 18138 20544 18144 20596
rect 18196 20584 18202 20596
rect 19061 20587 19119 20593
rect 19061 20584 19073 20587
rect 18196 20556 19073 20584
rect 18196 20544 18202 20556
rect 19061 20553 19073 20556
rect 19107 20553 19119 20587
rect 19061 20547 19119 20553
rect 19613 20587 19671 20593
rect 19613 20553 19625 20587
rect 19659 20584 19671 20587
rect 21634 20584 21640 20596
rect 19659 20556 21640 20584
rect 19659 20553 19671 20556
rect 19613 20547 19671 20553
rect 21634 20544 21640 20556
rect 21692 20544 21698 20596
rect 5316 20488 6684 20516
rect 6748 20488 8984 20516
rect 5316 20476 5322 20488
rect 3513 20451 3571 20457
rect 3513 20417 3525 20451
rect 3559 20448 3571 20451
rect 4430 20448 4436 20460
rect 3559 20420 4436 20448
rect 3559 20417 3571 20420
rect 3513 20411 3571 20417
rect 4430 20408 4436 20420
rect 4488 20408 4494 20460
rect 6656 20457 6684 20488
rect 5905 20451 5963 20457
rect 5905 20448 5917 20451
rect 4724 20420 5917 20448
rect 3099 20352 3188 20380
rect 3099 20349 3111 20352
rect 3053 20343 3111 20349
rect 3234 20340 3240 20392
rect 3292 20380 3298 20392
rect 3329 20383 3387 20389
rect 3329 20380 3341 20383
rect 3292 20352 3341 20380
rect 3292 20340 3298 20352
rect 3329 20349 3341 20352
rect 3375 20380 3387 20383
rect 3605 20383 3663 20389
rect 3605 20380 3617 20383
rect 3375 20352 3617 20380
rect 3375 20349 3387 20352
rect 3329 20343 3387 20349
rect 3605 20349 3617 20352
rect 3651 20349 3663 20383
rect 3605 20343 3663 20349
rect 3694 20340 3700 20392
rect 3752 20380 3758 20392
rect 3973 20383 4031 20389
rect 3973 20380 3985 20383
rect 3752 20352 3985 20380
rect 3752 20340 3758 20352
rect 3973 20349 3985 20352
rect 4019 20380 4031 20383
rect 4617 20383 4675 20389
rect 4617 20380 4629 20383
rect 4019 20352 4629 20380
rect 4019 20349 4031 20352
rect 3973 20343 4031 20349
rect 4617 20349 4629 20352
rect 4663 20349 4675 20383
rect 4617 20343 4675 20349
rect 1578 20312 1584 20324
rect 1539 20284 1584 20312
rect 1578 20272 1584 20284
rect 1636 20272 1642 20324
rect 1949 20315 2007 20321
rect 1949 20281 1961 20315
rect 1995 20312 2007 20315
rect 2130 20312 2136 20324
rect 1995 20284 2136 20312
rect 1995 20281 2007 20284
rect 1949 20275 2007 20281
rect 2130 20272 2136 20284
rect 2188 20272 2194 20324
rect 2314 20312 2320 20324
rect 2275 20284 2320 20312
rect 2314 20272 2320 20284
rect 2372 20272 2378 20324
rect 2590 20272 2596 20324
rect 2648 20312 2654 20324
rect 2685 20315 2743 20321
rect 2685 20312 2697 20315
rect 2648 20284 2697 20312
rect 2648 20272 2654 20284
rect 2685 20281 2697 20284
rect 2731 20281 2743 20315
rect 4341 20315 4399 20321
rect 4341 20312 4353 20315
rect 2685 20275 2743 20281
rect 3988 20284 4353 20312
rect 3988 20256 4016 20284
rect 4341 20281 4353 20284
rect 4387 20312 4399 20315
rect 4724 20312 4752 20420
rect 5905 20417 5917 20420
rect 5951 20417 5963 20451
rect 5905 20411 5963 20417
rect 6641 20451 6699 20457
rect 6641 20417 6653 20451
rect 6687 20417 6699 20451
rect 8956 20448 8984 20488
rect 9030 20476 9036 20528
rect 9088 20516 9094 20528
rect 10686 20516 10692 20528
rect 9088 20488 10692 20516
rect 9088 20476 9094 20488
rect 10686 20476 10692 20488
rect 10744 20476 10750 20528
rect 10870 20516 10876 20528
rect 10831 20488 10876 20516
rect 10870 20476 10876 20488
rect 10928 20476 10934 20528
rect 11238 20516 11244 20528
rect 11199 20488 11244 20516
rect 11238 20476 11244 20488
rect 11296 20476 11302 20528
rect 11698 20476 11704 20528
rect 11756 20516 11762 20528
rect 11885 20519 11943 20525
rect 11885 20516 11897 20519
rect 11756 20488 11897 20516
rect 11756 20476 11762 20488
rect 11885 20485 11897 20488
rect 11931 20485 11943 20519
rect 11885 20479 11943 20485
rect 12066 20476 12072 20528
rect 12124 20516 12130 20528
rect 12253 20519 12311 20525
rect 12253 20516 12265 20519
rect 12124 20488 12265 20516
rect 12124 20476 12130 20488
rect 12253 20485 12265 20488
rect 12299 20485 12311 20519
rect 12253 20479 12311 20485
rect 12434 20476 12440 20528
rect 12492 20516 12498 20528
rect 12621 20519 12679 20525
rect 12621 20516 12633 20519
rect 12492 20488 12633 20516
rect 12492 20476 12498 20488
rect 12621 20485 12633 20488
rect 12667 20485 12679 20519
rect 12621 20479 12679 20485
rect 12802 20476 12808 20528
rect 12860 20516 12866 20528
rect 12989 20519 13047 20525
rect 12989 20516 13001 20519
rect 12860 20488 13001 20516
rect 12860 20476 12866 20488
rect 12989 20485 13001 20488
rect 13035 20485 13047 20519
rect 12989 20479 13047 20485
rect 13170 20476 13176 20528
rect 13228 20516 13234 20528
rect 13357 20519 13415 20525
rect 13357 20516 13369 20519
rect 13228 20488 13369 20516
rect 13228 20476 13234 20488
rect 13357 20485 13369 20488
rect 13403 20485 13415 20519
rect 13357 20479 13415 20485
rect 13538 20476 13544 20528
rect 13596 20516 13602 20528
rect 13725 20519 13783 20525
rect 13725 20516 13737 20519
rect 13596 20488 13737 20516
rect 13596 20476 13602 20488
rect 13725 20485 13737 20488
rect 13771 20485 13783 20519
rect 13725 20479 13783 20485
rect 13998 20476 14004 20528
rect 14056 20516 14062 20528
rect 14093 20519 14151 20525
rect 14093 20516 14105 20519
rect 14056 20488 14105 20516
rect 14056 20476 14062 20488
rect 14093 20485 14105 20488
rect 14139 20485 14151 20519
rect 14734 20516 14740 20528
rect 14695 20488 14740 20516
rect 14093 20479 14151 20485
rect 14734 20476 14740 20488
rect 14792 20476 14798 20528
rect 15102 20516 15108 20528
rect 15063 20488 15108 20516
rect 15102 20476 15108 20488
rect 15160 20476 15166 20528
rect 15470 20516 15476 20528
rect 15431 20488 15476 20516
rect 15470 20476 15476 20488
rect 15528 20476 15534 20528
rect 15838 20516 15844 20528
rect 15799 20488 15844 20516
rect 15838 20476 15844 20488
rect 15896 20476 15902 20528
rect 16298 20516 16304 20528
rect 16259 20488 16304 20516
rect 16298 20476 16304 20488
rect 16356 20476 16362 20528
rect 16666 20516 16672 20528
rect 16627 20488 16672 20516
rect 16666 20476 16672 20488
rect 16724 20476 16730 20528
rect 17034 20476 17040 20528
rect 17092 20516 17098 20528
rect 17221 20519 17279 20525
rect 17221 20516 17233 20519
rect 17092 20488 17233 20516
rect 17092 20476 17098 20488
rect 17221 20485 17233 20488
rect 17267 20485 17279 20519
rect 17221 20479 17279 20485
rect 17402 20476 17408 20528
rect 17460 20516 17466 20528
rect 17589 20519 17647 20525
rect 17589 20516 17601 20519
rect 17460 20488 17601 20516
rect 17460 20476 17466 20488
rect 17589 20485 17601 20488
rect 17635 20485 17647 20519
rect 17954 20516 17960 20528
rect 17915 20488 17960 20516
rect 17589 20479 17647 20485
rect 17954 20476 17960 20488
rect 18012 20476 18018 20528
rect 18598 20516 18604 20528
rect 18559 20488 18604 20516
rect 18598 20476 18604 20488
rect 18656 20476 18662 20528
rect 20438 20516 20444 20528
rect 20399 20488 20444 20516
rect 20438 20476 20444 20488
rect 20496 20476 20502 20528
rect 20530 20476 20536 20528
rect 20588 20476 20594 20528
rect 20806 20516 20812 20528
rect 20767 20488 20812 20516
rect 20806 20476 20812 20488
rect 20864 20476 20870 20528
rect 18138 20448 18144 20460
rect 6641 20411 6699 20417
rect 8036 20420 8892 20448
rect 8956 20420 10916 20448
rect 4798 20340 4804 20392
rect 4856 20380 4862 20392
rect 4893 20383 4951 20389
rect 4893 20380 4905 20383
rect 4856 20352 4905 20380
rect 4856 20340 4862 20352
rect 4893 20349 4905 20352
rect 4939 20349 4951 20383
rect 4893 20343 4951 20349
rect 5166 20340 5172 20392
rect 5224 20380 5230 20392
rect 5353 20383 5411 20389
rect 5353 20380 5365 20383
rect 5224 20352 5365 20380
rect 5224 20340 5230 20352
rect 5353 20349 5365 20352
rect 5399 20349 5411 20383
rect 5353 20343 5411 20349
rect 5537 20383 5595 20389
rect 5537 20349 5549 20383
rect 5583 20380 5595 20383
rect 5626 20380 5632 20392
rect 5583 20352 5632 20380
rect 5583 20349 5595 20352
rect 5537 20343 5595 20349
rect 5626 20340 5632 20352
rect 5684 20340 5690 20392
rect 5721 20383 5779 20389
rect 5721 20349 5733 20383
rect 5767 20380 5779 20383
rect 5994 20380 6000 20392
rect 5767 20352 6000 20380
rect 5767 20349 5779 20352
rect 5721 20343 5779 20349
rect 5994 20340 6000 20352
rect 6052 20340 6058 20392
rect 6181 20383 6239 20389
rect 6181 20349 6193 20383
rect 6227 20380 6239 20383
rect 6270 20380 6276 20392
rect 6227 20352 6276 20380
rect 6227 20349 6239 20352
rect 6181 20343 6239 20349
rect 6270 20340 6276 20352
rect 6328 20340 6334 20392
rect 6362 20340 6368 20392
rect 6420 20380 6426 20392
rect 6420 20352 6465 20380
rect 6665 20352 7052 20380
rect 6420 20340 6426 20352
rect 4387 20284 4752 20312
rect 5077 20315 5135 20321
rect 4387 20281 4399 20284
rect 4341 20275 4399 20281
rect 5077 20281 5089 20315
rect 5123 20312 5135 20315
rect 5123 20284 5396 20312
rect 5123 20281 5135 20284
rect 5077 20275 5135 20281
rect 1486 20244 1492 20256
rect 1447 20216 1492 20244
rect 1486 20204 1492 20216
rect 1544 20204 1550 20256
rect 2498 20204 2504 20256
rect 2556 20244 2562 20256
rect 3326 20244 3332 20256
rect 2556 20216 3332 20244
rect 2556 20204 2562 20216
rect 3326 20204 3332 20216
rect 3384 20204 3390 20256
rect 3970 20204 3976 20256
rect 4028 20204 4034 20256
rect 4065 20247 4123 20253
rect 4065 20213 4077 20247
rect 4111 20244 4123 20247
rect 4706 20244 4712 20256
rect 4111 20216 4712 20244
rect 4111 20213 4123 20216
rect 4065 20207 4123 20213
rect 4706 20204 4712 20216
rect 4764 20204 4770 20256
rect 4890 20204 4896 20256
rect 4948 20244 4954 20256
rect 5261 20247 5319 20253
rect 5261 20244 5273 20247
rect 4948 20216 5273 20244
rect 4948 20204 4954 20216
rect 5261 20213 5273 20216
rect 5307 20213 5319 20247
rect 5368 20244 5396 20284
rect 5442 20272 5448 20324
rect 5500 20312 5506 20324
rect 6665 20312 6693 20352
rect 5500 20284 6693 20312
rect 5500 20272 5506 20284
rect 6730 20272 6736 20324
rect 6788 20312 6794 20324
rect 6917 20315 6975 20321
rect 6917 20312 6929 20315
rect 6788 20284 6929 20312
rect 6788 20272 6794 20284
rect 6917 20281 6929 20284
rect 6963 20281 6975 20315
rect 7024 20312 7052 20352
rect 7098 20340 7104 20392
rect 7156 20380 7162 20392
rect 7561 20383 7619 20389
rect 7561 20380 7573 20383
rect 7156 20352 7573 20380
rect 7156 20340 7162 20352
rect 7561 20349 7573 20352
rect 7607 20349 7619 20383
rect 7561 20343 7619 20349
rect 7834 20340 7840 20392
rect 7892 20380 7898 20392
rect 8036 20389 8064 20420
rect 8021 20383 8079 20389
rect 8021 20380 8033 20383
rect 7892 20352 8033 20380
rect 7892 20340 7898 20352
rect 8021 20349 8033 20352
rect 8067 20349 8079 20383
rect 8021 20343 8079 20349
rect 8110 20340 8116 20392
rect 8168 20380 8174 20392
rect 8205 20383 8263 20389
rect 8205 20380 8217 20383
rect 8168 20352 8217 20380
rect 8168 20340 8174 20352
rect 8205 20349 8217 20352
rect 8251 20349 8263 20383
rect 8205 20343 8263 20349
rect 8294 20340 8300 20392
rect 8352 20380 8358 20392
rect 8389 20383 8447 20389
rect 8389 20380 8401 20383
rect 8352 20352 8401 20380
rect 8352 20340 8358 20352
rect 8389 20349 8401 20352
rect 8435 20349 8447 20383
rect 8754 20380 8760 20392
rect 8715 20352 8760 20380
rect 8389 20343 8447 20349
rect 8754 20340 8760 20352
rect 8812 20340 8818 20392
rect 8864 20380 8892 20420
rect 9217 20383 9275 20389
rect 9217 20380 9229 20383
rect 8864 20352 9229 20380
rect 9217 20349 9229 20352
rect 9263 20349 9275 20383
rect 9217 20343 9275 20349
rect 9398 20340 9404 20392
rect 9456 20380 9462 20392
rect 9585 20383 9643 20389
rect 9585 20380 9597 20383
rect 9456 20352 9597 20380
rect 9456 20340 9462 20352
rect 9585 20349 9597 20352
rect 9631 20349 9643 20383
rect 9585 20343 9643 20349
rect 9766 20340 9772 20392
rect 9824 20380 9830 20392
rect 9953 20383 10011 20389
rect 9953 20380 9965 20383
rect 9824 20352 9965 20380
rect 9824 20340 9830 20352
rect 9953 20349 9965 20352
rect 9999 20349 10011 20383
rect 9953 20343 10011 20349
rect 10134 20340 10140 20392
rect 10192 20380 10198 20392
rect 10321 20383 10379 20389
rect 10321 20380 10333 20383
rect 10192 20352 10333 20380
rect 10192 20340 10198 20352
rect 10321 20349 10333 20352
rect 10367 20349 10379 20383
rect 10686 20380 10692 20392
rect 10647 20352 10692 20380
rect 10321 20343 10379 20349
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 7282 20312 7288 20324
rect 7024 20284 7288 20312
rect 6917 20275 6975 20281
rect 7282 20272 7288 20284
rect 7340 20272 7346 20324
rect 8846 20272 8852 20324
rect 8904 20312 8910 20324
rect 8941 20315 8999 20321
rect 8941 20312 8953 20315
rect 8904 20284 8953 20312
rect 8904 20272 8910 20284
rect 8941 20281 8953 20284
rect 8987 20281 8999 20315
rect 8941 20275 8999 20281
rect 9674 20272 9680 20324
rect 9732 20312 9738 20324
rect 9732 20284 10272 20312
rect 9732 20272 9738 20284
rect 6086 20244 6092 20256
rect 5368 20216 6092 20244
rect 5261 20207 5319 20213
rect 6086 20204 6092 20216
rect 6144 20204 6150 20256
rect 6825 20247 6883 20253
rect 6825 20213 6837 20247
rect 6871 20244 6883 20247
rect 7190 20244 7196 20256
rect 6871 20216 7196 20244
rect 6871 20213 6883 20216
rect 6825 20207 6883 20213
rect 7190 20204 7196 20216
rect 7248 20204 7254 20256
rect 7469 20247 7527 20253
rect 7469 20213 7481 20247
rect 7515 20244 7527 20247
rect 7742 20244 7748 20256
rect 7515 20216 7748 20244
rect 7515 20213 7527 20216
rect 7469 20207 7527 20213
rect 7742 20204 7748 20216
rect 7800 20204 7806 20256
rect 7929 20247 7987 20253
rect 7929 20213 7941 20247
rect 7975 20244 7987 20247
rect 8478 20244 8484 20256
rect 7975 20216 8484 20244
rect 7975 20213 7987 20216
rect 7929 20207 7987 20213
rect 8478 20204 8484 20216
rect 8536 20204 8542 20256
rect 8662 20244 8668 20256
rect 8623 20216 8668 20244
rect 8662 20204 8668 20216
rect 8720 20204 8726 20256
rect 9490 20244 9496 20256
rect 9451 20216 9496 20244
rect 9490 20204 9496 20216
rect 9548 20204 9554 20256
rect 9861 20247 9919 20253
rect 9861 20213 9873 20247
rect 9907 20244 9919 20247
rect 9950 20244 9956 20256
rect 9907 20216 9956 20244
rect 9907 20213 9919 20216
rect 9861 20207 9919 20213
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 10244 20253 10272 20284
rect 10229 20247 10287 20253
rect 10229 20213 10241 20247
rect 10275 20213 10287 20247
rect 10229 20207 10287 20213
rect 10505 20247 10563 20253
rect 10505 20213 10517 20247
rect 10551 20244 10563 20247
rect 10778 20244 10784 20256
rect 10551 20216 10784 20244
rect 10551 20213 10563 20216
rect 10505 20207 10563 20213
rect 10778 20204 10784 20216
rect 10836 20204 10842 20256
rect 10888 20244 10916 20420
rect 17880 20420 18144 20448
rect 17880 20392 17908 20420
rect 18138 20408 18144 20420
rect 18196 20448 18202 20460
rect 19702 20448 19708 20460
rect 18196 20420 19708 20448
rect 18196 20408 18202 20420
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 17862 20340 17868 20392
rect 17920 20340 17926 20392
rect 18325 20383 18383 20389
rect 18325 20349 18337 20383
rect 18371 20380 18383 20383
rect 18966 20380 18972 20392
rect 18371 20352 18972 20380
rect 18371 20349 18383 20352
rect 18325 20343 18383 20349
rect 18966 20340 18972 20352
rect 19024 20340 19030 20392
rect 19150 20380 19156 20392
rect 19111 20352 19156 20380
rect 19150 20340 19156 20352
rect 19208 20340 19214 20392
rect 19334 20340 19340 20392
rect 19392 20380 19398 20392
rect 19889 20383 19947 20389
rect 19889 20380 19901 20383
rect 19392 20352 19901 20380
rect 19392 20340 19398 20352
rect 19889 20349 19901 20352
rect 19935 20349 19947 20383
rect 20254 20380 20260 20392
rect 20215 20352 20260 20380
rect 19889 20343 19947 20349
rect 20254 20340 20260 20352
rect 20312 20340 20318 20392
rect 20548 20380 20576 20476
rect 21174 20448 21180 20460
rect 21135 20420 21180 20448
rect 21174 20408 21180 20420
rect 21232 20408 21238 20460
rect 20608 20383 20666 20389
rect 20608 20380 20620 20383
rect 20548 20352 20620 20380
rect 20608 20349 20620 20352
rect 20654 20349 20666 20383
rect 20990 20380 20996 20392
rect 20951 20352 20996 20380
rect 20608 20343 20666 20349
rect 20990 20340 20996 20352
rect 21048 20340 21054 20392
rect 22370 20380 22376 20392
rect 21100 20352 22376 20380
rect 11054 20312 11060 20324
rect 11015 20284 11060 20312
rect 11054 20272 11060 20284
rect 11112 20272 11118 20324
rect 11422 20312 11428 20324
rect 11383 20284 11428 20312
rect 11422 20272 11428 20284
rect 11480 20272 11486 20324
rect 12066 20312 12072 20324
rect 12027 20284 12072 20312
rect 12066 20272 12072 20284
rect 12124 20272 12130 20324
rect 12434 20272 12440 20324
rect 12492 20312 12498 20324
rect 12802 20312 12808 20324
rect 12492 20284 12537 20312
rect 12763 20284 12808 20312
rect 12492 20272 12498 20284
rect 12802 20272 12808 20284
rect 12860 20272 12866 20324
rect 13170 20312 13176 20324
rect 13131 20284 13176 20312
rect 13170 20272 13176 20284
rect 13228 20272 13234 20324
rect 13538 20312 13544 20324
rect 13499 20284 13544 20312
rect 13538 20272 13544 20284
rect 13596 20272 13602 20324
rect 13814 20272 13820 20324
rect 13872 20312 13878 20324
rect 13909 20315 13967 20321
rect 13909 20312 13921 20315
rect 13872 20284 13921 20312
rect 13872 20272 13878 20284
rect 13909 20281 13921 20284
rect 13955 20281 13967 20315
rect 14274 20312 14280 20324
rect 14235 20284 14280 20312
rect 13909 20275 13967 20281
rect 14274 20272 14280 20284
rect 14332 20272 14338 20324
rect 14642 20272 14648 20324
rect 14700 20312 14706 20324
rect 14921 20315 14979 20321
rect 14921 20312 14933 20315
rect 14700 20284 14933 20312
rect 14700 20272 14706 20284
rect 14921 20281 14933 20284
rect 14967 20281 14979 20315
rect 14921 20275 14979 20281
rect 15194 20272 15200 20324
rect 15252 20312 15258 20324
rect 15289 20315 15347 20321
rect 15289 20312 15301 20315
rect 15252 20284 15301 20312
rect 15252 20272 15258 20284
rect 15289 20281 15301 20284
rect 15335 20281 15347 20315
rect 15654 20312 15660 20324
rect 15615 20284 15660 20312
rect 15289 20275 15347 20281
rect 15654 20272 15660 20284
rect 15712 20272 15718 20324
rect 16022 20312 16028 20324
rect 15983 20284 16028 20312
rect 16022 20272 16028 20284
rect 16080 20272 16086 20324
rect 16482 20312 16488 20324
rect 16443 20284 16488 20312
rect 16482 20272 16488 20284
rect 16540 20272 16546 20324
rect 16850 20312 16856 20324
rect 16811 20284 16856 20312
rect 16850 20272 16856 20284
rect 16908 20272 16914 20324
rect 17402 20312 17408 20324
rect 17363 20284 17408 20312
rect 17402 20272 17408 20284
rect 17460 20272 17466 20324
rect 17770 20312 17776 20324
rect 17731 20284 17776 20312
rect 17770 20272 17776 20284
rect 17828 20272 17834 20324
rect 17954 20272 17960 20324
rect 18012 20312 18018 20324
rect 18141 20315 18199 20321
rect 18141 20312 18153 20315
rect 18012 20284 18153 20312
rect 18012 20272 18018 20284
rect 18141 20281 18153 20284
rect 18187 20281 18199 20315
rect 18785 20315 18843 20321
rect 18141 20275 18199 20281
rect 18248 20284 18644 20312
rect 15930 20244 15936 20256
rect 10888 20216 15936 20244
rect 15930 20204 15936 20216
rect 15988 20204 15994 20256
rect 17218 20204 17224 20256
rect 17276 20244 17282 20256
rect 18248 20244 18276 20284
rect 18506 20244 18512 20256
rect 17276 20216 18276 20244
rect 18467 20216 18512 20244
rect 17276 20204 17282 20216
rect 18506 20204 18512 20216
rect 18564 20204 18570 20256
rect 18616 20244 18644 20284
rect 18785 20281 18797 20315
rect 18831 20312 18843 20315
rect 18874 20312 18880 20324
rect 18831 20284 18880 20312
rect 18831 20281 18843 20284
rect 18785 20275 18843 20281
rect 18874 20272 18880 20284
rect 18932 20272 18938 20324
rect 19518 20312 19524 20324
rect 18984 20284 19334 20312
rect 19479 20284 19524 20312
rect 18984 20244 19012 20284
rect 18616 20216 19012 20244
rect 19306 20244 19334 20284
rect 19518 20272 19524 20284
rect 19576 20272 19582 20324
rect 21100 20312 21128 20352
rect 22370 20340 22376 20352
rect 22428 20340 22434 20392
rect 19628 20284 21128 20312
rect 21361 20315 21419 20321
rect 19628 20244 19656 20284
rect 21361 20281 21373 20315
rect 21407 20281 21419 20315
rect 21542 20312 21548 20324
rect 21503 20284 21548 20312
rect 21361 20275 21419 20281
rect 20070 20244 20076 20256
rect 19306 20216 19656 20244
rect 20031 20216 20076 20244
rect 20070 20204 20076 20216
rect 20128 20204 20134 20256
rect 20162 20204 20168 20256
rect 20220 20244 20226 20256
rect 21376 20244 21404 20275
rect 21542 20272 21548 20284
rect 21600 20272 21606 20324
rect 20220 20216 21404 20244
rect 20220 20204 20226 20216
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 1394 20000 1400 20052
rect 1452 20040 1458 20052
rect 1857 20043 1915 20049
rect 1857 20040 1869 20043
rect 1452 20012 1869 20040
rect 1452 20000 1458 20012
rect 1857 20009 1869 20012
rect 1903 20009 1915 20043
rect 1857 20003 1915 20009
rect 2038 20000 2044 20052
rect 2096 20040 2102 20052
rect 3050 20040 3056 20052
rect 2096 20012 3056 20040
rect 2096 20000 2102 20012
rect 3050 20000 3056 20012
rect 3108 20000 3114 20052
rect 3234 20000 3240 20052
rect 3292 20040 3298 20052
rect 5442 20040 5448 20052
rect 3292 20012 5448 20040
rect 3292 20000 3298 20012
rect 5442 20000 5448 20012
rect 5500 20000 5506 20052
rect 5629 20043 5687 20049
rect 5629 20009 5641 20043
rect 5675 20040 5687 20043
rect 7006 20040 7012 20052
rect 5675 20012 7012 20040
rect 5675 20009 5687 20012
rect 5629 20003 5687 20009
rect 7006 20000 7012 20012
rect 7064 20000 7070 20052
rect 7282 20000 7288 20052
rect 7340 20040 7346 20052
rect 8113 20043 8171 20049
rect 8113 20040 8125 20043
rect 7340 20012 8125 20040
rect 7340 20000 7346 20012
rect 8113 20009 8125 20012
rect 8159 20009 8171 20043
rect 8113 20003 8171 20009
rect 8754 20000 8760 20052
rect 8812 20040 8818 20052
rect 9309 20043 9367 20049
rect 9309 20040 9321 20043
rect 8812 20012 9321 20040
rect 8812 20000 8818 20012
rect 9309 20009 9321 20012
rect 9355 20009 9367 20043
rect 9309 20003 9367 20009
rect 9398 20000 9404 20052
rect 9456 20040 9462 20052
rect 9769 20043 9827 20049
rect 9769 20040 9781 20043
rect 9456 20012 9781 20040
rect 9456 20000 9462 20012
rect 9769 20009 9781 20012
rect 9815 20009 9827 20043
rect 9769 20003 9827 20009
rect 10505 20043 10563 20049
rect 10505 20009 10517 20043
rect 10551 20040 10563 20043
rect 11422 20040 11428 20052
rect 10551 20012 11428 20040
rect 10551 20009 10563 20012
rect 10505 20003 10563 20009
rect 11422 20000 11428 20012
rect 11480 20000 11486 20052
rect 11609 20043 11667 20049
rect 11609 20009 11621 20043
rect 11655 20040 11667 20043
rect 12802 20040 12808 20052
rect 11655 20012 12808 20040
rect 11655 20009 11667 20012
rect 11609 20003 11667 20009
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 16761 20043 16819 20049
rect 16761 20009 16773 20043
rect 16807 20040 16819 20043
rect 16942 20040 16948 20052
rect 16807 20012 16948 20040
rect 16807 20009 16819 20012
rect 16761 20003 16819 20009
rect 16942 20000 16948 20012
rect 17000 20000 17006 20052
rect 17218 20040 17224 20052
rect 17179 20012 17224 20040
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 18325 20043 18383 20049
rect 17420 20012 18276 20040
rect 1581 19975 1639 19981
rect 1581 19941 1593 19975
rect 1627 19972 1639 19975
rect 2222 19972 2228 19984
rect 1627 19944 2228 19972
rect 1627 19941 1639 19944
rect 1581 19935 1639 19941
rect 2222 19932 2228 19944
rect 2280 19932 2286 19984
rect 3878 19972 3884 19984
rect 2516 19944 3884 19972
rect 1949 19907 2007 19913
rect 1949 19873 1961 19907
rect 1995 19904 2007 19907
rect 2038 19904 2044 19916
rect 1995 19876 2044 19904
rect 1995 19873 2007 19876
rect 1949 19867 2007 19873
rect 2038 19864 2044 19876
rect 2096 19864 2102 19916
rect 2133 19907 2191 19913
rect 2133 19873 2145 19907
rect 2179 19873 2191 19907
rect 2406 19904 2412 19916
rect 2367 19876 2412 19904
rect 2133 19867 2191 19873
rect 198 19796 204 19848
rect 256 19836 262 19848
rect 1762 19836 1768 19848
rect 256 19808 1768 19836
rect 256 19796 262 19808
rect 1762 19796 1768 19808
rect 1820 19836 1826 19848
rect 2148 19836 2176 19867
rect 2406 19864 2412 19876
rect 2464 19864 2470 19916
rect 2516 19836 2544 19944
rect 3878 19932 3884 19944
rect 3936 19932 3942 19984
rect 3970 19932 3976 19984
rect 4028 19972 4034 19984
rect 4028 19944 5488 19972
rect 4028 19932 4034 19944
rect 2682 19904 2688 19916
rect 2643 19876 2688 19904
rect 2682 19864 2688 19876
rect 2740 19864 2746 19916
rect 2953 19907 3011 19913
rect 2953 19873 2965 19907
rect 2999 19904 3011 19907
rect 3050 19904 3056 19916
rect 2999 19876 3056 19904
rect 2999 19873 3011 19876
rect 2953 19867 3011 19873
rect 3050 19864 3056 19876
rect 3108 19864 3114 19916
rect 3237 19907 3295 19913
rect 3237 19873 3249 19907
rect 3283 19904 3295 19907
rect 3326 19904 3332 19916
rect 3283 19876 3332 19904
rect 3283 19873 3295 19876
rect 3237 19867 3295 19873
rect 3326 19864 3332 19876
rect 3384 19864 3390 19916
rect 3513 19907 3571 19913
rect 3513 19873 3525 19907
rect 3559 19904 3571 19907
rect 3694 19904 3700 19916
rect 3559 19876 3700 19904
rect 3559 19873 3571 19876
rect 3513 19867 3571 19873
rect 3694 19864 3700 19876
rect 3752 19904 3758 19916
rect 4062 19904 4068 19916
rect 3752 19876 4068 19904
rect 3752 19864 3758 19876
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 5097 19907 5155 19913
rect 5097 19873 5109 19907
rect 5143 19904 5155 19907
rect 5258 19904 5264 19916
rect 5143 19876 5264 19904
rect 5143 19873 5155 19876
rect 5097 19867 5155 19873
rect 5258 19864 5264 19876
rect 5316 19864 5322 19916
rect 5460 19913 5488 19944
rect 5534 19932 5540 19984
rect 5592 19972 5598 19984
rect 5994 19972 6000 19984
rect 5592 19944 6000 19972
rect 5592 19932 5598 19944
rect 5994 19932 6000 19944
rect 6052 19932 6058 19984
rect 6638 19932 6644 19984
rect 6696 19972 6702 19984
rect 7098 19972 7104 19984
rect 6696 19944 7104 19972
rect 6696 19932 6702 19944
rect 7098 19932 7104 19944
rect 7156 19972 7162 19984
rect 7377 19975 7435 19981
rect 7377 19972 7389 19975
rect 7156 19944 7389 19972
rect 7156 19932 7162 19944
rect 7377 19941 7389 19944
rect 7423 19941 7435 19975
rect 7377 19935 7435 19941
rect 7466 19932 7472 19984
rect 7524 19972 7530 19984
rect 7524 19944 8156 19972
rect 7524 19932 7530 19944
rect 5445 19907 5503 19913
rect 5445 19873 5457 19907
rect 5491 19873 5503 19907
rect 5445 19867 5503 19873
rect 6080 19907 6138 19913
rect 6080 19873 6092 19907
rect 6126 19904 6138 19907
rect 6546 19904 6552 19916
rect 6126 19876 6552 19904
rect 6126 19873 6138 19876
rect 6080 19867 6138 19873
rect 6546 19864 6552 19876
rect 6604 19904 6610 19916
rect 6822 19904 6828 19916
rect 6604 19876 6828 19904
rect 6604 19864 6610 19876
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 8021 19907 8079 19913
rect 8021 19873 8033 19907
rect 8067 19873 8079 19907
rect 8128 19904 8156 19944
rect 8294 19932 8300 19984
rect 8352 19972 8358 19984
rect 9125 19975 9183 19981
rect 9125 19972 9137 19975
rect 8352 19944 9137 19972
rect 8352 19932 8358 19944
rect 9125 19941 9137 19944
rect 9171 19941 9183 19975
rect 11333 19975 11391 19981
rect 11333 19972 11345 19975
rect 9125 19935 9183 19941
rect 10796 19944 11345 19972
rect 8665 19907 8723 19913
rect 8665 19904 8677 19907
rect 8128 19876 8677 19904
rect 8021 19867 8079 19873
rect 8665 19873 8677 19876
rect 8711 19904 8723 19907
rect 8757 19907 8815 19913
rect 8757 19904 8769 19907
rect 8711 19876 8769 19904
rect 8711 19873 8723 19876
rect 8665 19867 8723 19873
rect 8757 19873 8769 19876
rect 8803 19873 8815 19907
rect 8757 19867 8815 19873
rect 1820 19808 2176 19836
rect 2332 19808 2544 19836
rect 5353 19839 5411 19845
rect 1820 19796 1826 19808
rect 2332 19777 2360 19808
rect 5353 19805 5365 19839
rect 5399 19836 5411 19839
rect 5718 19836 5724 19848
rect 5399 19808 5724 19836
rect 5399 19805 5411 19808
rect 5353 19799 5411 19805
rect 5718 19796 5724 19808
rect 5776 19836 5782 19848
rect 5813 19839 5871 19845
rect 5813 19836 5825 19839
rect 5776 19808 5825 19836
rect 5776 19796 5782 19808
rect 5813 19805 5825 19808
rect 5859 19805 5871 19839
rect 5813 19799 5871 19805
rect 7374 19796 7380 19848
rect 7432 19836 7438 19848
rect 8036 19836 8064 19867
rect 9766 19864 9772 19916
rect 9824 19904 9830 19916
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9824 19876 10149 19904
rect 9824 19864 9830 19876
rect 10137 19873 10149 19876
rect 10183 19873 10195 19907
rect 10318 19904 10324 19916
rect 10279 19876 10324 19904
rect 10137 19867 10195 19873
rect 10318 19864 10324 19876
rect 10376 19864 10382 19916
rect 10502 19864 10508 19916
rect 10560 19904 10566 19916
rect 10796 19913 10824 19944
rect 11333 19941 11345 19944
rect 11379 19941 11391 19975
rect 14366 19972 14372 19984
rect 14327 19944 14372 19972
rect 11333 19935 11391 19941
rect 14366 19932 14372 19944
rect 14424 19932 14430 19984
rect 10781 19907 10839 19913
rect 10781 19904 10793 19907
rect 10560 19876 10793 19904
rect 10560 19864 10566 19876
rect 10781 19873 10793 19876
rect 10827 19873 10839 19907
rect 10781 19867 10839 19873
rect 11238 19864 11244 19916
rect 11296 19904 11302 19916
rect 11425 19907 11483 19913
rect 11425 19904 11437 19907
rect 11296 19876 11437 19904
rect 11296 19864 11302 19876
rect 11425 19873 11437 19876
rect 11471 19873 11483 19907
rect 11425 19867 11483 19873
rect 12161 19907 12219 19913
rect 12161 19873 12173 19907
rect 12207 19904 12219 19907
rect 12526 19904 12532 19916
rect 12207 19876 12532 19904
rect 12207 19873 12219 19876
rect 12161 19867 12219 19873
rect 12526 19864 12532 19876
rect 12584 19864 12590 19916
rect 14550 19904 14556 19916
rect 14511 19876 14556 19904
rect 14550 19864 14556 19876
rect 14608 19864 14614 19916
rect 17034 19904 17040 19916
rect 16995 19876 17040 19904
rect 17034 19864 17040 19876
rect 17092 19864 17098 19916
rect 17310 19904 17316 19916
rect 17271 19876 17316 19904
rect 17310 19864 17316 19876
rect 17368 19864 17374 19916
rect 7432 19808 8064 19836
rect 7432 19796 7438 19808
rect 8110 19796 8116 19848
rect 8168 19836 8174 19848
rect 8205 19839 8263 19845
rect 8205 19836 8217 19839
rect 8168 19808 8217 19836
rect 8168 19796 8174 19808
rect 8205 19805 8217 19808
rect 8251 19805 8263 19839
rect 17420 19836 17448 20012
rect 18248 19972 18276 20012
rect 18325 20009 18337 20043
rect 18371 20040 18383 20043
rect 18371 20012 18644 20040
rect 18371 20009 18383 20012
rect 18325 20003 18383 20009
rect 18248 19944 18460 19972
rect 17589 19907 17647 19913
rect 17589 19873 17601 19907
rect 17635 19904 17647 19907
rect 17678 19904 17684 19916
rect 17635 19876 17684 19904
rect 17635 19873 17647 19876
rect 17589 19867 17647 19873
rect 17678 19864 17684 19876
rect 17736 19864 17742 19916
rect 17862 19904 17868 19916
rect 17823 19876 17868 19904
rect 17862 19864 17868 19876
rect 17920 19864 17926 19916
rect 18046 19864 18052 19916
rect 18104 19904 18110 19916
rect 18141 19907 18199 19913
rect 18141 19904 18153 19907
rect 18104 19876 18153 19904
rect 18104 19864 18110 19876
rect 18141 19873 18153 19876
rect 18187 19873 18199 19907
rect 18141 19867 18199 19873
rect 8205 19799 8263 19805
rect 8312 19808 17448 19836
rect 2317 19771 2375 19777
rect 2317 19737 2329 19771
rect 2363 19737 2375 19771
rect 2317 19731 2375 19737
rect 2593 19771 2651 19777
rect 2593 19737 2605 19771
rect 2639 19768 2651 19771
rect 4062 19768 4068 19780
rect 2639 19740 4068 19768
rect 2639 19737 2651 19740
rect 2593 19731 2651 19737
rect 4062 19728 4068 19740
rect 4120 19728 4126 19780
rect 8312 19768 8340 19808
rect 6748 19740 8340 19768
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 2866 19700 2872 19712
rect 2827 19672 2872 19700
rect 2866 19660 2872 19672
rect 2924 19660 2930 19712
rect 3145 19703 3203 19709
rect 3145 19669 3157 19703
rect 3191 19700 3203 19703
rect 3234 19700 3240 19712
rect 3191 19672 3240 19700
rect 3191 19669 3203 19672
rect 3145 19663 3203 19669
rect 3234 19660 3240 19672
rect 3292 19660 3298 19712
rect 3418 19700 3424 19712
rect 3379 19672 3424 19700
rect 3418 19660 3424 19672
rect 3476 19660 3482 19712
rect 3697 19703 3755 19709
rect 3697 19669 3709 19703
rect 3743 19700 3755 19703
rect 3786 19700 3792 19712
rect 3743 19672 3792 19700
rect 3743 19669 3755 19672
rect 3697 19663 3755 19669
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 3973 19703 4031 19709
rect 3973 19669 3985 19703
rect 4019 19700 4031 19703
rect 4982 19700 4988 19712
rect 4019 19672 4988 19700
rect 4019 19669 4031 19672
rect 3973 19663 4031 19669
rect 4982 19660 4988 19672
rect 5040 19660 5046 19712
rect 6178 19660 6184 19712
rect 6236 19700 6242 19712
rect 6748 19700 6776 19740
rect 10134 19728 10140 19780
rect 10192 19768 10198 19780
rect 11057 19771 11115 19777
rect 11057 19768 11069 19771
rect 10192 19740 11069 19768
rect 10192 19728 10198 19740
rect 11057 19737 11069 19740
rect 11103 19737 11115 19771
rect 17494 19768 17500 19780
rect 17455 19740 17500 19768
rect 11057 19731 11115 19737
rect 17494 19728 17500 19740
rect 17552 19728 17558 19780
rect 18432 19777 18460 19944
rect 18616 19913 18644 20012
rect 19242 20000 19248 20052
rect 19300 20040 19306 20052
rect 19300 20012 20944 20040
rect 19300 20000 19306 20012
rect 19058 19932 19064 19984
rect 19116 19972 19122 19984
rect 20070 19972 20076 19984
rect 19116 19944 19932 19972
rect 20031 19944 20076 19972
rect 19116 19932 19122 19944
rect 19158 19913 19186 19944
rect 18601 19907 18659 19913
rect 18601 19873 18613 19907
rect 18647 19904 18659 19907
rect 19153 19907 19211 19913
rect 18647 19876 19104 19904
rect 18647 19873 18659 19876
rect 18601 19867 18659 19873
rect 19076 19848 19104 19876
rect 19153 19873 19165 19907
rect 19199 19873 19211 19907
rect 19153 19867 19211 19873
rect 19245 19907 19303 19913
rect 19245 19873 19257 19907
rect 19291 19904 19303 19907
rect 19426 19904 19432 19916
rect 19291 19876 19432 19904
rect 19291 19873 19303 19876
rect 19245 19867 19303 19873
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 19702 19904 19708 19916
rect 19663 19876 19708 19904
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 19904 19904 19932 19944
rect 20070 19932 20076 19944
rect 20128 19932 20134 19984
rect 20438 19932 20444 19984
rect 20496 19972 20502 19984
rect 20625 19975 20683 19981
rect 20496 19944 20541 19972
rect 20496 19932 20502 19944
rect 20625 19941 20637 19975
rect 20671 19972 20683 19975
rect 20714 19972 20720 19984
rect 20671 19944 20720 19972
rect 20671 19941 20683 19944
rect 20625 19935 20683 19941
rect 20714 19932 20720 19944
rect 20772 19932 20778 19984
rect 20916 19981 20944 20012
rect 20901 19975 20959 19981
rect 20901 19941 20913 19975
rect 20947 19941 20959 19975
rect 22002 19972 22008 19984
rect 20901 19935 20959 19941
rect 21284 19944 22008 19972
rect 20990 19904 20996 19916
rect 19904 19876 20996 19904
rect 20990 19864 20996 19876
rect 21048 19904 21054 19916
rect 21177 19907 21235 19913
rect 21177 19904 21189 19907
rect 21048 19876 21189 19904
rect 21048 19864 21054 19876
rect 21177 19873 21189 19876
rect 21223 19873 21235 19907
rect 21177 19867 21235 19873
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 18877 19839 18935 19845
rect 18877 19836 18889 19839
rect 18748 19808 18889 19836
rect 18748 19796 18754 19808
rect 18877 19805 18889 19808
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 19058 19796 19064 19848
rect 19116 19796 19122 19848
rect 19886 19836 19892 19848
rect 19847 19808 19892 19836
rect 19886 19796 19892 19808
rect 19944 19796 19950 19848
rect 20257 19839 20315 19845
rect 20257 19805 20269 19839
rect 20303 19836 20315 19839
rect 21284 19836 21312 19944
rect 22002 19932 22008 19944
rect 22060 19932 22066 19984
rect 21361 19907 21419 19913
rect 21361 19873 21373 19907
rect 21407 19873 21419 19907
rect 21361 19867 21419 19873
rect 20303 19808 21312 19836
rect 20303 19805 20315 19808
rect 20257 19799 20315 19805
rect 18417 19771 18475 19777
rect 18417 19737 18429 19771
rect 18463 19737 18475 19771
rect 18417 19731 18475 19737
rect 19429 19771 19487 19777
rect 19429 19737 19441 19771
rect 19475 19768 19487 19771
rect 20530 19768 20536 19780
rect 19475 19740 20536 19768
rect 19475 19737 19487 19740
rect 19429 19731 19487 19737
rect 20530 19728 20536 19740
rect 20588 19728 20594 19780
rect 21376 19768 21404 19867
rect 20732 19740 21404 19768
rect 6236 19672 6776 19700
rect 6236 19660 6242 19672
rect 6914 19660 6920 19712
rect 6972 19700 6978 19712
rect 7193 19703 7251 19709
rect 7193 19700 7205 19703
rect 6972 19672 7205 19700
rect 6972 19660 6978 19672
rect 7193 19669 7205 19672
rect 7239 19669 7251 19703
rect 7193 19663 7251 19669
rect 7282 19660 7288 19712
rect 7340 19700 7346 19712
rect 7469 19703 7527 19709
rect 7469 19700 7481 19703
rect 7340 19672 7481 19700
rect 7340 19660 7346 19672
rect 7469 19669 7481 19672
rect 7515 19669 7527 19703
rect 7650 19700 7656 19712
rect 7611 19672 7656 19700
rect 7469 19663 7527 19669
rect 7650 19660 7656 19672
rect 7708 19660 7714 19712
rect 7742 19660 7748 19712
rect 7800 19700 7806 19712
rect 8294 19700 8300 19712
rect 7800 19672 8300 19700
rect 7800 19660 7806 19672
rect 8294 19660 8300 19672
rect 8352 19660 8358 19712
rect 8481 19703 8539 19709
rect 8481 19669 8493 19703
rect 8527 19700 8539 19703
rect 9398 19700 9404 19712
rect 8527 19672 9404 19700
rect 8527 19669 8539 19672
rect 8481 19663 8539 19669
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 10226 19660 10232 19712
rect 10284 19700 10290 19712
rect 10597 19703 10655 19709
rect 10597 19700 10609 19703
rect 10284 19672 10609 19700
rect 10284 19660 10290 19672
rect 10597 19669 10609 19672
rect 10643 19669 10655 19703
rect 10597 19663 10655 19669
rect 10686 19660 10692 19712
rect 10744 19700 10750 19712
rect 10873 19703 10931 19709
rect 10873 19700 10885 19703
rect 10744 19672 10885 19700
rect 10744 19660 10750 19672
rect 10873 19669 10885 19672
rect 10919 19669 10931 19703
rect 11790 19700 11796 19712
rect 11751 19672 11796 19700
rect 10873 19663 10931 19669
rect 11790 19660 11796 19672
rect 11848 19660 11854 19712
rect 12345 19703 12403 19709
rect 12345 19669 12357 19703
rect 12391 19700 12403 19703
rect 13630 19700 13636 19712
rect 12391 19672 13636 19700
rect 12391 19669 12403 19672
rect 12345 19663 12403 19669
rect 13630 19660 13636 19672
rect 13688 19660 13694 19712
rect 17773 19703 17831 19709
rect 17773 19669 17785 19703
rect 17819 19700 17831 19703
rect 17862 19700 17868 19712
rect 17819 19672 17868 19700
rect 17819 19669 17831 19672
rect 17773 19663 17831 19669
rect 17862 19660 17868 19672
rect 17920 19660 17926 19712
rect 18049 19703 18107 19709
rect 18049 19669 18061 19703
rect 18095 19700 18107 19703
rect 18598 19700 18604 19712
rect 18095 19672 18604 19700
rect 18095 19669 18107 19672
rect 18049 19663 18107 19669
rect 18598 19660 18604 19672
rect 18656 19700 18662 19712
rect 19334 19700 19340 19712
rect 18656 19672 19340 19700
rect 18656 19660 18662 19672
rect 19334 19660 19340 19672
rect 19392 19660 19398 19712
rect 19794 19660 19800 19712
rect 19852 19700 19858 19712
rect 20732 19700 20760 19740
rect 21450 19700 21456 19712
rect 19852 19672 20760 19700
rect 21411 19672 21456 19700
rect 19852 19660 19858 19672
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 1578 19456 1584 19508
rect 1636 19496 1642 19508
rect 1765 19499 1823 19505
rect 1765 19496 1777 19499
rect 1636 19468 1777 19496
rect 1636 19456 1642 19468
rect 1765 19465 1777 19468
rect 1811 19465 1823 19499
rect 1765 19459 1823 19465
rect 2406 19456 2412 19508
rect 2464 19496 2470 19508
rect 3145 19499 3203 19505
rect 3145 19496 3157 19499
rect 2464 19468 3157 19496
rect 2464 19456 2470 19468
rect 3145 19465 3157 19468
rect 3191 19465 3203 19499
rect 3694 19496 3700 19508
rect 3655 19468 3700 19496
rect 3145 19459 3203 19465
rect 3694 19456 3700 19468
rect 3752 19456 3758 19508
rect 3970 19496 3976 19508
rect 3931 19468 3976 19496
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 6178 19496 6184 19508
rect 4632 19468 6184 19496
rect 2314 19388 2320 19440
rect 2372 19428 2378 19440
rect 4632 19428 4660 19468
rect 6178 19456 6184 19468
rect 6236 19456 6242 19508
rect 6270 19456 6276 19508
rect 6328 19496 6334 19508
rect 6825 19499 6883 19505
rect 6825 19496 6837 19499
rect 6328 19468 6837 19496
rect 6328 19456 6334 19468
rect 6825 19465 6837 19468
rect 6871 19465 6883 19499
rect 6825 19459 6883 19465
rect 7006 19456 7012 19508
rect 7064 19496 7070 19508
rect 10137 19499 10195 19505
rect 7064 19468 9260 19496
rect 7064 19456 7070 19468
rect 2372 19400 4660 19428
rect 2372 19388 2378 19400
rect 5994 19388 6000 19440
rect 6052 19428 6058 19440
rect 6457 19431 6515 19437
rect 6457 19428 6469 19431
rect 6052 19400 6469 19428
rect 6052 19388 6058 19400
rect 6457 19397 6469 19400
rect 6503 19397 6515 19431
rect 9232 19428 9260 19468
rect 10137 19465 10149 19499
rect 10183 19496 10195 19499
rect 10318 19496 10324 19508
rect 10183 19468 10324 19496
rect 10183 19465 10195 19468
rect 10137 19459 10195 19465
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 11238 19456 11244 19508
rect 11296 19496 11302 19508
rect 11425 19499 11483 19505
rect 11425 19496 11437 19499
rect 11296 19468 11437 19496
rect 11296 19456 11302 19468
rect 11425 19465 11437 19468
rect 11471 19465 11483 19499
rect 11425 19459 11483 19465
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 12529 19499 12587 19505
rect 12529 19496 12541 19499
rect 12492 19468 12541 19496
rect 12492 19456 12498 19468
rect 12529 19465 12541 19468
rect 12575 19465 12587 19499
rect 12529 19459 12587 19465
rect 12989 19499 13047 19505
rect 12989 19465 13001 19499
rect 13035 19496 13047 19499
rect 13170 19496 13176 19508
rect 13035 19468 13176 19496
rect 13035 19465 13047 19468
rect 12989 19459 13047 19465
rect 13170 19456 13176 19468
rect 13228 19456 13234 19508
rect 13265 19499 13323 19505
rect 13265 19465 13277 19499
rect 13311 19496 13323 19499
rect 13538 19496 13544 19508
rect 13311 19468 13544 19496
rect 13311 19465 13323 19468
rect 13265 19459 13323 19465
rect 13538 19456 13544 19468
rect 13596 19456 13602 19508
rect 13817 19499 13875 19505
rect 13817 19465 13829 19499
rect 13863 19496 13875 19499
rect 14274 19496 14280 19508
rect 13863 19468 14280 19496
rect 13863 19465 13875 19468
rect 13817 19459 13875 19465
rect 14274 19456 14280 19468
rect 14332 19456 14338 19508
rect 14553 19499 14611 19505
rect 14553 19465 14565 19499
rect 14599 19496 14611 19499
rect 14642 19496 14648 19508
rect 14599 19468 14648 19496
rect 14599 19465 14611 19468
rect 14553 19459 14611 19465
rect 14642 19456 14648 19468
rect 14700 19456 14706 19508
rect 15749 19499 15807 19505
rect 15749 19465 15761 19499
rect 15795 19496 15807 19499
rect 16482 19496 16488 19508
rect 15795 19468 16488 19496
rect 15795 19465 15807 19468
rect 15749 19459 15807 19465
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 16669 19499 16727 19505
rect 16669 19465 16681 19499
rect 16715 19496 16727 19499
rect 16850 19496 16856 19508
rect 16715 19468 16856 19496
rect 16715 19465 16727 19468
rect 16669 19459 16727 19465
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 17405 19499 17463 19505
rect 17405 19465 17417 19499
rect 17451 19496 17463 19499
rect 17770 19496 17776 19508
rect 17451 19468 17776 19496
rect 17451 19465 17463 19468
rect 17405 19459 17463 19465
rect 17770 19456 17776 19468
rect 17828 19456 17834 19508
rect 18049 19499 18107 19505
rect 18049 19465 18061 19499
rect 18095 19496 18107 19499
rect 19150 19496 19156 19508
rect 18095 19468 19156 19496
rect 18095 19465 18107 19468
rect 18049 19459 18107 19465
rect 19150 19456 19156 19468
rect 19208 19456 19214 19508
rect 21358 19496 21364 19508
rect 21319 19468 21364 19496
rect 21358 19456 21364 19468
rect 21416 19456 21422 19508
rect 12066 19428 12072 19440
rect 9232 19400 12072 19428
rect 6457 19391 6515 19397
rect 12066 19388 12072 19400
rect 12124 19388 12130 19440
rect 15289 19431 15347 19437
rect 15289 19397 15301 19431
rect 15335 19428 15347 19431
rect 16022 19428 16028 19440
rect 15335 19400 16028 19428
rect 15335 19397 15347 19400
rect 15289 19391 15347 19397
rect 16022 19388 16028 19400
rect 16080 19388 16086 19440
rect 17310 19388 17316 19440
rect 17368 19428 17374 19440
rect 18233 19431 18291 19437
rect 17368 19400 18184 19428
rect 17368 19388 17374 19400
rect 1780 19332 2084 19360
rect 1394 19292 1400 19304
rect 1355 19264 1400 19292
rect 1394 19252 1400 19264
rect 1452 19252 1458 19304
rect 1780 19292 1808 19332
rect 1946 19292 1952 19304
rect 1504 19264 1808 19292
rect 1907 19264 1952 19292
rect 1302 19184 1308 19236
rect 1360 19224 1366 19236
rect 1504 19224 1532 19264
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2056 19301 2084 19332
rect 2682 19320 2688 19372
rect 2740 19360 2746 19372
rect 2740 19332 3004 19360
rect 2740 19320 2746 19332
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19261 2099 19295
rect 2317 19295 2375 19301
rect 2317 19292 2329 19295
rect 2041 19255 2099 19261
rect 2148 19264 2329 19292
rect 1360 19196 1532 19224
rect 1581 19227 1639 19233
rect 1360 19184 1366 19196
rect 1581 19193 1593 19227
rect 1627 19224 1639 19227
rect 1854 19224 1860 19236
rect 1627 19196 1860 19224
rect 1627 19193 1639 19196
rect 1581 19187 1639 19193
rect 1854 19184 1860 19196
rect 1912 19184 1918 19236
rect 1670 19116 1676 19168
rect 1728 19156 1734 19168
rect 2148 19156 2176 19264
rect 2317 19261 2329 19264
rect 2363 19292 2375 19295
rect 2498 19292 2504 19304
rect 2363 19264 2504 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 2498 19252 2504 19264
rect 2556 19252 2562 19304
rect 2774 19292 2780 19304
rect 2735 19264 2780 19292
rect 2774 19252 2780 19264
rect 2832 19252 2838 19304
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19261 2927 19295
rect 2976 19292 3004 19332
rect 5626 19320 5632 19372
rect 5684 19360 5690 19372
rect 6546 19360 6552 19372
rect 5684 19332 6552 19360
rect 5684 19320 5690 19332
rect 6546 19320 6552 19332
rect 6604 19320 6610 19372
rect 9033 19363 9091 19369
rect 9033 19360 9045 19363
rect 8312 19332 9045 19360
rect 3329 19295 3387 19301
rect 3329 19292 3341 19295
rect 2976 19264 3341 19292
rect 2869 19255 2927 19261
rect 3329 19261 3341 19264
rect 3375 19261 3387 19295
rect 3329 19255 3387 19261
rect 3789 19295 3847 19301
rect 3789 19261 3801 19295
rect 3835 19292 3847 19295
rect 4890 19292 4896 19304
rect 3835 19264 4896 19292
rect 3835 19261 3847 19264
rect 3789 19255 3847 19261
rect 2682 19224 2688 19236
rect 2516 19196 2688 19224
rect 1728 19128 2176 19156
rect 2225 19159 2283 19165
rect 1728 19116 1734 19128
rect 2225 19125 2237 19159
rect 2271 19156 2283 19159
rect 2406 19156 2412 19168
rect 2271 19128 2412 19156
rect 2271 19125 2283 19128
rect 2225 19119 2283 19125
rect 2406 19116 2412 19128
rect 2464 19116 2470 19168
rect 2516 19165 2544 19196
rect 2682 19184 2688 19196
rect 2740 19184 2746 19236
rect 2884 19224 2912 19255
rect 4890 19252 4896 19264
rect 4948 19252 4954 19304
rect 4982 19252 4988 19304
rect 5040 19292 5046 19304
rect 5270 19295 5328 19301
rect 5270 19292 5282 19295
rect 5040 19264 5282 19292
rect 5040 19252 5046 19264
rect 5270 19261 5282 19264
rect 5316 19292 5328 19295
rect 5442 19292 5448 19304
rect 5316 19264 5448 19292
rect 5316 19261 5328 19264
rect 5270 19255 5328 19261
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 5537 19295 5595 19301
rect 5537 19261 5549 19295
rect 5583 19292 5595 19295
rect 5718 19292 5724 19304
rect 5583 19264 5724 19292
rect 5583 19261 5595 19264
rect 5537 19255 5595 19261
rect 5718 19252 5724 19264
rect 5776 19252 5782 19304
rect 5902 19292 5908 19304
rect 5863 19264 5908 19292
rect 5902 19252 5908 19264
rect 5960 19292 5966 19304
rect 6641 19295 6699 19301
rect 6641 19292 6653 19295
rect 5960 19264 6653 19292
rect 5960 19252 5966 19264
rect 6641 19261 6653 19264
rect 6687 19261 6699 19295
rect 8312 19292 8340 19332
rect 9033 19329 9045 19332
rect 9079 19329 9091 19363
rect 9033 19323 9091 19329
rect 10594 19320 10600 19372
rect 10652 19360 10658 19372
rect 10965 19363 11023 19369
rect 10965 19360 10977 19363
rect 10652 19332 10977 19360
rect 10652 19320 10658 19332
rect 10965 19329 10977 19332
rect 11011 19329 11023 19363
rect 11882 19360 11888 19372
rect 11843 19332 11888 19360
rect 10965 19323 11023 19329
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 14660 19332 14964 19360
rect 6641 19255 6699 19261
rect 8240 19264 8340 19292
rect 8389 19295 8447 19301
rect 3142 19224 3148 19236
rect 2884 19196 3148 19224
rect 3142 19184 3148 19196
rect 3200 19184 3206 19236
rect 4614 19184 4620 19236
rect 4672 19224 4678 19236
rect 5629 19227 5687 19233
rect 5629 19224 5641 19227
rect 4672 19196 5641 19224
rect 4672 19184 4678 19196
rect 5629 19193 5641 19196
rect 5675 19193 5687 19227
rect 6181 19227 6239 19233
rect 6181 19224 6193 19227
rect 5629 19187 5687 19193
rect 5736 19196 6193 19224
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19125 2559 19159
rect 2501 19119 2559 19125
rect 2593 19159 2651 19165
rect 2593 19125 2605 19159
rect 2639 19156 2651 19159
rect 2958 19156 2964 19168
rect 2639 19128 2964 19156
rect 2639 19125 2651 19128
rect 2593 19119 2651 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 3053 19159 3111 19165
rect 3053 19125 3065 19159
rect 3099 19156 3111 19159
rect 3786 19156 3792 19168
rect 3099 19128 3792 19156
rect 3099 19125 3111 19128
rect 3053 19119 3111 19125
rect 3786 19116 3792 19128
rect 3844 19116 3850 19168
rect 4154 19156 4160 19168
rect 4115 19128 4160 19156
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 5166 19116 5172 19168
rect 5224 19156 5230 19168
rect 5736 19156 5764 19196
rect 6181 19193 6193 19196
rect 6227 19193 6239 19227
rect 6181 19187 6239 19193
rect 7466 19184 7472 19236
rect 7524 19224 7530 19236
rect 8110 19224 8116 19236
rect 8168 19233 8174 19236
rect 7524 19196 8116 19224
rect 7524 19184 7530 19196
rect 8110 19184 8116 19196
rect 8168 19224 8180 19233
rect 8240 19224 8268 19264
rect 8389 19261 8401 19295
rect 8435 19292 8447 19295
rect 9306 19292 9312 19304
rect 8435 19264 9076 19292
rect 9267 19264 9312 19292
rect 8435 19261 8447 19264
rect 8389 19255 8447 19261
rect 9048 19236 9076 19264
rect 9306 19252 9312 19264
rect 9364 19252 9370 19304
rect 9677 19295 9735 19301
rect 9677 19292 9689 19295
rect 9508 19264 9689 19292
rect 8168 19196 8268 19224
rect 8168 19187 8180 19196
rect 8168 19184 8174 19187
rect 8846 19184 8852 19236
rect 8904 19224 8910 19236
rect 8904 19196 8949 19224
rect 8904 19184 8910 19196
rect 9030 19184 9036 19236
rect 9088 19184 9094 19236
rect 5224 19128 5764 19156
rect 5224 19116 5230 19128
rect 5994 19116 6000 19168
rect 6052 19156 6058 19168
rect 6089 19159 6147 19165
rect 6089 19156 6101 19159
rect 6052 19128 6101 19156
rect 6052 19116 6058 19128
rect 6089 19125 6101 19128
rect 6135 19125 6147 19159
rect 6089 19119 6147 19125
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 7009 19159 7067 19165
rect 7009 19156 7021 19159
rect 6880 19128 7021 19156
rect 6880 19116 6886 19128
rect 7009 19125 7021 19128
rect 7055 19125 7067 19159
rect 7009 19119 7067 19125
rect 7558 19116 7564 19168
rect 7616 19156 7622 19168
rect 8481 19159 8539 19165
rect 8481 19156 8493 19159
rect 7616 19128 8493 19156
rect 7616 19116 7622 19128
rect 8481 19125 8493 19128
rect 8527 19125 8539 19159
rect 8938 19156 8944 19168
rect 8899 19128 8944 19156
rect 8481 19119 8539 19125
rect 8938 19116 8944 19128
rect 8996 19116 9002 19168
rect 9508 19165 9536 19264
rect 9677 19261 9689 19264
rect 9723 19261 9735 19295
rect 9677 19255 9735 19261
rect 9858 19252 9864 19304
rect 9916 19292 9922 19304
rect 9953 19295 10011 19301
rect 9953 19292 9965 19295
rect 9916 19264 9965 19292
rect 9916 19252 9922 19264
rect 9953 19261 9965 19264
rect 9999 19261 10011 19295
rect 11054 19292 11060 19304
rect 9953 19255 10011 19261
rect 10428 19264 11060 19292
rect 10428 19224 10456 19264
rect 11054 19252 11060 19264
rect 11112 19252 11118 19304
rect 11238 19292 11244 19304
rect 11199 19264 11244 19292
rect 11238 19252 11244 19264
rect 11296 19252 11302 19304
rect 12250 19252 12256 19304
rect 12308 19292 12314 19304
rect 12713 19295 12771 19301
rect 12713 19292 12725 19295
rect 12308 19264 12725 19292
rect 12308 19252 12314 19264
rect 12713 19261 12725 19264
rect 12759 19261 12771 19295
rect 12713 19255 12771 19261
rect 12802 19252 12808 19304
rect 12860 19292 12866 19304
rect 13081 19295 13139 19301
rect 12860 19264 12905 19292
rect 12860 19252 12866 19264
rect 13081 19261 13093 19295
rect 13127 19261 13139 19295
rect 13081 19255 13139 19261
rect 13357 19295 13415 19301
rect 13357 19261 13369 19295
rect 13403 19261 13415 19295
rect 13630 19292 13636 19304
rect 13591 19264 13636 19292
rect 13357 19255 13415 19261
rect 9876 19196 10456 19224
rect 10781 19227 10839 19233
rect 9876 19165 9904 19196
rect 10781 19193 10793 19227
rect 10827 19224 10839 19227
rect 11790 19224 11796 19236
rect 10827 19196 11796 19224
rect 10827 19193 10839 19196
rect 10781 19187 10839 19193
rect 11790 19184 11796 19196
rect 11848 19184 11854 19236
rect 12894 19184 12900 19236
rect 12952 19224 12958 19236
rect 13096 19224 13124 19255
rect 12952 19196 13124 19224
rect 13372 19224 13400 19255
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 13998 19252 14004 19304
rect 14056 19292 14062 19304
rect 14277 19295 14335 19301
rect 14277 19292 14289 19295
rect 14056 19264 14289 19292
rect 14056 19252 14062 19264
rect 14277 19261 14289 19264
rect 14323 19292 14335 19295
rect 14369 19295 14427 19301
rect 14369 19292 14381 19295
rect 14323 19264 14381 19292
rect 14323 19261 14335 19264
rect 14277 19255 14335 19261
rect 14369 19261 14381 19264
rect 14415 19261 14427 19295
rect 14369 19255 14427 19261
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 14660 19292 14688 19332
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 14516 19264 14688 19292
rect 14752 19264 14841 19292
rect 14516 19252 14522 19264
rect 13372 19196 14044 19224
rect 12952 19184 12958 19196
rect 9493 19159 9551 19165
rect 9493 19125 9505 19159
rect 9539 19125 9551 19159
rect 9493 19119 9551 19125
rect 9861 19159 9919 19165
rect 9861 19125 9873 19159
rect 9907 19125 9919 19159
rect 10410 19156 10416 19168
rect 10371 19128 10416 19156
rect 9861 19119 9919 19125
rect 10410 19116 10416 19128
rect 10468 19116 10474 19168
rect 10870 19116 10876 19168
rect 10928 19156 10934 19168
rect 10928 19128 10973 19156
rect 10928 19116 10934 19128
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 11977 19159 12035 19165
rect 11977 19156 11989 19159
rect 11112 19128 11989 19156
rect 11112 19116 11118 19128
rect 11977 19125 11989 19128
rect 12023 19125 12035 19159
rect 11977 19119 12035 19125
rect 12066 19116 12072 19168
rect 12124 19156 12130 19168
rect 12437 19159 12495 19165
rect 12124 19128 12169 19156
rect 12124 19116 12130 19128
rect 12437 19125 12449 19159
rect 12483 19156 12495 19159
rect 12526 19156 12532 19168
rect 12483 19128 12532 19156
rect 12483 19125 12495 19128
rect 12437 19119 12495 19125
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 13541 19159 13599 19165
rect 13541 19125 13553 19159
rect 13587 19156 13599 19159
rect 13722 19156 13728 19168
rect 13587 19128 13728 19156
rect 13587 19125 13599 19128
rect 13541 19119 13599 19125
rect 13722 19116 13728 19128
rect 13780 19116 13786 19168
rect 14016 19165 14044 19196
rect 14752 19168 14780 19264
rect 14829 19261 14841 19264
rect 14875 19261 14887 19295
rect 14936 19292 14964 19332
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 18156 19360 18184 19400
rect 18233 19397 18245 19431
rect 18279 19428 18291 19431
rect 18966 19428 18972 19440
rect 18279 19400 18972 19428
rect 18279 19397 18291 19400
rect 18233 19391 18291 19397
rect 18966 19388 18972 19400
rect 19024 19388 19030 19440
rect 19058 19388 19064 19440
rect 19116 19428 19122 19440
rect 20530 19428 20536 19440
rect 19116 19400 20536 19428
rect 19116 19388 19122 19400
rect 20530 19388 20536 19400
rect 20588 19428 20594 19440
rect 20588 19400 21588 19428
rect 20588 19388 20594 19400
rect 20993 19363 21051 19369
rect 20993 19360 21005 19363
rect 17828 19332 18092 19360
rect 18156 19332 21005 19360
rect 17828 19320 17834 19332
rect 15105 19295 15163 19301
rect 15105 19292 15117 19295
rect 14936 19264 15117 19292
rect 14829 19255 14887 19261
rect 15105 19261 15117 19264
rect 15151 19292 15163 19295
rect 15381 19295 15439 19301
rect 15381 19292 15393 19295
rect 15151 19264 15393 19292
rect 15151 19261 15163 19264
rect 15105 19255 15163 19261
rect 15381 19261 15393 19264
rect 15427 19261 15439 19295
rect 15381 19255 15439 19261
rect 15470 19252 15476 19304
rect 15528 19292 15534 19304
rect 15565 19295 15623 19301
rect 15565 19292 15577 19295
rect 15528 19264 15577 19292
rect 15528 19252 15534 19264
rect 15565 19261 15577 19264
rect 15611 19261 15623 19295
rect 16114 19292 16120 19304
rect 16075 19264 16120 19292
rect 15565 19255 15623 19261
rect 15580 19224 15608 19255
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 16485 19295 16543 19301
rect 16485 19261 16497 19295
rect 16531 19292 16543 19295
rect 17218 19292 17224 19304
rect 16531 19264 17080 19292
rect 17179 19264 17224 19292
rect 16531 19261 16543 19264
rect 16485 19255 16543 19261
rect 16209 19227 16267 19233
rect 16209 19224 16221 19227
rect 15580 19196 16221 19224
rect 16209 19193 16221 19196
rect 16255 19193 16267 19227
rect 16209 19187 16267 19193
rect 17052 19168 17080 19264
rect 17218 19252 17224 19264
rect 17276 19252 17282 19304
rect 17494 19252 17500 19304
rect 17552 19292 17558 19304
rect 17589 19295 17647 19301
rect 17589 19292 17601 19295
rect 17552 19264 17601 19292
rect 17552 19252 17558 19264
rect 17589 19261 17601 19264
rect 17635 19261 17647 19295
rect 17589 19255 17647 19261
rect 17865 19295 17923 19301
rect 17865 19261 17877 19295
rect 17911 19261 17923 19295
rect 18064 19292 18092 19332
rect 20993 19329 21005 19332
rect 21039 19329 21051 19363
rect 20993 19323 21051 19329
rect 18509 19295 18567 19301
rect 18509 19292 18521 19295
rect 18064 19264 18521 19292
rect 17865 19255 17923 19261
rect 18509 19261 18521 19264
rect 18555 19261 18567 19295
rect 18509 19255 18567 19261
rect 17880 19224 17908 19255
rect 17604 19196 17908 19224
rect 17604 19168 17632 19196
rect 18046 19184 18052 19236
rect 18104 19224 18110 19236
rect 18325 19227 18383 19233
rect 18325 19224 18337 19227
rect 18104 19196 18337 19224
rect 18104 19184 18110 19196
rect 18325 19193 18337 19196
rect 18371 19193 18383 19227
rect 18524 19224 18552 19255
rect 18782 19252 18788 19304
rect 18840 19292 18846 19304
rect 18877 19295 18935 19301
rect 18877 19292 18889 19295
rect 18840 19264 18889 19292
rect 18840 19252 18846 19264
rect 18877 19261 18889 19264
rect 18923 19261 18935 19295
rect 18877 19255 18935 19261
rect 19150 19252 19156 19304
rect 19208 19292 19214 19304
rect 20714 19292 20720 19304
rect 19208 19264 20720 19292
rect 19208 19252 19214 19264
rect 20714 19252 20720 19264
rect 20772 19252 20778 19304
rect 20809 19295 20867 19301
rect 20809 19261 20821 19295
rect 20855 19292 20867 19295
rect 20898 19292 20904 19304
rect 20855 19264 20904 19292
rect 20855 19261 20867 19264
rect 20809 19255 20867 19261
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 21560 19301 21588 19400
rect 21545 19295 21603 19301
rect 21545 19261 21557 19295
rect 21591 19261 21603 19295
rect 21545 19255 21603 19261
rect 18969 19227 19027 19233
rect 18524 19196 18920 19224
rect 18325 19187 18383 19193
rect 14001 19159 14059 19165
rect 14001 19125 14013 19159
rect 14047 19156 14059 19159
rect 14458 19156 14464 19168
rect 14047 19128 14464 19156
rect 14047 19125 14059 19128
rect 14001 19119 14059 19125
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 14734 19156 14740 19168
rect 14695 19128 14740 19156
rect 14734 19116 14740 19128
rect 14792 19116 14798 19168
rect 15013 19159 15071 19165
rect 15013 19125 15025 19159
rect 15059 19156 15071 19159
rect 15194 19156 15200 19168
rect 15059 19128 15200 19156
rect 15059 19125 15071 19128
rect 15013 19119 15071 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 15930 19156 15936 19168
rect 15891 19128 15936 19156
rect 15930 19116 15936 19128
rect 15988 19116 15994 19168
rect 17034 19156 17040 19168
rect 16995 19128 17040 19156
rect 17034 19116 17040 19128
rect 17092 19116 17098 19168
rect 17586 19116 17592 19168
rect 17644 19116 17650 19168
rect 17773 19159 17831 19165
rect 17773 19125 17785 19159
rect 17819 19156 17831 19159
rect 17954 19156 17960 19168
rect 17819 19128 17960 19156
rect 17819 19125 17831 19128
rect 17773 19119 17831 19125
rect 17954 19116 17960 19128
rect 18012 19116 18018 19168
rect 18690 19156 18696 19168
rect 18651 19128 18696 19156
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 18892 19156 18920 19196
rect 18969 19193 18981 19227
rect 19015 19224 19027 19227
rect 19242 19224 19248 19236
rect 19015 19196 19248 19224
rect 19015 19193 19027 19196
rect 18969 19187 19027 19193
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 19886 19156 19892 19168
rect 18892 19128 19892 19156
rect 19886 19116 19892 19128
rect 19944 19116 19950 19168
rect 20070 19116 20076 19168
rect 20128 19156 20134 19168
rect 20257 19159 20315 19165
rect 20257 19156 20269 19159
rect 20128 19128 20269 19156
rect 20128 19116 20134 19128
rect 20257 19125 20269 19128
rect 20303 19125 20315 19159
rect 20257 19119 20315 19125
rect 20714 19116 20720 19168
rect 20772 19156 20778 19168
rect 21082 19156 21088 19168
rect 20772 19128 21088 19156
rect 20772 19116 20778 19128
rect 21082 19116 21088 19128
rect 21140 19116 21146 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1765 18955 1823 18961
rect 1765 18952 1777 18955
rect 1596 18924 1777 18952
rect 1394 18884 1400 18896
rect 1355 18856 1400 18884
rect 1394 18844 1400 18856
rect 1452 18844 1458 18896
rect 1596 18893 1624 18924
rect 1765 18921 1777 18924
rect 1811 18921 1823 18955
rect 1765 18915 1823 18921
rect 1854 18912 1860 18964
rect 1912 18952 1918 18964
rect 2041 18955 2099 18961
rect 2041 18952 2053 18955
rect 1912 18924 2053 18952
rect 1912 18912 1918 18924
rect 2041 18921 2053 18924
rect 2087 18921 2099 18955
rect 2041 18915 2099 18921
rect 2222 18912 2228 18964
rect 2280 18952 2286 18964
rect 2317 18955 2375 18961
rect 2317 18952 2329 18955
rect 2280 18924 2329 18952
rect 2280 18912 2286 18924
rect 2317 18921 2329 18924
rect 2363 18921 2375 18955
rect 2317 18915 2375 18921
rect 2498 18912 2504 18964
rect 2556 18952 2562 18964
rect 2961 18955 3019 18961
rect 2961 18952 2973 18955
rect 2556 18924 2973 18952
rect 2556 18912 2562 18924
rect 2961 18921 2973 18924
rect 3007 18921 3019 18955
rect 2961 18915 3019 18921
rect 3142 18912 3148 18964
rect 3200 18952 3206 18964
rect 3513 18955 3571 18961
rect 3513 18952 3525 18955
rect 3200 18924 3525 18952
rect 3200 18912 3206 18924
rect 3513 18921 3525 18924
rect 3559 18921 3571 18955
rect 3513 18915 3571 18921
rect 4062 18912 4068 18964
rect 4120 18952 4126 18964
rect 4801 18955 4859 18961
rect 4801 18952 4813 18955
rect 4120 18924 4813 18952
rect 4120 18912 4126 18924
rect 4801 18921 4813 18924
rect 4847 18921 4859 18955
rect 4801 18915 4859 18921
rect 5258 18912 5264 18964
rect 5316 18952 5322 18964
rect 5353 18955 5411 18961
rect 5353 18952 5365 18955
rect 5316 18924 5365 18952
rect 5316 18912 5322 18924
rect 5353 18921 5365 18924
rect 5399 18921 5411 18955
rect 5353 18915 5411 18921
rect 6454 18912 6460 18964
rect 6512 18952 6518 18964
rect 6914 18952 6920 18964
rect 6512 18924 6920 18952
rect 6512 18912 6518 18924
rect 6914 18912 6920 18924
rect 6972 18912 6978 18964
rect 7098 18952 7104 18964
rect 7059 18924 7104 18952
rect 7098 18912 7104 18924
rect 7156 18912 7162 18964
rect 7650 18952 7656 18964
rect 7611 18924 7656 18952
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 8021 18955 8079 18961
rect 8021 18921 8033 18955
rect 8067 18952 8079 18955
rect 8573 18955 8631 18961
rect 8573 18952 8585 18955
rect 8067 18924 8585 18952
rect 8067 18921 8079 18924
rect 8021 18915 8079 18921
rect 8573 18921 8585 18924
rect 8619 18921 8631 18955
rect 8573 18915 8631 18921
rect 10137 18955 10195 18961
rect 10137 18921 10149 18955
rect 10183 18952 10195 18955
rect 10410 18952 10416 18964
rect 10183 18924 10416 18952
rect 10183 18921 10195 18924
rect 10137 18915 10195 18921
rect 10410 18912 10416 18924
rect 10468 18912 10474 18964
rect 10505 18955 10563 18961
rect 10505 18921 10517 18955
rect 10551 18952 10563 18955
rect 11054 18952 11060 18964
rect 10551 18924 11060 18952
rect 10551 18921 10563 18924
rect 10505 18915 10563 18921
rect 11054 18912 11060 18924
rect 11112 18912 11118 18964
rect 11882 18912 11888 18964
rect 11940 18952 11946 18964
rect 11977 18955 12035 18961
rect 11977 18952 11989 18955
rect 11940 18924 11989 18952
rect 11940 18912 11946 18924
rect 11977 18921 11989 18924
rect 12023 18921 12035 18955
rect 11977 18915 12035 18921
rect 12713 18955 12771 18961
rect 12713 18921 12725 18955
rect 12759 18952 12771 18955
rect 12802 18952 12808 18964
rect 12759 18924 12808 18952
rect 12759 18921 12771 18924
rect 12713 18915 12771 18921
rect 12802 18912 12808 18924
rect 12860 18912 12866 18964
rect 14369 18955 14427 18961
rect 14369 18921 14381 18955
rect 14415 18952 14427 18955
rect 14550 18952 14556 18964
rect 14415 18924 14556 18952
rect 14415 18921 14427 18924
rect 14369 18915 14427 18921
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 18138 18952 18144 18964
rect 18099 18924 18144 18952
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 18414 18952 18420 18964
rect 18375 18924 18420 18952
rect 18414 18912 18420 18924
rect 18472 18912 18478 18964
rect 19242 18952 19248 18964
rect 19203 18924 19248 18952
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 19702 18952 19708 18964
rect 19663 18924 19708 18952
rect 19702 18912 19708 18924
rect 19760 18912 19766 18964
rect 19978 18912 19984 18964
rect 20036 18912 20042 18964
rect 20165 18955 20223 18961
rect 20165 18921 20177 18955
rect 20211 18952 20223 18955
rect 20438 18952 20444 18964
rect 20211 18924 20444 18952
rect 20211 18921 20223 18924
rect 20165 18915 20223 18921
rect 20438 18912 20444 18924
rect 20496 18912 20502 18964
rect 20717 18955 20775 18961
rect 20717 18921 20729 18955
rect 20763 18952 20775 18955
rect 22738 18952 22744 18964
rect 20763 18924 22744 18952
rect 20763 18921 20775 18924
rect 20717 18915 20775 18921
rect 22738 18912 22744 18924
rect 22796 18912 22802 18964
rect 1581 18887 1639 18893
rect 1581 18853 1593 18887
rect 1627 18853 1639 18887
rect 2593 18887 2651 18893
rect 2593 18884 2605 18887
rect 1581 18847 1639 18853
rect 1780 18856 2605 18884
rect 1780 18828 1808 18856
rect 2593 18853 2605 18856
rect 2639 18853 2651 18887
rect 3326 18884 3332 18896
rect 3287 18856 3332 18884
rect 2593 18847 2651 18853
rect 3326 18844 3332 18856
rect 3384 18844 3390 18896
rect 3878 18844 3884 18896
rect 3936 18884 3942 18896
rect 4893 18887 4951 18893
rect 4893 18884 4905 18887
rect 3936 18856 4905 18884
rect 3936 18844 3942 18856
rect 4893 18853 4905 18856
rect 4939 18884 4951 18887
rect 5626 18884 5632 18896
rect 4939 18856 5632 18884
rect 4939 18853 4951 18856
rect 4893 18847 4951 18853
rect 5626 18844 5632 18856
rect 5684 18844 5690 18896
rect 10962 18884 10968 18896
rect 5736 18856 10968 18884
rect 1762 18776 1768 18828
rect 1820 18776 1826 18828
rect 1946 18816 1952 18828
rect 1907 18788 1952 18816
rect 1946 18776 1952 18788
rect 2004 18776 2010 18828
rect 2225 18819 2283 18825
rect 2225 18785 2237 18819
rect 2271 18785 2283 18819
rect 2498 18816 2504 18828
rect 2459 18788 2504 18816
rect 2225 18779 2283 18785
rect 2240 18748 2268 18779
rect 2498 18776 2504 18788
rect 2556 18776 2562 18828
rect 3050 18776 3056 18828
rect 3108 18816 3114 18828
rect 3145 18819 3203 18825
rect 3145 18816 3157 18819
rect 3108 18788 3157 18816
rect 3108 18776 3114 18788
rect 3145 18785 3157 18788
rect 3191 18785 3203 18819
rect 3145 18779 3203 18785
rect 3970 18776 3976 18828
rect 4028 18816 4034 18828
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 4028 18788 4353 18816
rect 4028 18776 4034 18788
rect 4341 18785 4353 18788
rect 4387 18785 4399 18819
rect 5442 18816 5448 18828
rect 4341 18779 4399 18785
rect 5092 18788 5448 18816
rect 3510 18748 3516 18760
rect 2240 18720 3516 18748
rect 3510 18708 3516 18720
rect 3568 18748 3574 18760
rect 3697 18751 3755 18757
rect 3568 18720 3648 18748
rect 3568 18708 3574 18720
rect 2777 18683 2835 18689
rect 2777 18680 2789 18683
rect 2608 18652 2789 18680
rect 1302 18572 1308 18624
rect 1360 18612 1366 18624
rect 2608 18612 2636 18652
rect 2777 18649 2789 18652
rect 2823 18649 2835 18683
rect 3620 18680 3648 18720
rect 3697 18717 3709 18751
rect 3743 18748 3755 18751
rect 4246 18748 4252 18760
rect 3743 18720 4252 18748
rect 3743 18717 3755 18720
rect 3697 18711 3755 18717
rect 4246 18708 4252 18720
rect 4304 18708 4310 18760
rect 5092 18757 5120 18788
rect 5442 18776 5448 18788
rect 5500 18776 5506 18828
rect 5077 18751 5135 18757
rect 5077 18717 5089 18751
rect 5123 18717 5135 18751
rect 5077 18711 5135 18717
rect 3973 18683 4031 18689
rect 3973 18680 3985 18683
rect 3620 18652 3985 18680
rect 2777 18643 2835 18649
rect 3973 18649 3985 18652
rect 4019 18649 4031 18683
rect 3973 18643 4031 18649
rect 4430 18640 4436 18692
rect 4488 18680 4494 18692
rect 5736 18680 5764 18856
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 11992 18856 14044 18884
rect 11992 18828 12020 18856
rect 6178 18776 6184 18828
rect 6236 18816 6242 18828
rect 6454 18816 6460 18828
rect 6512 18825 6518 18828
rect 6236 18788 6460 18816
rect 6236 18776 6242 18788
rect 6454 18776 6460 18788
rect 6512 18779 6524 18825
rect 6512 18776 6518 18779
rect 6638 18776 6644 18828
rect 6696 18816 6702 18828
rect 6696 18788 7420 18816
rect 6696 18776 6702 18788
rect 7392 18757 7420 18788
rect 8202 18776 8208 18828
rect 8260 18816 8266 18828
rect 8481 18819 8539 18825
rect 8481 18816 8493 18819
rect 8260 18788 8493 18816
rect 8260 18776 8266 18788
rect 8481 18785 8493 18788
rect 8527 18785 8539 18819
rect 10864 18819 10922 18825
rect 10864 18816 10876 18819
rect 8481 18779 8539 18785
rect 9876 18788 10876 18816
rect 6733 18751 6791 18757
rect 6733 18717 6745 18751
rect 6779 18717 6791 18751
rect 6733 18711 6791 18717
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 7377 18751 7435 18757
rect 7377 18717 7389 18751
rect 7423 18717 7435 18751
rect 7558 18748 7564 18760
rect 7519 18720 7564 18748
rect 7377 18711 7435 18717
rect 4488 18652 4533 18680
rect 5368 18652 5764 18680
rect 4488 18640 4494 18652
rect 1360 18584 2636 18612
rect 1360 18572 1366 18584
rect 2682 18572 2688 18624
rect 2740 18612 2746 18624
rect 3697 18615 3755 18621
rect 3697 18612 3709 18615
rect 2740 18584 3709 18612
rect 2740 18572 2746 18584
rect 3697 18581 3709 18584
rect 3743 18581 3755 18615
rect 3697 18575 3755 18581
rect 3878 18572 3884 18624
rect 3936 18612 3942 18624
rect 4157 18615 4215 18621
rect 4157 18612 4169 18615
rect 3936 18584 4169 18612
rect 3936 18572 3942 18584
rect 4157 18581 4169 18584
rect 4203 18612 4215 18615
rect 5368 18612 5396 18652
rect 4203 18584 5396 18612
rect 4203 18581 4215 18584
rect 4157 18575 4215 18581
rect 5718 18572 5724 18624
rect 5776 18612 5782 18624
rect 6748 18612 6776 18711
rect 6840 18624 6868 18711
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 9876 18757 9904 18788
rect 10864 18785 10876 18788
rect 10910 18816 10922 18819
rect 11146 18816 11152 18828
rect 10910 18788 11152 18816
rect 10910 18785 10922 18788
rect 10864 18779 10922 18785
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 11974 18776 11980 18828
rect 12032 18776 12038 18828
rect 12250 18776 12256 18828
rect 12308 18816 12314 18828
rect 12345 18819 12403 18825
rect 12345 18816 12357 18819
rect 12308 18788 12357 18816
rect 12308 18776 12314 18788
rect 12345 18785 12357 18788
rect 12391 18785 12403 18819
rect 14016 18816 14044 18856
rect 18598 18844 18604 18896
rect 18656 18884 18662 18896
rect 19610 18884 19616 18896
rect 18656 18856 18920 18884
rect 18656 18844 18662 18856
rect 14553 18819 14611 18825
rect 14553 18816 14565 18819
rect 14016 18788 14565 18816
rect 12345 18779 12403 18785
rect 14553 18785 14565 18788
rect 14599 18816 14611 18819
rect 14645 18819 14703 18825
rect 14645 18816 14657 18819
rect 14599 18788 14657 18816
rect 14599 18785 14611 18788
rect 14553 18779 14611 18785
rect 14645 18785 14657 18788
rect 14691 18785 14703 18819
rect 14645 18779 14703 18785
rect 16114 18776 16120 18828
rect 16172 18816 16178 18828
rect 18892 18825 18920 18856
rect 19444 18856 19616 18884
rect 19444 18825 19472 18856
rect 19610 18844 19616 18856
rect 19668 18884 19674 18896
rect 19996 18884 20024 18912
rect 20530 18884 20536 18896
rect 19668 18856 20024 18884
rect 20456 18856 20536 18884
rect 19668 18844 19674 18856
rect 18877 18819 18935 18825
rect 16172 18788 18736 18816
rect 16172 18776 16178 18788
rect 8665 18751 8723 18757
rect 8665 18717 8677 18751
rect 8711 18717 8723 18751
rect 8665 18711 8723 18717
rect 9861 18751 9919 18757
rect 9861 18717 9873 18751
rect 9907 18717 9919 18751
rect 10042 18748 10048 18760
rect 10003 18720 10048 18748
rect 9861 18711 9919 18717
rect 7190 18640 7196 18692
rect 7248 18680 7254 18692
rect 8113 18683 8171 18689
rect 8113 18680 8125 18683
rect 7248 18652 8125 18680
rect 7248 18640 7254 18652
rect 8113 18649 8125 18652
rect 8159 18649 8171 18683
rect 8113 18643 8171 18649
rect 5776 18584 6776 18612
rect 5776 18572 5782 18584
rect 6822 18572 6828 18624
rect 6880 18572 6886 18624
rect 6914 18572 6920 18624
rect 6972 18612 6978 18624
rect 8680 18612 8708 18711
rect 10042 18708 10048 18720
rect 10100 18708 10106 18760
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 9030 18640 9036 18692
rect 9088 18680 9094 18692
rect 10612 18680 10640 18711
rect 11790 18708 11796 18760
rect 11848 18748 11854 18760
rect 17494 18748 17500 18760
rect 11848 18720 17500 18748
rect 11848 18708 11854 18720
rect 17494 18708 17500 18720
rect 17552 18748 17558 18760
rect 18598 18748 18604 18760
rect 17552 18720 18604 18748
rect 17552 18708 17558 18720
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 18708 18748 18736 18788
rect 18877 18785 18889 18819
rect 18923 18816 18935 18819
rect 19153 18819 19211 18825
rect 18923 18788 19104 18816
rect 18923 18785 18935 18788
rect 18877 18779 18935 18785
rect 18708 18720 19012 18748
rect 18984 18692 19012 18720
rect 12802 18680 12808 18692
rect 9088 18652 10640 18680
rect 12406 18652 12808 18680
rect 9088 18640 9094 18652
rect 6972 18584 8708 18612
rect 6972 18572 6978 18584
rect 9766 18572 9772 18624
rect 9824 18612 9830 18624
rect 12406 18612 12434 18652
rect 12802 18640 12808 18652
rect 12860 18640 12866 18692
rect 14642 18640 14648 18692
rect 14700 18680 14706 18692
rect 17586 18680 17592 18692
rect 14700 18652 17592 18680
rect 14700 18640 14706 18652
rect 17586 18640 17592 18652
rect 17644 18680 17650 18692
rect 17681 18683 17739 18689
rect 17681 18680 17693 18683
rect 17644 18652 17693 18680
rect 17644 18640 17650 18652
rect 17681 18649 17693 18652
rect 17727 18649 17739 18683
rect 18690 18680 18696 18692
rect 18651 18652 18696 18680
rect 17681 18643 17739 18649
rect 18690 18640 18696 18652
rect 18748 18640 18754 18692
rect 18966 18680 18972 18692
rect 18879 18652 18972 18680
rect 18966 18640 18972 18652
rect 19024 18640 19030 18692
rect 19076 18680 19104 18788
rect 19153 18785 19165 18819
rect 19199 18785 19211 18819
rect 19153 18779 19211 18785
rect 19429 18819 19487 18825
rect 19429 18785 19441 18819
rect 19475 18785 19487 18819
rect 19886 18816 19892 18828
rect 19847 18788 19892 18816
rect 19429 18779 19487 18785
rect 19168 18748 19196 18779
rect 19886 18776 19892 18788
rect 19944 18776 19950 18828
rect 19978 18776 19984 18828
rect 20036 18816 20042 18828
rect 20456 18825 20484 18856
rect 20530 18844 20536 18856
rect 20588 18844 20594 18896
rect 21177 18887 21235 18893
rect 21177 18853 21189 18887
rect 21223 18884 21235 18887
rect 21266 18884 21272 18896
rect 21223 18856 21272 18884
rect 21223 18853 21235 18856
rect 21177 18847 21235 18853
rect 21266 18844 21272 18856
rect 21324 18844 21330 18896
rect 20441 18819 20499 18825
rect 20036 18788 20081 18816
rect 20036 18776 20042 18788
rect 20441 18785 20453 18819
rect 20487 18785 20499 18819
rect 20622 18816 20628 18828
rect 20583 18788 20628 18816
rect 20441 18779 20499 18785
rect 20622 18776 20628 18788
rect 20680 18776 20686 18828
rect 20990 18816 20996 18828
rect 20951 18788 20996 18816
rect 20990 18776 20996 18788
rect 21048 18776 21054 18828
rect 21358 18816 21364 18828
rect 21319 18788 21364 18816
rect 21358 18776 21364 18788
rect 21416 18776 21422 18828
rect 21542 18816 21548 18828
rect 21503 18788 21548 18816
rect 21542 18776 21548 18788
rect 21600 18776 21606 18828
rect 19334 18748 19340 18760
rect 19168 18720 19340 18748
rect 19334 18708 19340 18720
rect 19392 18748 19398 18760
rect 20346 18748 20352 18760
rect 19392 18720 20352 18748
rect 19392 18708 19398 18720
rect 20346 18708 20352 18720
rect 20404 18708 20410 18760
rect 19076 18652 19472 18680
rect 12894 18612 12900 18624
rect 9824 18584 12434 18612
rect 12855 18584 12900 18612
rect 9824 18572 9830 18584
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 16574 18572 16580 18624
rect 16632 18612 16638 18624
rect 17037 18615 17095 18621
rect 17037 18612 17049 18615
rect 16632 18584 17049 18612
rect 16632 18572 16638 18584
rect 17037 18581 17049 18584
rect 17083 18612 17095 18615
rect 17218 18612 17224 18624
rect 17083 18584 17224 18612
rect 17083 18581 17095 18584
rect 17037 18575 17095 18581
rect 17218 18572 17224 18584
rect 17276 18572 17282 18624
rect 17954 18612 17960 18624
rect 17867 18584 17960 18612
rect 17954 18572 17960 18584
rect 18012 18612 18018 18624
rect 19150 18612 19156 18624
rect 18012 18584 19156 18612
rect 18012 18572 18018 18584
rect 19150 18572 19156 18584
rect 19208 18572 19214 18624
rect 19444 18612 19472 18652
rect 19518 18640 19524 18692
rect 19576 18680 19582 18692
rect 20257 18683 20315 18689
rect 20257 18680 20269 18683
rect 19576 18652 20269 18680
rect 19576 18640 19582 18652
rect 20257 18649 20269 18652
rect 20303 18649 20315 18683
rect 20257 18643 20315 18649
rect 19978 18612 19984 18624
rect 19444 18584 19984 18612
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 1854 18408 1860 18420
rect 1815 18380 1860 18408
rect 1854 18368 1860 18380
rect 1912 18368 1918 18420
rect 1946 18368 1952 18420
rect 2004 18408 2010 18420
rect 2685 18411 2743 18417
rect 2685 18408 2697 18411
rect 2004 18380 2697 18408
rect 2004 18368 2010 18380
rect 2685 18377 2697 18380
rect 2731 18377 2743 18411
rect 2685 18371 2743 18377
rect 2866 18368 2872 18420
rect 2924 18408 2930 18420
rect 5166 18408 5172 18420
rect 2924 18380 5172 18408
rect 2924 18368 2930 18380
rect 5166 18368 5172 18380
rect 5224 18368 5230 18420
rect 5445 18411 5503 18417
rect 5445 18377 5457 18411
rect 5491 18408 5503 18411
rect 6454 18408 6460 18420
rect 5491 18380 6460 18408
rect 5491 18377 5503 18380
rect 5445 18371 5503 18377
rect 6454 18368 6460 18380
rect 6512 18368 6518 18420
rect 8202 18408 8208 18420
rect 8163 18380 8208 18408
rect 8202 18368 8208 18380
rect 8260 18368 8266 18420
rect 13814 18408 13820 18420
rect 8312 18380 13820 18408
rect 2133 18343 2191 18349
rect 2133 18309 2145 18343
rect 2179 18309 2191 18343
rect 4154 18340 4160 18352
rect 2133 18303 2191 18309
rect 3804 18312 4160 18340
rect 1581 18207 1639 18213
rect 1581 18173 1593 18207
rect 1627 18204 1639 18207
rect 2148 18204 2176 18303
rect 3234 18232 3240 18284
rect 3292 18272 3298 18284
rect 3804 18281 3832 18312
rect 4154 18300 4160 18312
rect 4212 18340 4218 18352
rect 4212 18312 4568 18340
rect 4212 18300 4218 18312
rect 3605 18275 3663 18281
rect 3605 18272 3617 18275
rect 3292 18244 3617 18272
rect 3292 18232 3298 18244
rect 3605 18241 3617 18244
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 3789 18275 3847 18281
rect 3789 18241 3801 18275
rect 3835 18241 3847 18275
rect 3789 18235 3847 18241
rect 4338 18232 4344 18284
rect 4396 18272 4402 18284
rect 4540 18281 4568 18312
rect 4433 18275 4491 18281
rect 4433 18272 4445 18275
rect 4396 18244 4445 18272
rect 4396 18232 4402 18244
rect 4433 18241 4445 18244
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 4525 18275 4583 18281
rect 4525 18241 4537 18275
rect 4571 18272 4583 18275
rect 4982 18272 4988 18284
rect 4571 18244 4988 18272
rect 4571 18241 4583 18244
rect 4525 18235 4583 18241
rect 4982 18232 4988 18244
rect 5040 18232 5046 18284
rect 5721 18275 5779 18281
rect 5721 18241 5733 18275
rect 5767 18272 5779 18275
rect 6638 18272 6644 18284
rect 5767 18244 6644 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 6638 18232 6644 18244
rect 6696 18272 6702 18284
rect 7009 18275 7067 18281
rect 7009 18272 7021 18275
rect 6696 18244 7021 18272
rect 6696 18232 6702 18244
rect 7009 18241 7021 18244
rect 7055 18272 7067 18275
rect 7561 18275 7619 18281
rect 7561 18272 7573 18275
rect 7055 18244 7573 18272
rect 7055 18241 7067 18244
rect 7009 18235 7067 18241
rect 7561 18241 7573 18244
rect 7607 18241 7619 18275
rect 8312 18272 8340 18380
rect 13814 18368 13820 18380
rect 13872 18368 13878 18420
rect 14645 18411 14703 18417
rect 14645 18377 14657 18411
rect 14691 18408 14703 18411
rect 15654 18408 15660 18420
rect 14691 18380 15660 18408
rect 14691 18377 14703 18380
rect 14645 18371 14703 18377
rect 15654 18368 15660 18380
rect 15712 18368 15718 18420
rect 16577 18411 16635 18417
rect 16577 18377 16589 18411
rect 16623 18408 16635 18411
rect 17402 18408 17408 18420
rect 16623 18380 17408 18408
rect 16623 18377 16635 18380
rect 16577 18371 16635 18377
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 19334 18408 19340 18420
rect 19295 18380 19340 18408
rect 19334 18368 19340 18380
rect 19392 18368 19398 18420
rect 19610 18408 19616 18420
rect 19571 18380 19616 18408
rect 19610 18368 19616 18380
rect 19668 18368 19674 18420
rect 19889 18411 19947 18417
rect 19889 18377 19901 18411
rect 19935 18408 19947 18411
rect 20162 18408 20168 18420
rect 19935 18380 20168 18408
rect 19935 18377 19947 18380
rect 19889 18371 19947 18377
rect 20162 18368 20168 18380
rect 20220 18368 20226 18420
rect 20257 18411 20315 18417
rect 20257 18377 20269 18411
rect 20303 18408 20315 18411
rect 20622 18408 20628 18420
rect 20303 18380 20628 18408
rect 20303 18377 20315 18380
rect 20257 18371 20315 18377
rect 20622 18368 20628 18380
rect 20680 18368 20686 18420
rect 10873 18343 10931 18349
rect 10873 18309 10885 18343
rect 10919 18340 10931 18343
rect 11146 18340 11152 18352
rect 10919 18312 11152 18340
rect 10919 18309 10931 18312
rect 10873 18303 10931 18309
rect 11146 18300 11152 18312
rect 11204 18340 11210 18352
rect 11698 18340 11704 18352
rect 11204 18312 11704 18340
rect 11204 18300 11210 18312
rect 11698 18300 11704 18312
rect 11756 18300 11762 18352
rect 16025 18343 16083 18349
rect 16025 18309 16037 18343
rect 16071 18309 16083 18343
rect 16025 18303 16083 18309
rect 19061 18343 19119 18349
rect 19061 18309 19073 18343
rect 19107 18340 19119 18343
rect 19794 18340 19800 18352
rect 19107 18312 19800 18340
rect 19107 18309 19119 18312
rect 19061 18303 19119 18309
rect 7561 18235 7619 18241
rect 7668 18244 8340 18272
rect 8481 18275 8539 18281
rect 1627 18176 2176 18204
rect 2317 18207 2375 18213
rect 1627 18173 1639 18176
rect 1581 18167 1639 18173
rect 2317 18173 2329 18207
rect 2363 18204 2375 18207
rect 2593 18207 2651 18213
rect 2363 18176 2544 18204
rect 2363 18173 2375 18176
rect 2317 18167 2375 18173
rect 1949 18139 2007 18145
rect 1949 18105 1961 18139
rect 1995 18136 2007 18139
rect 1995 18108 2452 18136
rect 1995 18105 2007 18108
rect 1949 18099 2007 18105
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 2424 18077 2452 18108
rect 2409 18071 2467 18077
rect 2409 18037 2421 18071
rect 2455 18037 2467 18071
rect 2516 18068 2544 18176
rect 2593 18173 2605 18207
rect 2639 18173 2651 18207
rect 2593 18167 2651 18173
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 5350 18204 5356 18216
rect 2915 18176 5356 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 2608 18136 2636 18167
rect 5350 18164 5356 18176
rect 5408 18164 5414 18216
rect 5905 18207 5963 18213
rect 5905 18173 5917 18207
rect 5951 18204 5963 18207
rect 6270 18204 6276 18216
rect 5951 18176 6276 18204
rect 5951 18173 5963 18176
rect 5905 18167 5963 18173
rect 6270 18164 6276 18176
rect 6328 18164 6334 18216
rect 6454 18164 6460 18216
rect 6512 18204 6518 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6512 18176 6837 18204
rect 6512 18164 6518 18176
rect 6825 18173 6837 18176
rect 6871 18204 6883 18207
rect 7668 18204 7696 18244
rect 8481 18241 8493 18275
rect 8527 18272 8539 18275
rect 8846 18272 8852 18284
rect 8527 18244 8852 18272
rect 8527 18241 8539 18244
rect 8481 18235 8539 18241
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 6871 18176 7696 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 7742 18164 7748 18216
rect 7800 18204 7806 18216
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 7800 18176 7849 18204
rect 7800 18164 7806 18176
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 8570 18164 8576 18216
rect 8628 18204 8634 18216
rect 8665 18207 8723 18213
rect 8665 18204 8677 18207
rect 8628 18176 8677 18204
rect 8628 18164 8634 18176
rect 8665 18173 8677 18176
rect 8711 18173 8723 18207
rect 8665 18167 8723 18173
rect 9030 18164 9036 18216
rect 9088 18204 9094 18216
rect 9493 18207 9551 18213
rect 9493 18204 9505 18207
rect 9088 18176 9505 18204
rect 9088 18164 9094 18176
rect 9493 18173 9505 18176
rect 9539 18173 9551 18207
rect 9493 18167 9551 18173
rect 9582 18164 9588 18216
rect 9640 18204 9646 18216
rect 11606 18204 11612 18216
rect 9640 18176 11612 18204
rect 9640 18164 9646 18176
rect 11606 18164 11612 18176
rect 11664 18164 11670 18216
rect 11701 18207 11759 18213
rect 11701 18173 11713 18207
rect 11747 18204 11759 18207
rect 12434 18204 12440 18216
rect 11747 18176 12440 18204
rect 11747 18173 11759 18176
rect 11701 18167 11759 18173
rect 12434 18164 12440 18176
rect 12492 18164 12498 18216
rect 14458 18204 14464 18216
rect 14419 18176 14464 18204
rect 14458 18164 14464 18176
rect 14516 18164 14522 18216
rect 15838 18204 15844 18216
rect 15799 18176 15844 18204
rect 15838 18164 15844 18176
rect 15896 18164 15902 18216
rect 16040 18204 16068 18303
rect 19794 18300 19800 18312
rect 19852 18300 19858 18352
rect 20533 18343 20591 18349
rect 20533 18309 20545 18343
rect 20579 18340 20591 18343
rect 20990 18340 20996 18352
rect 20579 18312 20996 18340
rect 20579 18309 20591 18312
rect 20533 18303 20591 18309
rect 20990 18300 20996 18312
rect 21048 18300 21054 18352
rect 21174 18340 21180 18352
rect 21135 18312 21180 18340
rect 21174 18300 21180 18312
rect 21232 18300 21238 18352
rect 18966 18232 18972 18284
rect 19024 18272 19030 18284
rect 19024 18244 20392 18272
rect 19024 18232 19030 18244
rect 16393 18207 16451 18213
rect 16393 18204 16405 18207
rect 16040 18176 16405 18204
rect 16393 18173 16405 18176
rect 16439 18173 16451 18207
rect 16393 18167 16451 18173
rect 18785 18207 18843 18213
rect 18785 18173 18797 18207
rect 18831 18204 18843 18207
rect 18877 18207 18935 18213
rect 18877 18204 18889 18207
rect 18831 18176 18889 18204
rect 18831 18173 18843 18176
rect 18785 18167 18843 18173
rect 18877 18173 18889 18176
rect 18923 18173 18935 18207
rect 19702 18204 19708 18216
rect 19663 18176 19708 18204
rect 18877 18167 18935 18173
rect 3602 18136 3608 18148
rect 2608 18108 3608 18136
rect 3602 18096 3608 18108
rect 3660 18096 3666 18148
rect 4062 18096 4068 18148
rect 4120 18136 4126 18148
rect 8938 18136 8944 18148
rect 4120 18108 8944 18136
rect 4120 18096 4126 18108
rect 2958 18068 2964 18080
rect 2516 18040 2964 18068
rect 2409 18031 2467 18037
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 3142 18068 3148 18080
rect 3103 18040 3148 18068
rect 3142 18028 3148 18040
rect 3200 18028 3206 18080
rect 3418 18028 3424 18080
rect 3476 18068 3482 18080
rect 3513 18071 3571 18077
rect 3513 18068 3525 18071
rect 3476 18040 3525 18068
rect 3476 18028 3482 18040
rect 3513 18037 3525 18040
rect 3559 18068 3571 18071
rect 3694 18068 3700 18080
rect 3559 18040 3700 18068
rect 3559 18037 3571 18040
rect 3513 18031 3571 18037
rect 3694 18028 3700 18040
rect 3752 18028 3758 18080
rect 3970 18068 3976 18080
rect 3931 18040 3976 18068
rect 3970 18028 3976 18040
rect 4028 18028 4034 18080
rect 4341 18071 4399 18077
rect 4341 18037 4353 18071
rect 4387 18068 4399 18071
rect 5166 18068 5172 18080
rect 4387 18040 5172 18068
rect 4387 18037 4399 18040
rect 4341 18031 4399 18037
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 5813 18071 5871 18077
rect 5813 18037 5825 18071
rect 5859 18068 5871 18071
rect 6086 18068 6092 18080
rect 5859 18040 6092 18068
rect 5859 18037 5871 18040
rect 5813 18031 5871 18037
rect 6086 18028 6092 18040
rect 6144 18028 6150 18080
rect 6270 18068 6276 18080
rect 6231 18040 6276 18068
rect 6270 18028 6276 18040
rect 6328 18028 6334 18080
rect 6454 18068 6460 18080
rect 6415 18040 6460 18068
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 6914 18028 6920 18080
rect 6972 18068 6978 18080
rect 6972 18040 7017 18068
rect 6972 18028 6978 18040
rect 7650 18028 7656 18080
rect 7708 18068 7714 18080
rect 8588 18077 8616 18108
rect 8938 18096 8944 18108
rect 8996 18096 9002 18148
rect 9760 18139 9818 18145
rect 9760 18105 9772 18139
rect 9806 18136 9818 18139
rect 10594 18136 10600 18148
rect 9806 18108 10600 18136
rect 9806 18105 9818 18108
rect 9760 18099 9818 18105
rect 10594 18096 10600 18108
rect 10652 18096 10658 18148
rect 11882 18096 11888 18148
rect 11940 18145 11946 18148
rect 11940 18139 12004 18145
rect 11940 18105 11958 18139
rect 11992 18105 12004 18139
rect 18892 18136 18920 18167
rect 19702 18164 19708 18176
rect 19760 18164 19766 18216
rect 19886 18164 19892 18216
rect 19944 18204 19950 18216
rect 20364 18213 20392 18244
rect 20438 18232 20444 18284
rect 20496 18272 20502 18284
rect 20496 18244 21404 18272
rect 20496 18232 20502 18244
rect 21376 18213 21404 18244
rect 20073 18207 20131 18213
rect 20073 18204 20085 18207
rect 19944 18176 20085 18204
rect 19944 18164 19950 18176
rect 20073 18173 20085 18176
rect 20119 18173 20131 18207
rect 20073 18167 20131 18173
rect 20349 18207 20407 18213
rect 20349 18173 20361 18207
rect 20395 18173 20407 18207
rect 20625 18207 20683 18213
rect 20625 18204 20637 18207
rect 20349 18167 20407 18173
rect 20456 18176 20637 18204
rect 18966 18136 18972 18148
rect 18892 18108 18972 18136
rect 11940 18099 12004 18105
rect 11940 18096 11946 18099
rect 18966 18096 18972 18108
rect 19024 18096 19030 18148
rect 19978 18096 19984 18148
rect 20036 18136 20042 18148
rect 20456 18136 20484 18176
rect 20625 18173 20637 18176
rect 20671 18173 20683 18207
rect 20625 18167 20683 18173
rect 21361 18207 21419 18213
rect 21361 18173 21373 18207
rect 21407 18173 21419 18207
rect 21361 18167 21419 18173
rect 20993 18139 21051 18145
rect 20993 18136 21005 18139
rect 20036 18108 20484 18136
rect 20640 18108 21005 18136
rect 20036 18096 20042 18108
rect 20640 18080 20668 18108
rect 20993 18105 21005 18108
rect 21039 18105 21051 18139
rect 21542 18136 21548 18148
rect 21503 18108 21548 18136
rect 20993 18099 21051 18105
rect 21542 18096 21548 18108
rect 21600 18096 21606 18148
rect 7745 18071 7803 18077
rect 7745 18068 7757 18071
rect 7708 18040 7757 18068
rect 7708 18028 7714 18040
rect 7745 18037 7757 18040
rect 7791 18037 7803 18071
rect 7745 18031 7803 18037
rect 8573 18071 8631 18077
rect 8573 18037 8585 18071
rect 8619 18037 8631 18071
rect 8573 18031 8631 18037
rect 9033 18071 9091 18077
rect 9033 18037 9045 18071
rect 9079 18068 9091 18071
rect 10410 18068 10416 18080
rect 9079 18040 10416 18068
rect 9079 18037 9091 18040
rect 9033 18031 9091 18037
rect 10410 18028 10416 18040
rect 10468 18028 10474 18080
rect 10962 18028 10968 18080
rect 11020 18068 11026 18080
rect 11020 18040 11065 18068
rect 11020 18028 11026 18040
rect 12526 18028 12532 18080
rect 12584 18068 12590 18080
rect 13081 18071 13139 18077
rect 13081 18068 13093 18071
rect 12584 18040 13093 18068
rect 12584 18028 12590 18040
rect 13081 18037 13093 18040
rect 13127 18037 13139 18071
rect 13081 18031 13139 18037
rect 20622 18028 20628 18080
rect 20680 18028 20686 18080
rect 20809 18071 20867 18077
rect 20809 18037 20821 18071
rect 20855 18068 20867 18071
rect 21266 18068 21272 18080
rect 20855 18040 21272 18068
rect 20855 18037 20867 18040
rect 20809 18031 20867 18037
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 2593 17867 2651 17873
rect 2593 17833 2605 17867
rect 2639 17864 2651 17867
rect 3142 17864 3148 17876
rect 2639 17836 3148 17864
rect 2639 17833 2651 17836
rect 2593 17827 2651 17833
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3375 17836 4077 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 4246 17824 4252 17876
rect 4304 17864 4310 17876
rect 4433 17867 4491 17873
rect 4433 17864 4445 17867
rect 4304 17836 4445 17864
rect 4304 17824 4310 17836
rect 4433 17833 4445 17836
rect 4479 17833 4491 17867
rect 4433 17827 4491 17833
rect 1581 17799 1639 17805
rect 1581 17765 1593 17799
rect 1627 17796 1639 17799
rect 3234 17796 3240 17808
rect 1627 17768 3240 17796
rect 1627 17765 1639 17768
rect 1581 17759 1639 17765
rect 3234 17756 3240 17768
rect 3292 17756 3298 17808
rect 3421 17799 3479 17805
rect 3421 17765 3433 17799
rect 3467 17796 3479 17799
rect 3970 17796 3976 17808
rect 3467 17768 3976 17796
rect 3467 17765 3479 17768
rect 3421 17759 3479 17765
rect 3970 17756 3976 17768
rect 4028 17756 4034 17808
rect 4448 17796 4476 17827
rect 4522 17824 4528 17876
rect 4580 17864 4586 17876
rect 4890 17864 4896 17876
rect 4580 17836 4625 17864
rect 4851 17836 4896 17864
rect 4580 17824 4586 17836
rect 4890 17824 4896 17836
rect 4948 17824 4954 17876
rect 5258 17864 5264 17876
rect 5219 17836 5264 17864
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 6365 17867 6423 17873
rect 6365 17833 6377 17867
rect 6411 17864 6423 17867
rect 6454 17864 6460 17876
rect 6411 17836 6460 17864
rect 6411 17833 6423 17836
rect 6365 17827 6423 17833
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 6730 17824 6736 17876
rect 6788 17864 6794 17876
rect 6825 17867 6883 17873
rect 6825 17864 6837 17867
rect 6788 17836 6837 17864
rect 6788 17824 6794 17836
rect 6825 17833 6837 17836
rect 6871 17833 6883 17867
rect 6825 17827 6883 17833
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7009 17867 7067 17873
rect 7009 17864 7021 17867
rect 6972 17836 7021 17864
rect 6972 17824 6978 17836
rect 7009 17833 7021 17836
rect 7055 17833 7067 17867
rect 7009 17827 7067 17833
rect 7190 17824 7196 17876
rect 7248 17864 7254 17876
rect 7377 17867 7435 17873
rect 7377 17864 7389 17867
rect 7248 17836 7389 17864
rect 7248 17824 7254 17836
rect 7377 17833 7389 17836
rect 7423 17864 7435 17867
rect 7558 17864 7564 17876
rect 7423 17836 7564 17864
rect 7423 17833 7435 17836
rect 7377 17827 7435 17833
rect 7558 17824 7564 17836
rect 7616 17824 7622 17876
rect 7742 17824 7748 17876
rect 7800 17864 7806 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 7800 17836 7849 17864
rect 7800 17824 7806 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 8202 17864 8208 17876
rect 8163 17836 8208 17864
rect 7837 17827 7895 17833
rect 8202 17824 8208 17836
rect 8260 17864 8266 17876
rect 9125 17867 9183 17873
rect 9125 17864 9137 17867
rect 8260 17836 9137 17864
rect 8260 17824 8266 17836
rect 9125 17833 9137 17836
rect 9171 17864 9183 17867
rect 9766 17864 9772 17876
rect 9171 17836 9772 17864
rect 9171 17833 9183 17836
rect 9125 17827 9183 17833
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 9953 17867 10011 17873
rect 9953 17833 9965 17867
rect 9999 17864 10011 17867
rect 10042 17864 10048 17876
rect 9999 17836 10048 17864
rect 9999 17833 10011 17836
rect 9953 17827 10011 17833
rect 10042 17824 10048 17836
rect 10100 17824 10106 17876
rect 10410 17864 10416 17876
rect 10371 17836 10416 17864
rect 10410 17824 10416 17836
rect 10468 17824 10474 17876
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 10870 17864 10876 17876
rect 10827 17836 10876 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 11974 17864 11980 17876
rect 11164 17836 11980 17864
rect 5534 17796 5540 17808
rect 4448 17768 5540 17796
rect 5534 17756 5540 17768
rect 5592 17756 5598 17808
rect 5994 17756 6000 17808
rect 6052 17796 6058 17808
rect 8754 17796 8760 17808
rect 6052 17768 8760 17796
rect 6052 17756 6058 17768
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 11164 17805 11192 17836
rect 11974 17824 11980 17836
rect 12032 17824 12038 17876
rect 12066 17824 12072 17876
rect 12124 17864 12130 17876
rect 12345 17867 12403 17873
rect 12345 17864 12357 17867
rect 12124 17836 12357 17864
rect 12124 17824 12130 17836
rect 12345 17833 12357 17836
rect 12391 17833 12403 17867
rect 12345 17827 12403 17833
rect 13817 17867 13875 17873
rect 13817 17833 13829 17867
rect 13863 17864 13875 17867
rect 14458 17864 14464 17876
rect 13863 17836 14464 17864
rect 13863 17833 13875 17836
rect 13817 17827 13875 17833
rect 14458 17824 14464 17836
rect 14516 17824 14522 17876
rect 15105 17867 15163 17873
rect 15105 17833 15117 17867
rect 15151 17864 15163 17867
rect 15473 17867 15531 17873
rect 15473 17864 15485 17867
rect 15151 17836 15485 17864
rect 15151 17833 15163 17836
rect 15105 17827 15163 17833
rect 15473 17833 15485 17836
rect 15519 17833 15531 17867
rect 15473 17827 15531 17833
rect 15933 17867 15991 17873
rect 15933 17833 15945 17867
rect 15979 17864 15991 17867
rect 16485 17867 16543 17873
rect 16485 17864 16497 17867
rect 15979 17836 16497 17864
rect 15979 17833 15991 17836
rect 15933 17827 15991 17833
rect 16485 17833 16497 17836
rect 16531 17833 16543 17867
rect 16485 17827 16543 17833
rect 19429 17867 19487 17873
rect 19429 17833 19441 17867
rect 19475 17864 19487 17867
rect 19702 17864 19708 17876
rect 19475 17836 19708 17864
rect 19475 17833 19487 17836
rect 19429 17827 19487 17833
rect 19702 17824 19708 17836
rect 19760 17824 19766 17876
rect 20349 17867 20407 17873
rect 20349 17833 20361 17867
rect 20395 17864 20407 17867
rect 20438 17864 20444 17876
rect 20395 17836 20444 17864
rect 20395 17833 20407 17836
rect 20349 17827 20407 17833
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 20622 17864 20628 17876
rect 20583 17836 20628 17864
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 11149 17799 11207 17805
rect 11149 17796 11161 17799
rect 9876 17768 11161 17796
rect 9876 17740 9904 17768
rect 11149 17765 11161 17768
rect 11195 17765 11207 17799
rect 14737 17799 14795 17805
rect 14737 17796 14749 17799
rect 11149 17759 11207 17765
rect 11348 17768 12112 17796
rect 1946 17728 1952 17740
rect 1907 17700 1952 17728
rect 1946 17688 1952 17700
rect 2004 17688 2010 17740
rect 2501 17731 2559 17737
rect 2501 17697 2513 17731
rect 2547 17728 2559 17731
rect 4154 17728 4160 17740
rect 2547 17700 4160 17728
rect 2547 17697 2559 17700
rect 2501 17691 2559 17697
rect 4154 17688 4160 17700
rect 4212 17688 4218 17740
rect 6270 17688 6276 17740
rect 6328 17728 6334 17740
rect 6457 17731 6515 17737
rect 6457 17728 6469 17731
rect 6328 17700 6469 17728
rect 6328 17688 6334 17700
rect 6457 17697 6469 17700
rect 6503 17697 6515 17731
rect 6457 17691 6515 17697
rect 7469 17731 7527 17737
rect 7469 17697 7481 17731
rect 7515 17728 7527 17731
rect 9858 17728 9864 17740
rect 7515 17700 8984 17728
rect 9819 17700 9864 17728
rect 7515 17697 7527 17700
rect 7469 17691 7527 17697
rect 2406 17620 2412 17672
rect 2464 17660 2470 17672
rect 2685 17663 2743 17669
rect 2685 17660 2697 17663
rect 2464 17632 2697 17660
rect 2464 17620 2470 17632
rect 2685 17629 2697 17632
rect 2731 17660 2743 17663
rect 3513 17663 3571 17669
rect 2731 17632 3188 17660
rect 2731 17629 2743 17632
rect 2685 17623 2743 17629
rect 1762 17592 1768 17604
rect 1723 17564 1768 17592
rect 1762 17552 1768 17564
rect 1820 17552 1826 17604
rect 2590 17552 2596 17604
rect 2648 17592 2654 17604
rect 3160 17592 3188 17632
rect 3513 17629 3525 17663
rect 3559 17629 3571 17663
rect 3513 17623 3571 17629
rect 3528 17592 3556 17623
rect 3602 17620 3608 17672
rect 3660 17660 3666 17672
rect 3973 17663 4031 17669
rect 3973 17660 3985 17663
rect 3660 17632 3985 17660
rect 3660 17620 3666 17632
rect 3973 17629 3985 17632
rect 4019 17660 4031 17663
rect 4062 17660 4068 17672
rect 4019 17632 4068 17660
rect 4019 17629 4031 17632
rect 3973 17623 4031 17629
rect 4062 17620 4068 17632
rect 4120 17620 4126 17672
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17660 4767 17663
rect 4982 17660 4988 17672
rect 4755 17632 4988 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 5353 17663 5411 17669
rect 5353 17629 5365 17663
rect 5399 17629 5411 17663
rect 5353 17623 5411 17629
rect 5368 17592 5396 17623
rect 5442 17620 5448 17672
rect 5500 17660 5506 17672
rect 5994 17660 6000 17672
rect 5500 17632 5545 17660
rect 5644 17632 6000 17660
rect 5500 17620 5506 17632
rect 2648 17564 3096 17592
rect 3160 17564 3556 17592
rect 3620 17564 5396 17592
rect 2648 17552 2654 17564
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 2133 17527 2191 17533
rect 2133 17493 2145 17527
rect 2179 17524 2191 17527
rect 2222 17524 2228 17536
rect 2179 17496 2228 17524
rect 2179 17493 2191 17496
rect 2133 17487 2191 17493
rect 2222 17484 2228 17496
rect 2280 17484 2286 17536
rect 2314 17484 2320 17536
rect 2372 17524 2378 17536
rect 2961 17527 3019 17533
rect 2961 17524 2973 17527
rect 2372 17496 2973 17524
rect 2372 17484 2378 17496
rect 2961 17493 2973 17496
rect 3007 17493 3019 17527
rect 3068 17524 3096 17564
rect 3620 17524 3648 17564
rect 3068 17496 3648 17524
rect 2961 17487 3019 17493
rect 3694 17484 3700 17536
rect 3752 17524 3758 17536
rect 5644 17524 5672 17632
rect 5994 17620 6000 17632
rect 6052 17620 6058 17672
rect 6178 17660 6184 17672
rect 6139 17632 6184 17660
rect 6178 17620 6184 17632
rect 6236 17620 6242 17672
rect 7558 17660 7564 17672
rect 7519 17632 7564 17660
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 8956 17669 8984 17700
rect 9858 17688 9864 17700
rect 9916 17688 9922 17740
rect 10318 17728 10324 17740
rect 10279 17700 10324 17728
rect 10318 17688 10324 17700
rect 10376 17688 10382 17740
rect 11348 17728 11376 17768
rect 11974 17728 11980 17740
rect 10796 17700 11376 17728
rect 11935 17700 11980 17728
rect 8297 17663 8355 17669
rect 8297 17660 8309 17663
rect 7800 17632 8309 17660
rect 7800 17620 7806 17632
rect 8297 17629 8309 17632
rect 8343 17629 8355 17663
rect 8297 17623 8355 17629
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17629 8447 17663
rect 8389 17623 8447 17629
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17660 8999 17663
rect 9766 17660 9772 17672
rect 8987 17632 9772 17660
rect 8987 17629 8999 17632
rect 8941 17623 8999 17629
rect 7576 17592 7604 17620
rect 8404 17592 8432 17623
rect 9766 17620 9772 17632
rect 9824 17620 9830 17672
rect 10594 17660 10600 17672
rect 10555 17632 10600 17660
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 10796 17660 10824 17700
rect 11974 17688 11980 17700
rect 12032 17688 12038 17740
rect 12084 17728 12112 17768
rect 13096 17768 14749 17796
rect 13096 17728 13124 17768
rect 14737 17765 14749 17768
rect 14783 17765 14795 17799
rect 14737 17759 14795 17765
rect 19797 17799 19855 17805
rect 19797 17765 19809 17799
rect 19843 17796 19855 17799
rect 19843 17768 20944 17796
rect 19843 17765 19855 17768
rect 19797 17759 19855 17765
rect 20916 17740 20944 17768
rect 12084 17700 13124 17728
rect 13173 17731 13231 17737
rect 13173 17697 13185 17731
rect 13219 17728 13231 17731
rect 13538 17728 13544 17740
rect 13219 17700 13544 17728
rect 13219 17697 13231 17700
rect 13173 17691 13231 17697
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 13633 17731 13691 17737
rect 13633 17697 13645 17731
rect 13679 17697 13691 17731
rect 15286 17728 15292 17740
rect 13633 17691 13691 17697
rect 14568 17700 15292 17728
rect 10704 17632 10824 17660
rect 10704 17592 10732 17632
rect 11146 17620 11152 17672
rect 11204 17660 11210 17672
rect 11241 17663 11299 17669
rect 11241 17660 11253 17663
rect 11204 17632 11253 17660
rect 11204 17620 11210 17632
rect 11241 17629 11253 17632
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 11330 17620 11336 17672
rect 11388 17660 11394 17672
rect 11698 17660 11704 17672
rect 11388 17632 11433 17660
rect 11659 17632 11704 17660
rect 11388 17620 11394 17632
rect 11698 17620 11704 17632
rect 11756 17620 11762 17672
rect 11885 17663 11943 17669
rect 11885 17629 11897 17663
rect 11931 17629 11943 17663
rect 11885 17623 11943 17629
rect 12897 17663 12955 17669
rect 12897 17629 12909 17663
rect 12943 17629 12955 17663
rect 13078 17660 13084 17672
rect 13039 17632 13084 17660
rect 12897 17623 12955 17629
rect 7576 17564 8432 17592
rect 8496 17564 10732 17592
rect 3752 17496 5672 17524
rect 5997 17527 6055 17533
rect 3752 17484 3758 17496
rect 5997 17493 6009 17527
rect 6043 17524 6055 17527
rect 7190 17524 7196 17536
rect 6043 17496 7196 17524
rect 6043 17493 6055 17496
rect 5997 17487 6055 17493
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 8496 17524 8524 17564
rect 10778 17552 10784 17604
rect 10836 17592 10842 17604
rect 11900 17592 11928 17623
rect 10836 17564 11928 17592
rect 10836 17552 10842 17564
rect 12342 17552 12348 17604
rect 12400 17592 12406 17604
rect 12437 17595 12495 17601
rect 12437 17592 12449 17595
rect 12400 17564 12449 17592
rect 12400 17552 12406 17564
rect 12437 17561 12449 17564
rect 12483 17561 12495 17595
rect 12912 17592 12940 17623
rect 13078 17620 13084 17632
rect 13136 17620 13142 17672
rect 13648 17660 13676 17691
rect 14568 17669 14596 17700
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 15562 17728 15568 17740
rect 15523 17700 15568 17728
rect 15562 17688 15568 17700
rect 15620 17688 15626 17740
rect 16390 17728 16396 17740
rect 16351 17700 16396 17728
rect 16390 17688 16396 17700
rect 16448 17688 16454 17740
rect 19889 17731 19947 17737
rect 19889 17697 19901 17731
rect 19935 17697 19947 17731
rect 20162 17728 20168 17740
rect 20123 17700 20168 17728
rect 19889 17691 19947 17697
rect 13556 17632 13676 17660
rect 14553 17663 14611 17669
rect 13446 17592 13452 17604
rect 12912 17564 13452 17592
rect 12437 17555 12495 17561
rect 13446 17552 13452 17564
rect 13504 17552 13510 17604
rect 13556 17601 13584 17632
rect 14553 17629 14565 17663
rect 14599 17629 14611 17663
rect 14553 17623 14611 17629
rect 14645 17663 14703 17669
rect 14645 17629 14657 17663
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 15381 17663 15439 17669
rect 15381 17629 15393 17663
rect 15427 17660 15439 17663
rect 15746 17660 15752 17672
rect 15427 17632 15752 17660
rect 15427 17629 15439 17632
rect 15381 17623 15439 17629
rect 13541 17595 13599 17601
rect 13541 17561 13553 17595
rect 13587 17561 13599 17595
rect 13541 17555 13599 17561
rect 7432 17496 8524 17524
rect 7432 17484 7438 17496
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 8665 17527 8723 17533
rect 8665 17524 8677 17527
rect 8628 17496 8677 17524
rect 8628 17484 8634 17496
rect 8665 17493 8677 17496
rect 8711 17493 8723 17527
rect 8665 17487 8723 17493
rect 9214 17484 9220 17536
rect 9272 17524 9278 17536
rect 14660 17524 14688 17623
rect 15746 17620 15752 17632
rect 15804 17620 15810 17672
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17660 16727 17663
rect 16758 17660 16764 17672
rect 16715 17632 16764 17660
rect 16715 17629 16727 17632
rect 16669 17623 16727 17629
rect 16758 17620 16764 17632
rect 16816 17620 16822 17672
rect 19904 17660 19932 17691
rect 20162 17688 20168 17700
rect 20220 17688 20226 17740
rect 20441 17731 20499 17737
rect 20441 17697 20453 17731
rect 20487 17728 20499 17731
rect 20530 17728 20536 17740
rect 20487 17700 20536 17728
rect 20487 17697 20499 17700
rect 20441 17691 20499 17697
rect 20530 17688 20536 17700
rect 20588 17688 20594 17740
rect 20898 17688 20904 17740
rect 20956 17728 20962 17740
rect 21177 17731 21235 17737
rect 21177 17728 21189 17731
rect 20956 17700 21189 17728
rect 20956 17688 20962 17700
rect 21177 17697 21189 17700
rect 21223 17697 21235 17731
rect 21177 17691 21235 17697
rect 21361 17731 21419 17737
rect 21361 17697 21373 17731
rect 21407 17728 21419 17731
rect 22005 17731 22063 17737
rect 22005 17728 22017 17731
rect 21407 17700 22017 17728
rect 21407 17697 21419 17700
rect 21361 17691 21419 17697
rect 22005 17697 22017 17700
rect 22051 17697 22063 17731
rect 22005 17691 22063 17697
rect 20346 17660 20352 17672
rect 19904 17632 20352 17660
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20993 17663 21051 17669
rect 20993 17629 21005 17663
rect 21039 17660 21051 17663
rect 21039 17632 22048 17660
rect 21039 17629 21051 17632
rect 20993 17623 21051 17629
rect 22020 17604 22048 17632
rect 15838 17552 15844 17604
rect 15896 17592 15902 17604
rect 16025 17595 16083 17601
rect 16025 17592 16037 17595
rect 15896 17564 16037 17592
rect 15896 17552 15902 17564
rect 16025 17561 16037 17564
rect 16071 17561 16083 17595
rect 21542 17592 21548 17604
rect 21503 17564 21548 17592
rect 16025 17555 16083 17561
rect 21542 17552 21548 17564
rect 21600 17552 21606 17604
rect 22002 17552 22008 17604
rect 22060 17552 22066 17604
rect 20070 17524 20076 17536
rect 9272 17496 14688 17524
rect 20031 17496 20076 17524
rect 9272 17484 9278 17496
rect 20070 17484 20076 17496
rect 20128 17484 20134 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 3326 17320 3332 17332
rect 1596 17292 3332 17320
rect 1596 17125 1624 17292
rect 3326 17280 3332 17292
rect 3384 17280 3390 17332
rect 4065 17323 4123 17329
rect 4065 17289 4077 17323
rect 4111 17320 4123 17323
rect 4338 17320 4344 17332
rect 4111 17292 4344 17320
rect 4111 17289 4123 17292
rect 4065 17283 4123 17289
rect 4338 17280 4344 17292
rect 4396 17320 4402 17332
rect 5442 17320 5448 17332
rect 4396 17292 5448 17320
rect 4396 17280 4402 17292
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 7374 17320 7380 17332
rect 5552 17292 7380 17320
rect 2590 17252 2596 17264
rect 2551 17224 2596 17252
rect 2590 17212 2596 17224
rect 2648 17212 2654 17264
rect 4154 17252 4160 17264
rect 4115 17224 4160 17252
rect 4154 17212 4160 17224
rect 4212 17212 4218 17264
rect 5552 17252 5580 17292
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 7650 17280 7656 17332
rect 7708 17320 7714 17332
rect 7929 17323 7987 17329
rect 7929 17320 7941 17323
rect 7708 17292 7941 17320
rect 7708 17280 7714 17292
rect 7929 17289 7941 17292
rect 7975 17289 7987 17323
rect 9030 17320 9036 17332
rect 7929 17283 7987 17289
rect 8772 17292 9036 17320
rect 4632 17224 5580 17252
rect 2041 17187 2099 17193
rect 2041 17153 2053 17187
rect 2087 17153 2099 17187
rect 2041 17147 2099 17153
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17184 2191 17187
rect 2314 17184 2320 17196
rect 2179 17156 2320 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17085 1639 17119
rect 1581 17079 1639 17085
rect 1762 17008 1768 17060
rect 1820 17048 1826 17060
rect 2056 17048 2084 17147
rect 2314 17144 2320 17156
rect 2372 17144 2378 17196
rect 3786 17144 3792 17196
rect 3844 17184 3850 17196
rect 4632 17193 4660 17224
rect 5718 17212 5724 17264
rect 5776 17252 5782 17264
rect 7837 17255 7895 17261
rect 5776 17224 6224 17252
rect 5776 17212 5782 17224
rect 6196 17196 6224 17224
rect 7837 17221 7849 17255
rect 7883 17252 7895 17255
rect 8386 17252 8392 17264
rect 7883 17224 8392 17252
rect 7883 17221 7895 17224
rect 7837 17215 7895 17221
rect 8386 17212 8392 17224
rect 8444 17212 8450 17264
rect 4617 17187 4675 17193
rect 4617 17184 4629 17187
rect 3844 17156 4629 17184
rect 3844 17144 3850 17156
rect 4617 17153 4629 17156
rect 4663 17153 4675 17187
rect 4617 17147 4675 17153
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17184 4859 17187
rect 4982 17184 4988 17196
rect 4847 17156 4988 17184
rect 4847 17153 4859 17156
rect 4801 17147 4859 17153
rect 4982 17144 4988 17156
rect 5040 17144 5046 17196
rect 5445 17187 5503 17193
rect 5445 17153 5457 17187
rect 5491 17184 5503 17187
rect 5810 17184 5816 17196
rect 5491 17156 5816 17184
rect 5491 17153 5503 17156
rect 5445 17147 5503 17153
rect 5810 17144 5816 17156
rect 5868 17144 5874 17196
rect 6178 17144 6184 17196
rect 6236 17184 6242 17196
rect 6457 17187 6515 17193
rect 6457 17184 6469 17187
rect 6236 17156 6469 17184
rect 6236 17144 6242 17156
rect 6457 17153 6469 17156
rect 6503 17153 6515 17187
rect 6457 17147 6515 17153
rect 7558 17144 7564 17196
rect 7616 17184 7622 17196
rect 8772 17193 8800 17292
rect 9030 17280 9036 17292
rect 9088 17280 9094 17332
rect 11241 17323 11299 17329
rect 11241 17289 11253 17323
rect 11287 17320 11299 17323
rect 11974 17320 11980 17332
rect 11287 17292 11980 17320
rect 11287 17289 11299 17292
rect 11241 17283 11299 17289
rect 11974 17280 11980 17292
rect 12032 17280 12038 17332
rect 13446 17280 13452 17332
rect 13504 17320 13510 17332
rect 13817 17323 13875 17329
rect 13817 17320 13829 17323
rect 13504 17292 13829 17320
rect 13504 17280 13510 17292
rect 13817 17289 13829 17292
rect 13863 17289 13875 17323
rect 16758 17320 16764 17332
rect 16719 17292 16764 17320
rect 13817 17283 13875 17289
rect 16758 17280 16764 17292
rect 16816 17280 16822 17332
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 21358 17320 21364 17332
rect 21039 17292 21364 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 21358 17280 21364 17292
rect 21416 17280 21422 17332
rect 10137 17255 10195 17261
rect 10137 17221 10149 17255
rect 10183 17221 10195 17255
rect 10137 17215 10195 17221
rect 8481 17187 8539 17193
rect 8481 17184 8493 17187
rect 7616 17156 8493 17184
rect 7616 17144 7622 17156
rect 8481 17153 8493 17156
rect 8527 17153 8539 17187
rect 8481 17147 8539 17153
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 10042 17144 10048 17196
rect 10100 17184 10106 17196
rect 10152 17184 10180 17215
rect 11146 17212 11152 17264
rect 11204 17252 11210 17264
rect 12342 17252 12348 17264
rect 11204 17224 12348 17252
rect 11204 17212 11210 17224
rect 12342 17212 12348 17224
rect 12400 17212 12406 17264
rect 20717 17255 20775 17261
rect 20717 17221 20729 17255
rect 20763 17252 20775 17255
rect 21634 17252 21640 17264
rect 20763 17224 21640 17252
rect 20763 17221 20775 17224
rect 20717 17215 20775 17221
rect 21634 17212 21640 17224
rect 21692 17212 21698 17264
rect 10594 17184 10600 17196
rect 10100 17156 10600 17184
rect 10100 17144 10106 17156
rect 10594 17144 10600 17156
rect 10652 17144 10658 17196
rect 11790 17144 11796 17196
rect 11848 17184 11854 17196
rect 12434 17184 12440 17196
rect 11848 17156 12440 17184
rect 11848 17144 11854 17156
rect 12434 17144 12440 17156
rect 12492 17144 12498 17196
rect 13446 17144 13452 17196
rect 13504 17184 13510 17196
rect 13504 17156 14044 17184
rect 13504 17144 13510 17156
rect 2222 17116 2228 17128
rect 2183 17088 2228 17116
rect 2222 17076 2228 17088
rect 2280 17076 2286 17128
rect 2685 17119 2743 17125
rect 2685 17085 2697 17119
rect 2731 17116 2743 17119
rect 5537 17119 5595 17125
rect 2731 17088 3188 17116
rect 2731 17085 2743 17088
rect 2685 17079 2743 17085
rect 3160 17060 3188 17088
rect 5537 17085 5549 17119
rect 5583 17116 5595 17119
rect 5626 17116 5632 17128
rect 5583 17088 5632 17116
rect 5583 17085 5595 17088
rect 5537 17079 5595 17085
rect 5626 17076 5632 17088
rect 5684 17116 5690 17128
rect 6546 17116 6552 17128
rect 5684 17088 6552 17116
rect 5684 17076 5690 17088
rect 6546 17076 6552 17088
rect 6604 17076 6610 17128
rect 8297 17119 8355 17125
rect 8297 17085 8309 17119
rect 8343 17116 8355 17119
rect 8570 17116 8576 17128
rect 8343 17088 8576 17116
rect 8343 17085 8355 17088
rect 8297 17079 8355 17085
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 8846 17076 8852 17128
rect 8904 17116 8910 17128
rect 9013 17119 9071 17125
rect 9013 17116 9025 17119
rect 8904 17088 9025 17116
rect 8904 17076 8910 17088
rect 9013 17085 9025 17088
rect 9059 17116 9071 17119
rect 9582 17116 9588 17128
rect 9059 17088 9588 17116
rect 9059 17085 9071 17088
rect 9013 17079 9071 17085
rect 9582 17076 9588 17088
rect 9640 17076 9646 17128
rect 10873 17119 10931 17125
rect 10873 17085 10885 17119
rect 10919 17116 10931 17119
rect 10962 17116 10968 17128
rect 10919 17088 10968 17116
rect 10919 17085 10931 17088
rect 10873 17079 10931 17085
rect 10962 17076 10968 17088
rect 11020 17076 11026 17128
rect 11698 17076 11704 17128
rect 11756 17076 11762 17128
rect 12452 17116 12480 17144
rect 13906 17116 13912 17128
rect 12452 17088 13912 17116
rect 13906 17076 13912 17088
rect 13964 17076 13970 17128
rect 14016 17116 14044 17156
rect 20898 17144 20904 17196
rect 20956 17184 20962 17196
rect 21085 17187 21143 17193
rect 21085 17184 21097 17187
rect 20956 17156 21097 17184
rect 20956 17144 20962 17156
rect 21085 17153 21097 17156
rect 21131 17153 21143 17187
rect 21542 17184 21548 17196
rect 21503 17156 21548 17184
rect 21085 17147 21143 17153
rect 21542 17144 21548 17156
rect 21600 17144 21606 17196
rect 14165 17119 14223 17125
rect 14165 17116 14177 17119
rect 14016 17088 14177 17116
rect 14165 17085 14177 17088
rect 14211 17085 14223 17119
rect 14165 17079 14223 17085
rect 15381 17119 15439 17125
rect 15381 17085 15393 17119
rect 15427 17116 15439 17119
rect 17402 17116 17408 17128
rect 15427 17088 17408 17116
rect 15427 17085 15439 17088
rect 15381 17079 15439 17085
rect 17402 17076 17408 17088
rect 17460 17076 17466 17128
rect 19886 17076 19892 17128
rect 19944 17116 19950 17128
rect 20533 17119 20591 17125
rect 20533 17116 20545 17119
rect 19944 17088 20545 17116
rect 19944 17076 19950 17088
rect 20533 17085 20545 17088
rect 20579 17085 20591 17119
rect 20806 17116 20812 17128
rect 20767 17088 20812 17116
rect 20533 17079 20591 17085
rect 20806 17076 20812 17088
rect 20864 17076 20870 17128
rect 2930 17051 2988 17057
rect 2930 17048 2942 17051
rect 1820 17020 2942 17048
rect 1820 17008 1826 17020
rect 2930 17017 2942 17020
rect 2976 17017 2988 17051
rect 2930 17011 2988 17017
rect 3142 17008 3148 17060
rect 3200 17008 3206 17060
rect 4430 17008 4436 17060
rect 4488 17048 4494 17060
rect 4525 17051 4583 17057
rect 4525 17048 4537 17051
rect 4488 17020 4537 17048
rect 4488 17008 4494 17020
rect 4525 17017 4537 17020
rect 4571 17048 4583 17051
rect 4985 17051 5043 17057
rect 4985 17048 4997 17051
rect 4571 17020 4997 17048
rect 4571 17017 4583 17020
rect 4525 17011 4583 17017
rect 4985 17017 4997 17020
rect 5031 17017 5043 17051
rect 4985 17011 5043 17017
rect 5166 17008 5172 17060
rect 5224 17048 5230 17060
rect 6724 17051 6782 17057
rect 5224 17020 6224 17048
rect 5224 17008 5230 17020
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 5644 16989 5672 17020
rect 5629 16983 5687 16989
rect 5629 16949 5641 16983
rect 5675 16949 5687 16983
rect 5629 16943 5687 16949
rect 5718 16940 5724 16992
rect 5776 16980 5782 16992
rect 5997 16983 6055 16989
rect 5997 16980 6009 16983
rect 5776 16952 6009 16980
rect 5776 16940 5782 16952
rect 5997 16949 6009 16952
rect 6043 16949 6055 16983
rect 6196 16980 6224 17020
rect 6724 17017 6736 17051
rect 6770 17048 6782 17051
rect 6914 17048 6920 17060
rect 6770 17020 6920 17048
rect 6770 17017 6782 17020
rect 6724 17011 6782 17017
rect 6914 17008 6920 17020
rect 6972 17008 6978 17060
rect 11606 17048 11612 17060
rect 7024 17020 11612 17048
rect 7024 16980 7052 17020
rect 11606 17008 11612 17020
rect 11664 17008 11670 17060
rect 11716 17048 11744 17076
rect 11882 17048 11888 17060
rect 11716 17020 11888 17048
rect 11882 17008 11888 17020
rect 11940 17008 11946 17060
rect 12704 17051 12762 17057
rect 12704 17017 12716 17051
rect 12750 17048 12762 17051
rect 13262 17048 13268 17060
rect 12750 17020 13268 17048
rect 12750 17017 12762 17020
rect 12704 17011 12762 17017
rect 13262 17008 13268 17020
rect 13320 17008 13326 17060
rect 13814 17008 13820 17060
rect 13872 17048 13878 17060
rect 15648 17051 15706 17057
rect 13872 17020 15424 17048
rect 13872 17008 13878 17020
rect 6196 16952 7052 16980
rect 8389 16983 8447 16989
rect 5997 16943 6055 16949
rect 8389 16949 8401 16983
rect 8435 16980 8447 16983
rect 8938 16980 8944 16992
rect 8435 16952 8944 16980
rect 8435 16949 8447 16952
rect 8389 16943 8447 16949
rect 8938 16940 8944 16952
rect 8996 16940 9002 16992
rect 9214 16940 9220 16992
rect 9272 16980 9278 16992
rect 9398 16980 9404 16992
rect 9272 16952 9404 16980
rect 9272 16940 9278 16952
rect 9398 16940 9404 16952
rect 9456 16940 9462 16992
rect 10413 16983 10471 16989
rect 10413 16949 10425 16983
rect 10459 16980 10471 16983
rect 10594 16980 10600 16992
rect 10459 16952 10600 16980
rect 10459 16949 10471 16952
rect 10413 16943 10471 16949
rect 10594 16940 10600 16952
rect 10652 16980 10658 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 10652 16952 10793 16980
rect 10652 16940 10658 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 10781 16943 10839 16949
rect 10962 16940 10968 16992
rect 11020 16980 11026 16992
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 11020 16952 11713 16980
rect 11020 16940 11026 16952
rect 11701 16949 11713 16952
rect 11747 16949 11759 16983
rect 15286 16980 15292 16992
rect 15247 16952 15292 16980
rect 11701 16943 11759 16949
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 15396 16980 15424 17020
rect 15648 17017 15660 17051
rect 15694 17048 15706 17051
rect 15746 17048 15752 17060
rect 15694 17020 15752 17048
rect 15694 17017 15706 17020
rect 15648 17011 15706 17017
rect 15746 17008 15752 17020
rect 15804 17008 15810 17060
rect 21358 17048 21364 17060
rect 21319 17020 21364 17048
rect 21358 17008 21364 17020
rect 21416 17008 21422 17060
rect 19981 16983 20039 16989
rect 19981 16980 19993 16983
rect 15396 16952 19993 16980
rect 19981 16949 19993 16952
rect 20027 16980 20039 16983
rect 20162 16980 20168 16992
rect 20027 16952 20168 16980
rect 20027 16949 20039 16952
rect 19981 16943 20039 16949
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 20349 16983 20407 16989
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 20530 16980 20536 16992
rect 20395 16952 20536 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 1762 16776 1768 16788
rect 1723 16748 1768 16776
rect 1762 16736 1768 16748
rect 1820 16736 1826 16788
rect 1946 16736 1952 16788
rect 2004 16776 2010 16788
rect 3513 16779 3571 16785
rect 3513 16776 3525 16779
rect 2004 16748 3525 16776
rect 2004 16736 2010 16748
rect 3513 16745 3525 16748
rect 3559 16745 3571 16779
rect 3513 16739 3571 16745
rect 3973 16779 4031 16785
rect 3973 16745 3985 16779
rect 4019 16776 4031 16779
rect 7282 16776 7288 16788
rect 4019 16748 7288 16776
rect 4019 16745 4031 16748
rect 3973 16739 4031 16745
rect 1581 16711 1639 16717
rect 1581 16677 1593 16711
rect 1627 16708 1639 16711
rect 3234 16708 3240 16720
rect 1627 16680 3240 16708
rect 1627 16677 1639 16680
rect 1581 16671 1639 16677
rect 3234 16668 3240 16680
rect 3292 16668 3298 16720
rect 2314 16600 2320 16652
rect 2372 16640 2378 16652
rect 2878 16643 2936 16649
rect 2878 16640 2890 16643
rect 2372 16612 2890 16640
rect 2372 16600 2378 16612
rect 2878 16609 2890 16612
rect 2924 16609 2936 16643
rect 3418 16640 3424 16652
rect 3379 16612 3424 16640
rect 2878 16603 2936 16609
rect 3418 16600 3424 16612
rect 3476 16600 3482 16652
rect 3697 16643 3755 16649
rect 3697 16609 3709 16643
rect 3743 16640 3755 16643
rect 3988 16640 4016 16739
rect 7282 16736 7288 16748
rect 7340 16736 7346 16788
rect 7377 16779 7435 16785
rect 7377 16745 7389 16779
rect 7423 16776 7435 16779
rect 7558 16776 7564 16788
rect 7423 16748 7564 16776
rect 7423 16745 7435 16748
rect 7377 16739 7435 16745
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 8628 16748 9137 16776
rect 8628 16736 8634 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9125 16739 9183 16745
rect 9769 16779 9827 16785
rect 9769 16745 9781 16779
rect 9815 16776 9827 16779
rect 10229 16779 10287 16785
rect 10229 16776 10241 16779
rect 9815 16748 10241 16776
rect 9815 16745 9827 16748
rect 9769 16739 9827 16745
rect 10229 16745 10241 16748
rect 10275 16776 10287 16779
rect 10502 16776 10508 16788
rect 10275 16748 10508 16776
rect 10275 16745 10287 16748
rect 10229 16739 10287 16745
rect 10502 16736 10508 16748
rect 10560 16736 10566 16788
rect 10597 16779 10655 16785
rect 10597 16745 10609 16779
rect 10643 16776 10655 16779
rect 10778 16776 10784 16788
rect 10643 16748 10784 16776
rect 10643 16745 10655 16748
rect 10597 16739 10655 16745
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 10962 16736 10968 16788
rect 11020 16776 11026 16788
rect 11149 16779 11207 16785
rect 11149 16776 11161 16779
rect 11020 16748 11161 16776
rect 11020 16736 11026 16748
rect 11149 16745 11161 16748
rect 11195 16745 11207 16779
rect 11149 16739 11207 16745
rect 11606 16736 11612 16788
rect 11664 16776 11670 16788
rect 11793 16779 11851 16785
rect 11793 16776 11805 16779
rect 11664 16748 11805 16776
rect 11664 16736 11670 16748
rect 11793 16745 11805 16748
rect 11839 16745 11851 16779
rect 11793 16739 11851 16745
rect 12253 16779 12311 16785
rect 12253 16745 12265 16779
rect 12299 16776 12311 16779
rect 12621 16779 12679 16785
rect 12621 16776 12633 16779
rect 12299 16748 12633 16776
rect 12299 16745 12311 16748
rect 12253 16739 12311 16745
rect 12621 16745 12633 16748
rect 12667 16745 12679 16779
rect 12621 16739 12679 16745
rect 13081 16779 13139 16785
rect 13081 16745 13093 16779
rect 13127 16776 13139 16779
rect 13633 16779 13691 16785
rect 13633 16776 13645 16779
rect 13127 16748 13645 16776
rect 13127 16745 13139 16748
rect 13081 16739 13139 16745
rect 13633 16745 13645 16748
rect 13679 16745 13691 16779
rect 15746 16776 15752 16788
rect 15707 16748 15752 16776
rect 13633 16739 13691 16745
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 16025 16779 16083 16785
rect 16025 16745 16037 16779
rect 16071 16745 16083 16779
rect 16025 16739 16083 16745
rect 20165 16779 20223 16785
rect 20165 16745 20177 16779
rect 20211 16776 20223 16779
rect 20806 16776 20812 16788
rect 20211 16748 20812 16776
rect 20211 16745 20223 16748
rect 20165 16739 20223 16745
rect 4338 16717 4344 16720
rect 4332 16708 4344 16717
rect 4299 16680 4344 16708
rect 4332 16671 4344 16680
rect 4338 16668 4344 16671
rect 4396 16668 4402 16720
rect 5552 16680 5948 16708
rect 5552 16649 5580 16680
rect 5537 16643 5595 16649
rect 5537 16640 5549 16643
rect 3743 16612 4016 16640
rect 4080 16612 5549 16640
rect 3743 16609 3755 16612
rect 3697 16603 3755 16609
rect 3142 16572 3148 16584
rect 3055 16544 3148 16572
rect 3142 16532 3148 16544
rect 3200 16572 3206 16584
rect 4080 16581 4108 16612
rect 5537 16609 5549 16612
rect 5583 16609 5595 16643
rect 5537 16603 5595 16609
rect 5626 16600 5632 16652
rect 5684 16640 5690 16652
rect 5793 16643 5851 16649
rect 5793 16640 5805 16643
rect 5684 16612 5805 16640
rect 5684 16600 5690 16612
rect 5793 16609 5805 16612
rect 5839 16609 5851 16643
rect 5920 16640 5948 16680
rect 5994 16668 6000 16720
rect 6052 16708 6058 16720
rect 6052 16680 6316 16708
rect 6052 16668 6058 16680
rect 6288 16652 6316 16680
rect 8386 16668 8392 16720
rect 8444 16708 8450 16720
rect 8490 16711 8548 16717
rect 8490 16708 8502 16711
rect 8444 16680 8502 16708
rect 8444 16668 8450 16680
rect 8490 16677 8502 16680
rect 8536 16677 8548 16711
rect 8490 16671 8548 16677
rect 8588 16680 9536 16708
rect 6178 16640 6184 16652
rect 5920 16612 6184 16640
rect 5793 16603 5851 16609
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 6270 16600 6276 16652
rect 6328 16640 6334 16652
rect 8588 16640 8616 16680
rect 6328 16612 8616 16640
rect 9508 16640 9536 16680
rect 9582 16668 9588 16720
rect 9640 16708 9646 16720
rect 10410 16708 10416 16720
rect 9640 16680 10416 16708
rect 9640 16668 9646 16680
rect 10410 16668 10416 16680
rect 10468 16668 10474 16720
rect 11057 16711 11115 16717
rect 11057 16677 11069 16711
rect 11103 16708 11115 16711
rect 11698 16708 11704 16720
rect 11103 16680 11704 16708
rect 11103 16677 11115 16680
rect 11057 16671 11115 16677
rect 11698 16668 11704 16680
rect 11756 16668 11762 16720
rect 14636 16711 14694 16717
rect 14636 16677 14648 16711
rect 14682 16708 14694 16711
rect 15286 16708 15292 16720
rect 14682 16680 15292 16708
rect 14682 16677 14694 16680
rect 14636 16671 14694 16677
rect 15286 16668 15292 16680
rect 15344 16668 15350 16720
rect 9858 16640 9864 16652
rect 9508 16612 9864 16640
rect 6328 16600 6334 16612
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 10318 16600 10324 16652
rect 10376 16640 10382 16652
rect 10376 16612 10548 16640
rect 10376 16600 10382 16612
rect 4065 16575 4123 16581
rect 4065 16572 4077 16575
rect 3200 16544 4077 16572
rect 3200 16532 3206 16544
rect 3712 16516 3740 16544
rect 4065 16541 4077 16544
rect 4111 16541 4123 16575
rect 4065 16535 4123 16541
rect 8757 16575 8815 16581
rect 8757 16541 8769 16575
rect 8803 16572 8815 16575
rect 9030 16572 9036 16584
rect 8803 16544 9036 16572
rect 8803 16541 8815 16544
rect 8757 16535 8815 16541
rect 9030 16532 9036 16544
rect 9088 16532 9094 16584
rect 10042 16572 10048 16584
rect 10003 16544 10048 16572
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 10137 16575 10195 16581
rect 10137 16541 10149 16575
rect 10183 16572 10195 16575
rect 10410 16572 10416 16584
rect 10183 16544 10416 16572
rect 10183 16541 10195 16544
rect 10137 16535 10195 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 10520 16572 10548 16612
rect 11146 16600 11152 16652
rect 11204 16640 11210 16652
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 11204 16612 11897 16640
rect 11204 16600 11210 16612
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 12526 16640 12532 16652
rect 11885 16603 11943 16609
rect 12360 16612 12532 16640
rect 10520 16544 10732 16572
rect 3237 16507 3295 16513
rect 3237 16473 3249 16507
rect 3283 16504 3295 16507
rect 3510 16504 3516 16516
rect 3283 16476 3516 16504
rect 3283 16473 3295 16476
rect 3237 16467 3295 16473
rect 3510 16464 3516 16476
rect 3568 16464 3574 16516
rect 3694 16464 3700 16516
rect 3752 16464 3758 16516
rect 8938 16504 8944 16516
rect 8899 16476 8944 16504
rect 8938 16464 8944 16476
rect 8996 16464 9002 16516
rect 10704 16513 10732 16544
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 11241 16575 11299 16581
rect 11241 16572 11253 16575
rect 11112 16544 11253 16572
rect 11112 16532 11118 16544
rect 11241 16541 11253 16544
rect 11287 16541 11299 16575
rect 11241 16535 11299 16541
rect 11701 16575 11759 16581
rect 11701 16541 11713 16575
rect 11747 16572 11759 16575
rect 12360 16572 12388 16612
rect 12526 16600 12532 16612
rect 12584 16600 12590 16652
rect 12710 16640 12716 16652
rect 12671 16612 12716 16640
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 13078 16600 13084 16652
rect 13136 16640 13142 16652
rect 13541 16643 13599 16649
rect 13136 16612 13216 16640
rect 13136 16600 13142 16612
rect 11747 16544 12388 16572
rect 11747 16541 11759 16544
rect 11701 16535 11759 16541
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 12492 16544 12537 16572
rect 12492 16532 12498 16544
rect 13188 16513 13216 16612
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 13814 16640 13820 16652
rect 13587 16612 13820 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 13906 16600 13912 16652
rect 13964 16640 13970 16652
rect 14369 16643 14427 16649
rect 14369 16640 14381 16643
rect 13964 16612 14381 16640
rect 13964 16600 13970 16612
rect 14369 16609 14381 16612
rect 14415 16609 14427 16643
rect 16040 16640 16068 16739
rect 20806 16736 20812 16748
rect 20864 16736 20870 16788
rect 20993 16779 21051 16785
rect 20993 16745 21005 16779
rect 21039 16745 21051 16779
rect 20993 16739 21051 16745
rect 16758 16668 16764 16720
rect 16816 16708 16822 16720
rect 17138 16711 17196 16717
rect 17138 16708 17150 16711
rect 16816 16680 17150 16708
rect 16816 16668 16822 16680
rect 17138 16677 17150 16680
rect 17184 16677 17196 16711
rect 17138 16671 17196 16677
rect 19886 16668 19892 16720
rect 19944 16708 19950 16720
rect 20349 16711 20407 16717
rect 20349 16708 20361 16711
rect 19944 16680 20361 16708
rect 19944 16668 19950 16680
rect 20349 16677 20361 16680
rect 20395 16708 20407 16711
rect 21008 16708 21036 16739
rect 21361 16711 21419 16717
rect 21361 16708 21373 16711
rect 20395 16680 20576 16708
rect 21008 16680 21373 16708
rect 20395 16677 20407 16680
rect 20349 16671 20407 16677
rect 17402 16640 17408 16652
rect 14369 16603 14427 16609
rect 14476 16612 16068 16640
rect 17363 16612 17408 16640
rect 13262 16532 13268 16584
rect 13320 16572 13326 16584
rect 13725 16575 13783 16581
rect 13725 16572 13737 16575
rect 13320 16544 13737 16572
rect 13320 16532 13326 16544
rect 13725 16541 13737 16544
rect 13771 16541 13783 16575
rect 13725 16535 13783 16541
rect 14274 16532 14280 16584
rect 14332 16572 14338 16584
rect 14476 16572 14504 16612
rect 17402 16600 17408 16612
rect 17460 16600 17466 16652
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 20548 16649 20576 16680
rect 21361 16677 21373 16680
rect 21407 16677 21419 16711
rect 21542 16708 21548 16720
rect 21503 16680 21548 16708
rect 21361 16671 21419 16677
rect 21542 16668 21548 16680
rect 21600 16668 21606 16720
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 19392 16612 19993 16640
rect 19392 16600 19398 16612
rect 19981 16609 19993 16612
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 20533 16643 20591 16649
rect 20533 16609 20545 16643
rect 20579 16609 20591 16643
rect 20533 16603 20591 16609
rect 20809 16643 20867 16649
rect 20809 16609 20821 16643
rect 20855 16609 20867 16643
rect 22005 16643 22063 16649
rect 22005 16640 22017 16643
rect 20809 16603 20867 16609
rect 20916 16612 22017 16640
rect 20824 16572 20852 16603
rect 14332 16544 14504 16572
rect 20640 16544 20852 16572
rect 14332 16532 14338 16544
rect 10689 16507 10747 16513
rect 10689 16473 10701 16507
rect 10735 16473 10747 16507
rect 10689 16467 10747 16473
rect 13173 16507 13231 16513
rect 13173 16473 13185 16507
rect 13219 16473 13231 16507
rect 13173 16467 13231 16473
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 2406 16396 2412 16448
rect 2464 16436 2470 16448
rect 5258 16436 5264 16448
rect 2464 16408 5264 16436
rect 2464 16396 2470 16408
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 5445 16439 5503 16445
rect 5445 16405 5457 16439
rect 5491 16436 5503 16439
rect 6178 16436 6184 16448
rect 5491 16408 6184 16436
rect 5491 16405 5503 16408
rect 5445 16399 5503 16405
rect 6178 16396 6184 16408
rect 6236 16396 6242 16448
rect 6914 16436 6920 16448
rect 6875 16408 6920 16436
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 13722 16396 13728 16448
rect 13780 16436 13786 16448
rect 14001 16439 14059 16445
rect 14001 16436 14013 16439
rect 13780 16408 14013 16436
rect 13780 16396 13786 16408
rect 14001 16405 14013 16408
rect 14047 16405 14059 16439
rect 14001 16399 14059 16405
rect 15378 16396 15384 16448
rect 15436 16436 15442 16448
rect 20640 16436 20668 16544
rect 20717 16507 20775 16513
rect 20717 16473 20729 16507
rect 20763 16504 20775 16507
rect 20916 16504 20944 16612
rect 22005 16609 22017 16612
rect 22051 16609 22063 16643
rect 22005 16603 22063 16609
rect 20763 16476 20944 16504
rect 20763 16473 20775 16476
rect 20717 16467 20775 16473
rect 21085 16439 21143 16445
rect 21085 16436 21097 16439
rect 15436 16408 21097 16436
rect 15436 16396 15442 16408
rect 21085 16405 21097 16408
rect 21131 16405 21143 16439
rect 21085 16399 21143 16405
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 2317 16235 2375 16241
rect 2317 16201 2329 16235
rect 2363 16232 2375 16235
rect 2406 16232 2412 16244
rect 2363 16204 2412 16232
rect 2363 16201 2375 16204
rect 2317 16195 2375 16201
rect 2406 16192 2412 16204
rect 2464 16192 2470 16244
rect 3234 16232 3240 16244
rect 3195 16204 3240 16232
rect 3234 16192 3240 16204
rect 3292 16192 3298 16244
rect 3326 16192 3332 16244
rect 3384 16232 3390 16244
rect 3513 16235 3571 16241
rect 3513 16232 3525 16235
rect 3384 16204 3525 16232
rect 3384 16192 3390 16204
rect 3513 16201 3525 16204
rect 3559 16201 3571 16235
rect 3513 16195 3571 16201
rect 4709 16235 4767 16241
rect 4709 16201 4721 16235
rect 4755 16232 4767 16235
rect 8941 16235 8999 16241
rect 4755 16204 8616 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 3789 16167 3847 16173
rect 3789 16164 3801 16167
rect 1872 16136 3801 16164
rect 1762 16096 1768 16108
rect 1723 16068 1768 16096
rect 1762 16056 1768 16068
rect 1820 16056 1826 16108
rect 1872 16105 1900 16136
rect 3789 16133 3801 16136
rect 3835 16133 3847 16167
rect 3789 16127 3847 16133
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16065 1915 16099
rect 1857 16059 1915 16065
rect 2314 16056 2320 16108
rect 2372 16096 2378 16108
rect 3053 16099 3111 16105
rect 3053 16096 3065 16099
rect 2372 16068 3065 16096
rect 2372 16056 2378 16068
rect 3053 16065 3065 16068
rect 3099 16096 3111 16099
rect 4341 16099 4399 16105
rect 4341 16096 4353 16099
rect 3099 16068 4353 16096
rect 3099 16065 3111 16068
rect 3053 16059 3111 16065
rect 4341 16065 4353 16068
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 3421 16031 3479 16037
rect 3421 15997 3433 16031
rect 3467 15997 3479 16031
rect 3421 15991 3479 15997
rect 3697 16031 3755 16037
rect 3697 15997 3709 16031
rect 3743 16028 3755 16031
rect 4724 16028 4752 16195
rect 7285 16167 7343 16173
rect 7285 16133 7297 16167
rect 7331 16164 7343 16167
rect 8588 16164 8616 16204
rect 8941 16201 8953 16235
rect 8987 16232 8999 16235
rect 9306 16232 9312 16244
rect 8987 16204 9312 16232
rect 8987 16201 8999 16204
rect 8941 16195 8999 16201
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 9582 16192 9588 16244
rect 9640 16232 9646 16244
rect 9677 16235 9735 16241
rect 9677 16232 9689 16235
rect 9640 16204 9689 16232
rect 9640 16192 9646 16204
rect 9677 16201 9689 16204
rect 9723 16201 9735 16235
rect 9677 16195 9735 16201
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 12250 16232 12256 16244
rect 10376 16204 12256 16232
rect 10376 16192 10382 16204
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 13262 16232 13268 16244
rect 13223 16204 13268 16232
rect 13262 16192 13268 16204
rect 13320 16192 13326 16244
rect 13538 16192 13544 16244
rect 13596 16232 13602 16244
rect 14185 16235 14243 16241
rect 14185 16232 14197 16235
rect 13596 16204 14197 16232
rect 13596 16192 13602 16204
rect 14185 16201 14197 16204
rect 14231 16201 14243 16235
rect 14185 16195 14243 16201
rect 15289 16235 15347 16241
rect 15289 16201 15301 16235
rect 15335 16232 15347 16235
rect 15562 16232 15568 16244
rect 15335 16204 15568 16232
rect 15335 16201 15347 16204
rect 15289 16195 15347 16201
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 20809 16235 20867 16241
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 21358 16232 21364 16244
rect 20855 16204 21364 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 21358 16192 21364 16204
rect 21416 16192 21422 16244
rect 9858 16164 9864 16176
rect 7331 16136 8524 16164
rect 8588 16136 9864 16164
rect 7331 16133 7343 16136
rect 7285 16127 7343 16133
rect 5353 16099 5411 16105
rect 5353 16065 5365 16099
rect 5399 16065 5411 16099
rect 5534 16096 5540 16108
rect 5495 16068 5540 16096
rect 5353 16059 5411 16065
rect 3743 16000 4752 16028
rect 5368 16028 5396 16059
rect 5534 16056 5540 16068
rect 5592 16096 5598 16108
rect 6454 16096 6460 16108
rect 5592 16068 6460 16096
rect 5592 16056 5598 16068
rect 6454 16056 6460 16068
rect 6512 16056 6518 16108
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16096 6791 16099
rect 6914 16096 6920 16108
rect 6779 16068 6920 16096
rect 6779 16065 6791 16068
rect 6733 16059 6791 16065
rect 6914 16056 6920 16068
rect 6972 16096 6978 16108
rect 7469 16099 7527 16105
rect 7469 16096 7481 16099
rect 6972 16068 7481 16096
rect 6972 16056 6978 16068
rect 7469 16065 7481 16068
rect 7515 16065 7527 16099
rect 8386 16096 8392 16108
rect 8347 16068 8392 16096
rect 7469 16059 7527 16065
rect 8386 16056 8392 16068
rect 8444 16056 8450 16108
rect 8496 16105 8524 16136
rect 9858 16124 9864 16136
rect 9916 16124 9922 16176
rect 13280 16164 13308 16192
rect 21542 16164 21548 16176
rect 13280 16136 14780 16164
rect 21503 16136 21548 16164
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 11790 16056 11796 16108
rect 11848 16096 11854 16108
rect 14752 16105 14780 16136
rect 21542 16124 21548 16136
rect 21600 16124 21606 16176
rect 11885 16099 11943 16105
rect 11885 16096 11897 16099
rect 11848 16068 11897 16096
rect 11848 16056 11854 16068
rect 11885 16065 11897 16068
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 13449 16099 13507 16105
rect 13449 16065 13461 16099
rect 13495 16065 13507 16099
rect 13449 16059 13507 16065
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 5810 16028 5816 16040
rect 5368 16000 5816 16028
rect 3743 15997 3755 16000
rect 3697 15991 3755 15997
rect 1949 15963 2007 15969
rect 1949 15929 1961 15963
rect 1995 15960 2007 15963
rect 2866 15960 2872 15972
rect 1995 15932 2452 15960
rect 2827 15932 2872 15960
rect 1995 15929 2007 15932
rect 1949 15923 2007 15929
rect 2424 15901 2452 15932
rect 2866 15920 2872 15932
rect 2924 15920 2930 15972
rect 3436 15960 3464 15991
rect 5552 15972 5580 16000
rect 5810 15988 5816 16000
rect 5868 15988 5874 16040
rect 6270 16028 6276 16040
rect 6104 16000 6276 16028
rect 3786 15960 3792 15972
rect 3436 15932 3792 15960
rect 3786 15920 3792 15932
rect 3844 15920 3850 15972
rect 4157 15963 4215 15969
rect 4157 15929 4169 15963
rect 4203 15960 4215 15963
rect 4430 15960 4436 15972
rect 4203 15932 4436 15960
rect 4203 15929 4215 15932
rect 4157 15923 4215 15929
rect 4430 15920 4436 15932
rect 4488 15920 4494 15972
rect 5534 15920 5540 15972
rect 5592 15920 5598 15972
rect 5629 15963 5687 15969
rect 5629 15929 5641 15963
rect 5675 15960 5687 15963
rect 6104 15960 6132 16000
rect 6270 15988 6276 16000
rect 6328 15988 6334 16040
rect 9950 15988 9956 16040
rect 10008 16028 10014 16040
rect 10226 16028 10232 16040
rect 10008 16000 10232 16028
rect 10008 15988 10014 16000
rect 10226 15988 10232 16000
rect 10284 15988 10290 16040
rect 11057 16031 11115 16037
rect 11057 16028 11069 16031
rect 10336 16000 11069 16028
rect 5675 15932 6132 15960
rect 6181 15963 6239 15969
rect 5675 15929 5687 15932
rect 5629 15923 5687 15929
rect 6181 15929 6193 15963
rect 6227 15960 6239 15963
rect 6638 15960 6644 15972
rect 6227 15932 6644 15960
rect 6227 15929 6239 15932
rect 6181 15923 6239 15929
rect 6638 15920 6644 15932
rect 6696 15920 6702 15972
rect 7650 15960 7656 15972
rect 7611 15932 7656 15960
rect 7650 15920 7656 15932
rect 7708 15920 7714 15972
rect 8573 15963 8631 15969
rect 8573 15960 8585 15963
rect 8128 15932 8585 15960
rect 2409 15895 2467 15901
rect 2409 15861 2421 15895
rect 2455 15861 2467 15895
rect 2409 15855 2467 15861
rect 2774 15852 2780 15904
rect 2832 15892 2838 15904
rect 4246 15892 4252 15904
rect 2832 15864 2877 15892
rect 4207 15864 4252 15892
rect 2832 15852 2838 15864
rect 4246 15852 4252 15864
rect 4304 15852 4310 15904
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5994 15892 6000 15904
rect 5955 15864 6000 15892
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 6270 15852 6276 15904
rect 6328 15892 6334 15904
rect 6825 15895 6883 15901
rect 6825 15892 6837 15895
rect 6328 15864 6837 15892
rect 6328 15852 6334 15864
rect 6825 15861 6837 15864
rect 6871 15861 6883 15895
rect 6825 15855 6883 15861
rect 6914 15852 6920 15904
rect 6972 15892 6978 15904
rect 7742 15892 7748 15904
rect 6972 15864 7017 15892
rect 7703 15864 7748 15892
rect 6972 15852 6978 15864
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 8128 15901 8156 15932
rect 8573 15929 8585 15932
rect 8619 15929 8631 15963
rect 8573 15923 8631 15929
rect 9030 15920 9036 15972
rect 9088 15960 9094 15972
rect 10336 15960 10364 16000
rect 11057 15997 11069 16000
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 12152 16031 12210 16037
rect 12152 15997 12164 16031
rect 12198 16028 12210 16031
rect 12434 16028 12440 16040
rect 12198 16000 12440 16028
rect 12198 15997 12210 16000
rect 12152 15991 12210 15997
rect 12434 15988 12440 16000
rect 12492 16028 12498 16040
rect 13170 16028 13176 16040
rect 12492 16000 13176 16028
rect 12492 15988 12498 16000
rect 13170 15988 13176 16000
rect 13228 16028 13234 16040
rect 13464 16028 13492 16059
rect 15286 16056 15292 16108
rect 15344 16096 15350 16108
rect 15841 16099 15899 16105
rect 15841 16096 15853 16099
rect 15344 16068 15853 16096
rect 15344 16056 15350 16068
rect 15841 16065 15853 16068
rect 15887 16065 15899 16099
rect 15841 16059 15899 16065
rect 13228 16000 13492 16028
rect 13633 16031 13691 16037
rect 13228 15988 13234 16000
rect 13633 15997 13645 16031
rect 13679 16028 13691 16031
rect 13722 16028 13728 16040
rect 13679 16000 13728 16028
rect 13679 15997 13691 16000
rect 13633 15991 13691 15997
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 20622 16028 20628 16040
rect 13832 16000 15700 16028
rect 20583 16000 20628 16028
rect 10778 15960 10784 15972
rect 10836 15969 10842 15972
rect 9088 15932 10364 15960
rect 10748 15932 10784 15960
rect 9088 15920 9094 15932
rect 10778 15920 10784 15932
rect 10836 15923 10848 15969
rect 13832 15960 13860 16000
rect 15672 15969 15700 16000
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 14553 15963 14611 15969
rect 14553 15960 14565 15963
rect 10879 15932 13860 15960
rect 14108 15932 14565 15960
rect 10836 15920 10842 15923
rect 8113 15895 8171 15901
rect 8113 15861 8125 15895
rect 8159 15861 8171 15895
rect 8113 15855 8171 15861
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 9490 15892 9496 15904
rect 8444 15864 9496 15892
rect 8444 15852 8450 15864
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10879 15892 10907 15932
rect 11698 15892 11704 15904
rect 9916 15864 10907 15892
rect 11659 15864 11704 15892
rect 9916 15852 9922 15864
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 13725 15895 13783 15901
rect 13725 15861 13737 15895
rect 13771 15892 13783 15895
rect 13906 15892 13912 15904
rect 13771 15864 13912 15892
rect 13771 15861 13783 15864
rect 13725 15855 13783 15861
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 14108 15901 14136 15932
rect 14553 15929 14565 15932
rect 14599 15929 14611 15963
rect 14553 15923 14611 15929
rect 15657 15963 15715 15969
rect 15657 15929 15669 15963
rect 15703 15960 15715 15963
rect 15703 15932 16344 15960
rect 15703 15929 15715 15932
rect 15657 15923 15715 15929
rect 16316 15904 16344 15932
rect 20714 15920 20720 15972
rect 20772 15960 20778 15972
rect 20993 15963 21051 15969
rect 20993 15960 21005 15963
rect 20772 15932 21005 15960
rect 20772 15920 20778 15932
rect 20993 15929 21005 15932
rect 21039 15929 21051 15963
rect 21174 15960 21180 15972
rect 21135 15932 21180 15960
rect 20993 15923 21051 15929
rect 21174 15920 21180 15932
rect 21232 15920 21238 15972
rect 21361 15963 21419 15969
rect 21361 15929 21373 15963
rect 21407 15929 21419 15963
rect 21361 15923 21419 15929
rect 14093 15895 14151 15901
rect 14093 15861 14105 15895
rect 14139 15861 14151 15895
rect 14093 15855 14151 15861
rect 14274 15852 14280 15904
rect 14332 15892 14338 15904
rect 14645 15895 14703 15901
rect 14645 15892 14657 15895
rect 14332 15864 14657 15892
rect 14332 15852 14338 15864
rect 14645 15861 14657 15864
rect 14691 15861 14703 15895
rect 14645 15855 14703 15861
rect 15749 15895 15807 15901
rect 15749 15861 15761 15895
rect 15795 15892 15807 15895
rect 15838 15892 15844 15904
rect 15795 15864 15844 15892
rect 15795 15861 15807 15864
rect 15749 15855 15807 15861
rect 15838 15852 15844 15864
rect 15896 15852 15902 15904
rect 16114 15892 16120 15904
rect 16075 15864 16120 15892
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 16298 15852 16304 15904
rect 16356 15892 16362 15904
rect 16393 15895 16451 15901
rect 16393 15892 16405 15895
rect 16356 15864 16405 15892
rect 16356 15852 16362 15864
rect 16393 15861 16405 15864
rect 16439 15861 16451 15895
rect 16393 15855 16451 15861
rect 20898 15852 20904 15904
rect 20956 15892 20962 15904
rect 21376 15892 21404 15923
rect 20956 15864 21404 15892
rect 20956 15852 20962 15864
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1854 15688 1860 15700
rect 1815 15660 1860 15688
rect 1854 15648 1860 15660
rect 1912 15648 1918 15700
rect 2314 15688 2320 15700
rect 2275 15660 2320 15688
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 3418 15648 3424 15700
rect 3476 15688 3482 15700
rect 3881 15691 3939 15697
rect 3881 15688 3893 15691
rect 3476 15660 3893 15688
rect 3476 15648 3482 15660
rect 3881 15657 3893 15660
rect 3927 15657 3939 15691
rect 4430 15688 4436 15700
rect 4391 15660 4436 15688
rect 3881 15651 3939 15657
rect 4430 15648 4436 15660
rect 4488 15648 4494 15700
rect 5629 15691 5687 15697
rect 5629 15657 5641 15691
rect 5675 15688 5687 15691
rect 5994 15688 6000 15700
rect 5675 15660 6000 15688
rect 5675 15657 5687 15660
rect 5629 15651 5687 15657
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 6454 15688 6460 15700
rect 6415 15660 6460 15688
rect 6454 15648 6460 15660
rect 6512 15648 6518 15700
rect 7653 15691 7711 15697
rect 7653 15657 7665 15691
rect 7699 15688 7711 15691
rect 7742 15688 7748 15700
rect 7699 15660 7748 15688
rect 7699 15657 7711 15660
rect 7653 15651 7711 15657
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 8938 15648 8944 15700
rect 8996 15688 9002 15700
rect 11146 15688 11152 15700
rect 8996 15660 11152 15688
rect 8996 15648 9002 15660
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 11238 15648 11244 15700
rect 11296 15688 11302 15700
rect 11333 15691 11391 15697
rect 11333 15688 11345 15691
rect 11296 15660 11345 15688
rect 11296 15648 11302 15660
rect 11333 15657 11345 15660
rect 11379 15657 11391 15691
rect 11333 15651 11391 15657
rect 11882 15648 11888 15700
rect 11940 15688 11946 15700
rect 12621 15691 12679 15697
rect 12621 15688 12633 15691
rect 11940 15660 12633 15688
rect 11940 15648 11946 15660
rect 12621 15657 12633 15660
rect 12667 15657 12679 15691
rect 12621 15651 12679 15657
rect 12710 15648 12716 15700
rect 12768 15688 12774 15700
rect 12989 15691 13047 15697
rect 12989 15688 13001 15691
rect 12768 15660 13001 15688
rect 12768 15648 12774 15660
rect 12989 15657 13001 15660
rect 13035 15657 13047 15691
rect 13906 15688 13912 15700
rect 13867 15660 13912 15688
rect 12989 15651 13047 15657
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 14366 15648 14372 15700
rect 14424 15688 14430 15700
rect 14921 15691 14979 15697
rect 14921 15688 14933 15691
rect 14424 15660 14933 15688
rect 14424 15648 14430 15660
rect 14921 15657 14933 15660
rect 14967 15657 14979 15691
rect 14921 15651 14979 15657
rect 15749 15691 15807 15697
rect 15749 15657 15761 15691
rect 15795 15688 15807 15691
rect 16114 15688 16120 15700
rect 15795 15660 16120 15688
rect 15795 15657 15807 15660
rect 15749 15651 15807 15657
rect 16114 15648 16120 15660
rect 16172 15648 16178 15700
rect 19886 15688 19892 15700
rect 16592 15660 19892 15688
rect 3234 15580 3240 15632
rect 3292 15580 3298 15632
rect 4893 15623 4951 15629
rect 4893 15589 4905 15623
rect 4939 15620 4951 15623
rect 5166 15620 5172 15632
rect 4939 15592 5172 15620
rect 4939 15589 4951 15592
rect 4893 15583 4951 15589
rect 5166 15580 5172 15592
rect 5224 15580 5230 15632
rect 5537 15623 5595 15629
rect 5537 15589 5549 15623
rect 5583 15620 5595 15623
rect 5718 15620 5724 15632
rect 5583 15592 5724 15620
rect 5583 15589 5595 15592
rect 5537 15583 5595 15589
rect 5718 15580 5724 15592
rect 5776 15580 5782 15632
rect 6365 15623 6423 15629
rect 6365 15589 6377 15623
rect 6411 15620 6423 15623
rect 6546 15620 6552 15632
rect 6411 15592 6552 15620
rect 6411 15589 6423 15592
rect 6365 15583 6423 15589
rect 6546 15580 6552 15592
rect 6604 15580 6610 15632
rect 8956 15620 8984 15648
rect 7208 15592 8984 15620
rect 9392 15623 9450 15629
rect 1578 15552 1584 15564
rect 1539 15524 1584 15552
rect 1578 15512 1584 15524
rect 1636 15512 1642 15564
rect 1946 15552 1952 15564
rect 1907 15524 1952 15552
rect 1946 15512 1952 15524
rect 2004 15512 2010 15564
rect 3252 15552 3280 15580
rect 3430 15555 3488 15561
rect 3430 15552 3442 15555
rect 3252 15524 3442 15552
rect 3430 15521 3442 15524
rect 3476 15521 3488 15555
rect 3430 15515 3488 15521
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4706 15552 4712 15564
rect 4111 15524 4712 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 5902 15552 5908 15564
rect 4847 15524 5908 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 5902 15512 5908 15524
rect 5960 15512 5966 15564
rect 7208 15552 7236 15592
rect 9392 15589 9404 15623
rect 9438 15620 9450 15623
rect 9490 15620 9496 15632
rect 9438 15592 9496 15620
rect 9438 15589 9450 15592
rect 9392 15583 9450 15589
rect 9490 15580 9496 15592
rect 9548 15580 9554 15632
rect 15286 15620 15292 15632
rect 9600 15592 14504 15620
rect 6012 15524 7236 15552
rect 7285 15555 7343 15561
rect 3694 15484 3700 15496
rect 3607 15456 3700 15484
rect 3694 15444 3700 15456
rect 3752 15484 3758 15496
rect 4154 15484 4160 15496
rect 3752 15456 4160 15484
rect 3752 15444 3758 15456
rect 4154 15444 4160 15456
rect 4212 15444 4218 15496
rect 4982 15484 4988 15496
rect 4943 15456 4988 15484
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 5445 15487 5503 15493
rect 5445 15453 5457 15487
rect 5491 15484 5503 15487
rect 5626 15484 5632 15496
rect 5491 15456 5632 15484
rect 5491 15453 5503 15456
rect 5445 15447 5503 15453
rect 5626 15444 5632 15456
rect 5684 15444 5690 15496
rect 6012 15484 6040 15524
rect 7285 15521 7297 15555
rect 7331 15552 7343 15555
rect 7745 15555 7803 15561
rect 7745 15552 7757 15555
rect 7331 15524 7757 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 7745 15521 7757 15524
rect 7791 15521 7803 15555
rect 7745 15515 7803 15521
rect 8570 15512 8576 15564
rect 8628 15552 8634 15564
rect 9030 15552 9036 15564
rect 8628 15524 9036 15552
rect 8628 15512 8634 15524
rect 9030 15512 9036 15524
rect 9088 15552 9094 15564
rect 9125 15555 9183 15561
rect 9125 15552 9137 15555
rect 9088 15524 9137 15552
rect 9088 15512 9094 15524
rect 9125 15521 9137 15524
rect 9171 15521 9183 15555
rect 9600 15552 9628 15592
rect 9125 15515 9183 15521
rect 9232 15524 9628 15552
rect 6178 15484 6184 15496
rect 5920 15456 6040 15484
rect 6139 15456 6184 15484
rect 1394 15416 1400 15428
rect 1355 15388 1400 15416
rect 1394 15376 1400 15388
rect 1452 15376 1458 15428
rect 3786 15376 3792 15428
rect 3844 15416 3850 15428
rect 4249 15419 4307 15425
rect 4249 15416 4261 15419
rect 3844 15388 4261 15416
rect 3844 15376 3850 15388
rect 4249 15385 4261 15388
rect 4295 15416 4307 15419
rect 5920 15416 5948 15456
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 6730 15444 6736 15496
rect 6788 15484 6794 15496
rect 7009 15487 7067 15493
rect 7009 15484 7021 15487
rect 6788 15456 7021 15484
rect 6788 15444 6794 15456
rect 7009 15453 7021 15456
rect 7055 15453 7067 15487
rect 7190 15484 7196 15496
rect 7103 15456 7196 15484
rect 7009 15447 7067 15453
rect 7190 15444 7196 15456
rect 7248 15484 7254 15496
rect 9232 15484 9260 15524
rect 10226 15512 10232 15564
rect 10284 15552 10290 15564
rect 10965 15555 11023 15561
rect 10965 15552 10977 15555
rect 10284 15524 10977 15552
rect 10284 15512 10290 15524
rect 10965 15521 10977 15524
rect 11011 15521 11023 15555
rect 10965 15515 11023 15521
rect 11146 15512 11152 15564
rect 11204 15552 11210 15564
rect 12529 15555 12587 15561
rect 12529 15552 12541 15555
rect 11204 15524 12541 15552
rect 11204 15512 11210 15524
rect 12529 15521 12541 15524
rect 12575 15552 12587 15555
rect 13262 15552 13268 15564
rect 12575 15524 13268 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 13446 15552 13452 15564
rect 13359 15524 13452 15552
rect 13446 15512 13452 15524
rect 13504 15552 13510 15564
rect 14090 15552 14096 15564
rect 13504 15524 14096 15552
rect 13504 15512 13510 15524
rect 14090 15512 14096 15524
rect 14148 15512 14154 15564
rect 10778 15484 10784 15496
rect 7248 15456 9260 15484
rect 10520 15456 10784 15484
rect 7248 15444 7254 15456
rect 4295 15388 5948 15416
rect 5997 15419 6055 15425
rect 4295 15385 4307 15388
rect 4249 15379 4307 15385
rect 5997 15385 6009 15419
rect 6043 15416 6055 15419
rect 6270 15416 6276 15428
rect 6043 15388 6276 15416
rect 6043 15385 6055 15388
rect 5997 15379 6055 15385
rect 6270 15376 6276 15388
rect 6328 15376 6334 15428
rect 10520 15425 10548 15456
rect 10778 15444 10784 15456
rect 10836 15444 10842 15496
rect 10870 15444 10876 15496
rect 10928 15484 10934 15496
rect 11974 15484 11980 15496
rect 10928 15456 10973 15484
rect 11935 15456 11980 15484
rect 10928 15444 10934 15456
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 12434 15444 12440 15496
rect 12492 15484 12498 15496
rect 12894 15484 12900 15496
rect 12492 15456 12537 15484
rect 12728 15456 12900 15484
rect 12492 15444 12498 15456
rect 10505 15419 10563 15425
rect 6380 15388 8340 15416
rect 2038 15308 2044 15360
rect 2096 15348 2102 15360
rect 2133 15351 2191 15357
rect 2133 15348 2145 15351
rect 2096 15320 2145 15348
rect 2096 15308 2102 15320
rect 2133 15317 2145 15320
rect 2179 15317 2191 15351
rect 2133 15311 2191 15317
rect 5166 15308 5172 15360
rect 5224 15348 5230 15360
rect 5442 15348 5448 15360
rect 5224 15320 5448 15348
rect 5224 15308 5230 15320
rect 5442 15308 5448 15320
rect 5500 15348 5506 15360
rect 6380 15348 6408 15388
rect 5500 15320 6408 15348
rect 6825 15351 6883 15357
rect 5500 15308 5506 15320
rect 6825 15317 6837 15351
rect 6871 15348 6883 15351
rect 8202 15348 8208 15360
rect 6871 15320 8208 15348
rect 6871 15317 6883 15320
rect 6825 15311 6883 15317
rect 8202 15308 8208 15320
rect 8260 15308 8266 15360
rect 8312 15348 8340 15388
rect 10505 15385 10517 15419
rect 10551 15385 10563 15419
rect 12728 15416 12756 15456
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 13170 15484 13176 15496
rect 13131 15456 13176 15484
rect 13170 15444 13176 15456
rect 13228 15444 13234 15496
rect 13357 15487 13415 15493
rect 13357 15484 13369 15487
rect 13280 15456 13369 15484
rect 10505 15379 10563 15385
rect 10612 15388 12756 15416
rect 10612 15348 10640 15388
rect 8312 15320 10640 15348
rect 11793 15351 11851 15357
rect 11793 15317 11805 15351
rect 11839 15348 11851 15351
rect 11882 15348 11888 15360
rect 11839 15320 11888 15348
rect 11839 15317 11851 15320
rect 11793 15311 11851 15317
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 12069 15351 12127 15357
rect 12069 15348 12081 15351
rect 12032 15320 12081 15348
rect 12032 15308 12038 15320
rect 12069 15317 12081 15320
rect 12115 15348 12127 15351
rect 13280 15348 13308 15456
rect 13357 15453 13369 15456
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 13817 15419 13875 15425
rect 13817 15385 13829 15419
rect 13863 15416 13875 15419
rect 14274 15416 14280 15428
rect 13863 15388 14280 15416
rect 13863 15385 13875 15388
rect 13817 15379 13875 15385
rect 14274 15376 14280 15388
rect 14332 15376 14338 15428
rect 14476 15416 14504 15592
rect 14844 15592 15292 15620
rect 14844 15552 14872 15592
rect 15286 15580 15292 15592
rect 15344 15580 15350 15632
rect 14752 15524 14872 15552
rect 14752 15493 14780 15524
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 14826 15444 14832 15496
rect 14884 15484 14890 15496
rect 15304 15484 15332 15580
rect 15378 15512 15384 15564
rect 15436 15552 15442 15564
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 15436 15524 15669 15552
rect 15436 15512 15442 15524
rect 15657 15521 15669 15524
rect 15703 15521 15715 15555
rect 15657 15515 15715 15521
rect 15473 15487 15531 15493
rect 15473 15484 15485 15487
rect 14884 15456 14929 15484
rect 15304 15456 15485 15484
rect 14884 15444 14890 15456
rect 15473 15453 15485 15456
rect 15519 15453 15531 15487
rect 15473 15447 15531 15453
rect 16592 15416 16620 15660
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 20165 15691 20223 15697
rect 20165 15657 20177 15691
rect 20211 15688 20223 15691
rect 20254 15688 20260 15700
rect 20211 15660 20260 15688
rect 20211 15657 20223 15660
rect 20165 15651 20223 15657
rect 20254 15648 20260 15660
rect 20312 15648 20318 15700
rect 20441 15691 20499 15697
rect 20441 15657 20453 15691
rect 20487 15657 20499 15691
rect 20714 15688 20720 15700
rect 20675 15660 20720 15688
rect 20441 15651 20499 15657
rect 17494 15580 17500 15632
rect 17552 15620 17558 15632
rect 19797 15623 19855 15629
rect 19797 15620 19809 15623
rect 17552 15592 19809 15620
rect 17552 15580 17558 15592
rect 19797 15589 19809 15592
rect 19843 15589 19855 15623
rect 20456 15620 20484 15651
rect 20714 15648 20720 15660
rect 20772 15648 20778 15700
rect 20993 15691 21051 15697
rect 20993 15657 21005 15691
rect 21039 15657 21051 15691
rect 20993 15651 21051 15657
rect 20898 15620 20904 15632
rect 20456 15592 20904 15620
rect 19797 15583 19855 15589
rect 18233 15555 18291 15561
rect 18233 15521 18245 15555
rect 18279 15552 18291 15555
rect 19610 15552 19616 15564
rect 18279 15524 19616 15552
rect 18279 15521 18291 15524
rect 18233 15515 18291 15521
rect 19610 15512 19616 15524
rect 19668 15512 19674 15564
rect 19812 15552 19840 15583
rect 20898 15580 20904 15592
rect 20956 15580 20962 15632
rect 21008 15620 21036 15651
rect 21361 15623 21419 15629
rect 21361 15620 21373 15623
rect 21008 15592 21373 15620
rect 21361 15589 21373 15592
rect 21407 15589 21419 15623
rect 21361 15583 21419 15589
rect 19981 15555 20039 15561
rect 19981 15552 19993 15555
rect 19812 15524 19993 15552
rect 19981 15521 19993 15524
rect 20027 15521 20039 15555
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 19981 15515 20039 15521
rect 20088 15524 20269 15552
rect 17954 15484 17960 15496
rect 17915 15456 17960 15484
rect 17954 15444 17960 15456
rect 18012 15444 18018 15496
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 18141 15487 18199 15493
rect 18141 15484 18153 15487
rect 18104 15456 18153 15484
rect 18104 15444 18110 15456
rect 18141 15453 18153 15456
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 19705 15487 19763 15493
rect 19705 15453 19717 15487
rect 19751 15484 19763 15487
rect 20088 15484 20116 15524
rect 20257 15521 20269 15524
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 20438 15512 20444 15564
rect 20496 15552 20502 15564
rect 20533 15555 20591 15561
rect 20533 15552 20545 15555
rect 20496 15524 20545 15552
rect 20496 15512 20502 15524
rect 20533 15521 20545 15524
rect 20579 15521 20591 15555
rect 20533 15515 20591 15521
rect 20809 15555 20867 15561
rect 20809 15521 20821 15555
rect 20855 15521 20867 15555
rect 20809 15515 20867 15521
rect 19751 15456 20116 15484
rect 19751 15453 19763 15456
rect 19705 15447 19763 15453
rect 19720 15416 19748 15447
rect 20162 15444 20168 15496
rect 20220 15484 20226 15496
rect 20824 15484 20852 15515
rect 20220 15456 20852 15484
rect 20220 15444 20226 15456
rect 21542 15416 21548 15428
rect 14476 15388 16620 15416
rect 16684 15388 19748 15416
rect 21503 15388 21548 15416
rect 12115 15320 13308 15348
rect 14461 15351 14519 15357
rect 12115 15317 12127 15320
rect 12069 15311 12127 15317
rect 14461 15317 14473 15351
rect 14507 15348 14519 15351
rect 15194 15348 15200 15360
rect 14507 15320 15200 15348
rect 14507 15317 14519 15320
rect 14461 15311 14519 15317
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 15289 15351 15347 15357
rect 15289 15317 15301 15351
rect 15335 15348 15347 15351
rect 15930 15348 15936 15360
rect 15335 15320 15936 15348
rect 15335 15317 15347 15320
rect 15289 15311 15347 15317
rect 15930 15308 15936 15320
rect 15988 15308 15994 15360
rect 16114 15348 16120 15360
rect 16075 15320 16120 15348
rect 16114 15308 16120 15320
rect 16172 15308 16178 15360
rect 16206 15308 16212 15360
rect 16264 15348 16270 15360
rect 16684 15348 16712 15388
rect 21542 15376 21548 15388
rect 21600 15376 21606 15428
rect 16264 15320 16712 15348
rect 18601 15351 18659 15357
rect 16264 15308 16270 15320
rect 18601 15317 18613 15351
rect 18647 15348 18659 15351
rect 19518 15348 19524 15360
rect 18647 15320 19524 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 20438 15308 20444 15360
rect 20496 15348 20502 15360
rect 21085 15351 21143 15357
rect 21085 15348 21097 15351
rect 20496 15320 21097 15348
rect 20496 15308 20502 15320
rect 21085 15317 21097 15320
rect 21131 15317 21143 15351
rect 21085 15311 21143 15317
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 1946 15104 1952 15156
rect 2004 15144 2010 15156
rect 2317 15147 2375 15153
rect 2317 15144 2329 15147
rect 2004 15116 2329 15144
rect 2004 15104 2010 15116
rect 2317 15113 2329 15116
rect 2363 15113 2375 15147
rect 2317 15107 2375 15113
rect 2685 15147 2743 15153
rect 2685 15113 2697 15147
rect 2731 15144 2743 15147
rect 2866 15144 2872 15156
rect 2731 15116 2872 15144
rect 2731 15113 2743 15116
rect 2685 15107 2743 15113
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 4065 15147 4123 15153
rect 4065 15113 4077 15147
rect 4111 15144 4123 15147
rect 4246 15144 4252 15156
rect 4111 15116 4252 15144
rect 4111 15113 4123 15116
rect 4065 15107 4123 15113
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 5626 15104 5632 15156
rect 5684 15144 5690 15156
rect 6273 15147 6331 15153
rect 6273 15144 6285 15147
rect 5684 15116 6285 15144
rect 5684 15104 5690 15116
rect 6273 15113 6285 15116
rect 6319 15144 6331 15147
rect 6730 15144 6736 15156
rect 6319 15116 6736 15144
rect 6319 15113 6331 15116
rect 6273 15107 6331 15113
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 6825 15147 6883 15153
rect 6825 15113 6837 15147
rect 6871 15144 6883 15147
rect 7190 15144 7196 15156
rect 6871 15116 7196 15144
rect 6871 15113 6883 15116
rect 6825 15107 6883 15113
rect 1578 15036 1584 15088
rect 1636 15076 1642 15088
rect 2041 15079 2099 15085
rect 2041 15076 2053 15079
rect 1636 15048 2053 15076
rect 1636 15036 1642 15048
rect 2041 15045 2053 15048
rect 2087 15045 2099 15079
rect 3970 15076 3976 15088
rect 2041 15039 2099 15045
rect 2746 15048 3976 15076
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 14968 1458 15020
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2038 14940 2044 14952
rect 1995 14912 2044 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2038 14900 2044 14912
rect 2096 14900 2102 14952
rect 2222 14940 2228 14952
rect 2183 14912 2228 14940
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2501 14943 2559 14949
rect 2501 14909 2513 14943
rect 2547 14940 2559 14943
rect 2746 14940 2774 15048
rect 3970 15036 3976 15048
rect 4028 15036 4034 15088
rect 6546 15036 6552 15088
rect 6604 15076 6610 15088
rect 6840 15076 6868 15107
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 9401 15147 9459 15153
rect 9401 15113 9413 15147
rect 9447 15144 9459 15147
rect 10870 15144 10876 15156
rect 9447 15116 10876 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 11241 15147 11299 15153
rect 11241 15113 11253 15147
rect 11287 15144 11299 15147
rect 12342 15144 12348 15156
rect 11287 15116 12348 15144
rect 11287 15113 11299 15116
rect 11241 15107 11299 15113
rect 6604 15048 6868 15076
rect 6604 15036 6610 15048
rect 8202 15036 8208 15088
rect 8260 15076 8266 15088
rect 10321 15079 10379 15085
rect 10321 15076 10333 15079
rect 8260 15048 9996 15076
rect 8260 15036 8266 15048
rect 3234 15008 3240 15020
rect 3195 14980 3240 15008
rect 3234 14968 3240 14980
rect 3292 15008 3298 15020
rect 4617 15011 4675 15017
rect 4617 15008 4629 15011
rect 3292 14980 4629 15008
rect 3292 14968 3298 14980
rect 4617 14977 4629 14980
rect 4663 15008 4675 15011
rect 7742 15008 7748 15020
rect 4663 14980 5028 15008
rect 4663 14977 4675 14980
rect 4617 14971 4675 14977
rect 5000 14952 5028 14980
rect 6665 14980 7748 15008
rect 2547 14912 2774 14940
rect 3053 14943 3111 14949
rect 2547 14909 2559 14912
rect 2501 14903 2559 14909
rect 3053 14909 3065 14943
rect 3099 14940 3111 14943
rect 3099 14912 3832 14940
rect 3099 14909 3111 14912
rect 3053 14903 3111 14909
rect 1581 14875 1639 14881
rect 1581 14841 1593 14875
rect 1627 14872 1639 14875
rect 3145 14875 3203 14881
rect 3145 14872 3157 14875
rect 1627 14844 1808 14872
rect 1627 14841 1639 14844
rect 1581 14835 1639 14841
rect 1780 14813 1808 14844
rect 2746 14844 3157 14872
rect 1765 14807 1823 14813
rect 1765 14773 1777 14807
rect 1811 14773 1823 14807
rect 1765 14767 1823 14773
rect 2498 14764 2504 14816
rect 2556 14804 2562 14816
rect 2746 14804 2774 14844
rect 3145 14841 3157 14844
rect 3191 14841 3203 14875
rect 3145 14835 3203 14841
rect 3804 14816 3832 14912
rect 4154 14900 4160 14952
rect 4212 14940 4218 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4212 14912 4905 14940
rect 4212 14900 4218 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 4982 14900 4988 14952
rect 5040 14900 5046 14952
rect 5160 14943 5218 14949
rect 5160 14909 5172 14943
rect 5206 14940 5218 14943
rect 5534 14940 5540 14952
rect 5206 14912 5540 14940
rect 5206 14909 5218 14912
rect 5160 14903 5218 14909
rect 5534 14900 5540 14912
rect 5592 14940 5598 14952
rect 6665 14940 6693 14980
rect 7742 14968 7748 14980
rect 7800 15008 7806 15020
rect 7837 15011 7895 15017
rect 7837 15008 7849 15011
rect 7800 14980 7849 15008
rect 7800 14968 7806 14980
rect 7837 14977 7849 14980
rect 7883 14977 7895 15011
rect 7837 14971 7895 14977
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 15008 8907 15011
rect 9490 15008 9496 15020
rect 8895 14980 9496 15008
rect 8895 14977 8907 14980
rect 8849 14971 8907 14977
rect 9490 14968 9496 14980
rect 9548 14968 9554 15020
rect 9968 15017 9996 15048
rect 10060 15048 10333 15076
rect 9953 15011 10011 15017
rect 9953 14977 9965 15011
rect 9999 14977 10011 15011
rect 9953 14971 10011 14977
rect 5592 14912 6693 14940
rect 5592 14900 5598 14912
rect 7006 14900 7012 14952
rect 7064 14940 7070 14952
rect 8389 14943 8447 14949
rect 8389 14940 8401 14943
rect 7064 14912 8401 14940
rect 7064 14900 7070 14912
rect 8389 14909 8401 14912
rect 8435 14909 8447 14943
rect 8389 14903 8447 14909
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14940 9091 14943
rect 10060 14940 10088 15048
rect 10321 15045 10333 15048
rect 10367 15045 10379 15079
rect 10321 15039 10379 15045
rect 10137 15011 10195 15017
rect 10137 14977 10149 15011
rect 10183 15008 10195 15011
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 10183 14980 10977 15008
rect 10183 14977 10195 14980
rect 10137 14971 10195 14977
rect 10965 14977 10977 14980
rect 11011 15008 11023 15011
rect 11054 15008 11060 15020
rect 11011 14980 11060 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 9079 14912 10088 14940
rect 10689 14943 10747 14949
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 10689 14909 10701 14943
rect 10735 14940 10747 14943
rect 11256 14940 11284 15107
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 13909 15147 13967 15153
rect 13909 15144 13921 15147
rect 13872 15116 13921 15144
rect 13872 15104 13878 15116
rect 13909 15113 13921 15116
rect 13955 15113 13967 15147
rect 13909 15107 13967 15113
rect 14090 15104 14096 15156
rect 14148 15144 14154 15156
rect 16206 15144 16212 15156
rect 14148 15116 16212 15144
rect 14148 15104 14154 15116
rect 16206 15104 16212 15116
rect 16264 15104 16270 15156
rect 16390 15144 16396 15156
rect 16351 15116 16396 15144
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 20162 15144 20168 15156
rect 16500 15116 18460 15144
rect 20123 15116 20168 15144
rect 13078 15036 13084 15088
rect 13136 15076 13142 15088
rect 14829 15079 14887 15085
rect 14829 15076 14841 15079
rect 13136 15048 14841 15076
rect 13136 15036 13142 15048
rect 14829 15045 14841 15048
rect 14875 15045 14887 15079
rect 16500 15076 16528 15116
rect 14829 15039 14887 15045
rect 14936 15048 16528 15076
rect 18432 15076 18460 15116
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 20441 15147 20499 15153
rect 20441 15113 20453 15147
rect 20487 15144 20499 15147
rect 20622 15144 20628 15156
rect 20487 15116 20628 15144
rect 20487 15113 20499 15116
rect 20441 15107 20499 15113
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 18432 15048 20300 15076
rect 13170 14968 13176 15020
rect 13228 15008 13234 15020
rect 13265 15011 13323 15017
rect 13265 15008 13277 15011
rect 13228 14980 13277 15008
rect 13228 14968 13234 14980
rect 13265 14977 13277 14980
rect 13311 14977 13323 15011
rect 13449 15011 13507 15017
rect 13449 15008 13461 15011
rect 13265 14971 13323 14977
rect 13372 14980 13461 15008
rect 10735 14912 11284 14940
rect 10735 14909 10747 14912
rect 10689 14903 10747 14909
rect 11330 14900 11336 14952
rect 11388 14940 11394 14952
rect 11701 14943 11759 14949
rect 11701 14940 11713 14943
rect 11388 14912 11713 14940
rect 11388 14900 11394 14912
rect 11701 14909 11713 14912
rect 11747 14940 11759 14943
rect 11790 14940 11796 14952
rect 11747 14912 11796 14940
rect 11747 14909 11759 14912
rect 11701 14903 11759 14909
rect 11790 14900 11796 14912
rect 11848 14900 11854 14952
rect 11968 14943 12026 14949
rect 11968 14909 11980 14943
rect 12014 14940 12026 14943
rect 12434 14940 12440 14952
rect 12014 14912 12440 14940
rect 12014 14909 12026 14912
rect 11968 14903 12026 14909
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 12986 14900 12992 14952
rect 13044 14940 13050 14952
rect 13372 14940 13400 14980
rect 13449 14977 13461 14980
rect 13495 14977 13507 15011
rect 13449 14971 13507 14977
rect 13538 14968 13544 15020
rect 13596 15008 13602 15020
rect 14936 15008 14964 15048
rect 15470 15008 15476 15020
rect 13596 14980 14964 15008
rect 15431 14980 15476 15008
rect 13596 14968 13602 14980
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 15746 15008 15752 15020
rect 15707 14980 15752 15008
rect 15746 14968 15752 14980
rect 15804 14968 15810 15020
rect 15930 15008 15936 15020
rect 15891 14980 15936 15008
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 17402 14968 17408 15020
rect 17460 15008 17466 15020
rect 17497 15011 17555 15017
rect 17497 15008 17509 15011
rect 17460 14980 17509 15008
rect 17460 14968 17466 14980
rect 17497 14977 17509 14980
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 14553 14943 14611 14949
rect 14553 14940 14565 14943
rect 13044 14912 13400 14940
rect 14108 14912 14565 14940
rect 13044 14900 13050 14912
rect 14108 14884 14136 14912
rect 14553 14909 14565 14912
rect 14599 14940 14611 14943
rect 14642 14940 14648 14952
rect 14599 14912 14648 14940
rect 14599 14909 14611 14912
rect 14553 14903 14611 14909
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 16025 14943 16083 14949
rect 16025 14909 16037 14943
rect 16071 14940 16083 14943
rect 16114 14940 16120 14952
rect 16071 14912 16120 14940
rect 16071 14909 16083 14912
rect 16025 14903 16083 14909
rect 16114 14900 16120 14912
rect 16172 14900 16178 14952
rect 19518 14900 19524 14952
rect 19576 14940 19582 14952
rect 20272 14949 20300 15048
rect 21542 15008 21548 15020
rect 21503 14980 21548 15008
rect 21542 14968 21548 14980
rect 21600 14968 21606 15020
rect 19981 14943 20039 14949
rect 19981 14940 19993 14943
rect 19576 14912 19993 14940
rect 19576 14900 19582 14912
rect 19981 14909 19993 14912
rect 20027 14909 20039 14943
rect 19981 14903 20039 14909
rect 20257 14943 20315 14949
rect 20257 14909 20269 14943
rect 20303 14909 20315 14943
rect 20257 14903 20315 14909
rect 20809 14943 20867 14949
rect 20809 14909 20821 14943
rect 20855 14909 20867 14943
rect 20809 14903 20867 14909
rect 7193 14875 7251 14881
rect 7193 14841 7205 14875
rect 7239 14872 7251 14875
rect 7653 14875 7711 14881
rect 7653 14872 7665 14875
rect 7239 14844 7665 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 7653 14841 7665 14844
rect 7699 14872 7711 14875
rect 7834 14872 7840 14884
rect 7699 14844 7840 14872
rect 7699 14841 7711 14844
rect 7653 14835 7711 14841
rect 7834 14832 7840 14844
rect 7892 14832 7898 14884
rect 9582 14832 9588 14884
rect 9640 14872 9646 14884
rect 10318 14872 10324 14884
rect 9640 14844 10324 14872
rect 9640 14832 9646 14844
rect 10318 14832 10324 14844
rect 10376 14832 10382 14884
rect 10594 14832 10600 14884
rect 10652 14872 10658 14884
rect 10652 14844 11100 14872
rect 10652 14832 10658 14844
rect 3510 14804 3516 14816
rect 2556 14776 2774 14804
rect 3471 14776 3516 14804
rect 2556 14764 2562 14776
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 3786 14804 3792 14816
rect 3747 14776 3792 14804
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 4430 14804 4436 14816
rect 4120 14776 4436 14804
rect 4120 14764 4126 14776
rect 4430 14764 4436 14776
rect 4488 14764 4494 14816
rect 4525 14807 4583 14813
rect 4525 14773 4537 14807
rect 4571 14804 4583 14807
rect 5258 14804 5264 14816
rect 4571 14776 5264 14804
rect 4571 14773 4583 14776
rect 4525 14767 4583 14773
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 5994 14764 6000 14816
rect 6052 14804 6058 14816
rect 6638 14804 6644 14816
rect 6052 14776 6644 14804
rect 6052 14764 6058 14776
rect 6638 14764 6644 14776
rect 6696 14764 6702 14816
rect 7282 14804 7288 14816
rect 7243 14776 7288 14804
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 7374 14764 7380 14816
rect 7432 14804 7438 14816
rect 7745 14807 7803 14813
rect 7745 14804 7757 14807
rect 7432 14776 7757 14804
rect 7432 14764 7438 14776
rect 7745 14773 7757 14776
rect 7791 14804 7803 14807
rect 8113 14807 8171 14813
rect 8113 14804 8125 14807
rect 7791 14776 8125 14804
rect 7791 14773 7803 14776
rect 7745 14767 7803 14773
rect 8113 14773 8125 14776
rect 8159 14773 8171 14807
rect 8570 14804 8576 14816
rect 8531 14776 8576 14804
rect 8113 14767 8171 14773
rect 8570 14764 8576 14776
rect 8628 14764 8634 14816
rect 8941 14807 8999 14813
rect 8941 14773 8953 14807
rect 8987 14804 8999 14807
rect 9493 14807 9551 14813
rect 9493 14804 9505 14807
rect 8987 14776 9505 14804
rect 8987 14773 8999 14776
rect 8941 14767 8999 14773
rect 9493 14773 9505 14776
rect 9539 14773 9551 14807
rect 9858 14804 9864 14816
rect 9819 14776 9864 14804
rect 9493 14767 9551 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 10778 14804 10784 14816
rect 10739 14776 10784 14804
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11072 14804 11100 14844
rect 11146 14832 11152 14884
rect 11204 14872 11210 14884
rect 11425 14875 11483 14881
rect 11425 14872 11437 14875
rect 11204 14844 11437 14872
rect 11204 14832 11210 14844
rect 11425 14841 11437 14844
rect 11471 14872 11483 14875
rect 12158 14872 12164 14884
rect 11471 14844 12164 14872
rect 11471 14841 11483 14844
rect 11425 14835 11483 14841
rect 12158 14832 12164 14844
rect 12216 14832 12222 14884
rect 13541 14875 13599 14881
rect 13541 14841 13553 14875
rect 13587 14872 13599 14875
rect 14090 14872 14096 14884
rect 13587 14844 14096 14872
rect 13587 14841 13599 14844
rect 13541 14835 13599 14841
rect 14090 14832 14096 14844
rect 14148 14832 14154 14884
rect 14826 14872 14832 14884
rect 14200 14844 14832 14872
rect 14200 14816 14228 14844
rect 14826 14832 14832 14844
rect 14884 14832 14890 14884
rect 15197 14875 15255 14881
rect 15197 14841 15209 14875
rect 15243 14872 15255 14875
rect 16942 14872 16948 14884
rect 15243 14844 16948 14872
rect 15243 14841 15255 14844
rect 15197 14835 15255 14841
rect 16942 14832 16948 14844
rect 17000 14832 17006 14884
rect 17218 14832 17224 14884
rect 17276 14872 17282 14884
rect 17742 14875 17800 14881
rect 17742 14872 17754 14875
rect 17276 14844 17754 14872
rect 17276 14832 17282 14844
rect 17742 14841 17754 14844
rect 17788 14841 17800 14875
rect 17742 14835 17800 14841
rect 20824 14816 20852 14903
rect 21361 14875 21419 14881
rect 21361 14841 21373 14875
rect 21407 14841 21419 14875
rect 21361 14835 21419 14841
rect 12342 14804 12348 14816
rect 11072 14776 12348 14804
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 13081 14807 13139 14813
rect 13081 14773 13093 14807
rect 13127 14804 13139 14807
rect 13170 14804 13176 14816
rect 13127 14776 13176 14804
rect 13127 14773 13139 14776
rect 13081 14767 13139 14773
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 13906 14804 13912 14816
rect 13320 14776 13912 14804
rect 13320 14764 13326 14776
rect 13906 14764 13912 14776
rect 13964 14804 13970 14816
rect 14001 14807 14059 14813
rect 14001 14804 14013 14807
rect 13964 14776 14013 14804
rect 13964 14764 13970 14776
rect 14001 14773 14013 14776
rect 14047 14773 14059 14807
rect 14182 14804 14188 14816
rect 14143 14776 14188 14804
rect 14001 14767 14059 14773
rect 14182 14764 14188 14776
rect 14240 14764 14246 14816
rect 14366 14804 14372 14816
rect 14327 14776 14372 14804
rect 14366 14764 14372 14776
rect 14424 14764 14430 14816
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15930 14804 15936 14816
rect 15335 14776 15936 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15930 14764 15936 14776
rect 15988 14764 15994 14816
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18877 14807 18935 14813
rect 18877 14804 18889 14807
rect 18012 14776 18889 14804
rect 18012 14764 18018 14776
rect 18877 14773 18889 14776
rect 18923 14773 18935 14807
rect 18877 14767 18935 14773
rect 20717 14807 20775 14813
rect 20717 14773 20729 14807
rect 20763 14804 20775 14807
rect 20806 14804 20812 14816
rect 20763 14776 20812 14804
rect 20763 14773 20775 14776
rect 20717 14767 20775 14773
rect 20806 14764 20812 14776
rect 20864 14764 20870 14816
rect 20993 14807 21051 14813
rect 20993 14773 21005 14807
rect 21039 14804 21051 14807
rect 21376 14804 21404 14835
rect 21039 14776 21404 14804
rect 21039 14773 21051 14776
rect 20993 14767 21051 14773
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 2133 14603 2191 14609
rect 2133 14600 2145 14603
rect 1964 14572 2145 14600
rect 1964 14541 1992 14572
rect 2133 14569 2145 14572
rect 2179 14569 2191 14603
rect 2133 14563 2191 14569
rect 2593 14603 2651 14609
rect 2593 14569 2605 14603
rect 2639 14600 2651 14603
rect 2774 14600 2780 14612
rect 2639 14572 2780 14600
rect 2639 14569 2651 14572
rect 2593 14563 2651 14569
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 2961 14603 3019 14609
rect 2961 14569 2973 14603
rect 3007 14600 3019 14603
rect 3510 14600 3516 14612
rect 3007 14572 3516 14600
rect 3007 14569 3019 14572
rect 2961 14563 3019 14569
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 6457 14603 6515 14609
rect 6457 14600 6469 14603
rect 4212 14572 6469 14600
rect 4212 14560 4218 14572
rect 6457 14569 6469 14572
rect 6503 14569 6515 14603
rect 6457 14563 6515 14569
rect 6733 14603 6791 14609
rect 6733 14569 6745 14603
rect 6779 14600 6791 14603
rect 6914 14600 6920 14612
rect 6779 14572 6920 14600
rect 6779 14569 6791 14572
rect 6733 14563 6791 14569
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 7101 14603 7159 14609
rect 7101 14569 7113 14603
rect 7147 14600 7159 14603
rect 7282 14600 7288 14612
rect 7147 14572 7288 14600
rect 7147 14569 7159 14572
rect 7101 14563 7159 14569
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 10965 14603 11023 14609
rect 10965 14600 10977 14603
rect 7484 14572 10977 14600
rect 1949 14535 2007 14541
rect 1949 14501 1961 14535
rect 1995 14501 2007 14535
rect 1949 14495 2007 14501
rect 2038 14492 2044 14544
rect 2096 14532 2102 14544
rect 2866 14532 2872 14544
rect 2096 14504 2872 14532
rect 2096 14492 2102 14504
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 3053 14535 3111 14541
rect 3053 14501 3065 14535
rect 3099 14532 3111 14535
rect 3142 14532 3148 14544
rect 3099 14504 3148 14532
rect 3099 14501 3111 14504
rect 3053 14495 3111 14501
rect 3142 14492 3148 14504
rect 3200 14492 3206 14544
rect 3421 14535 3479 14541
rect 3421 14501 3433 14535
rect 3467 14532 3479 14535
rect 3694 14532 3700 14544
rect 3467 14504 3700 14532
rect 3467 14501 3479 14504
rect 3421 14495 3479 14501
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14433 1639 14467
rect 1581 14427 1639 14433
rect 2317 14467 2375 14473
rect 2317 14433 2329 14467
rect 2363 14464 2375 14467
rect 3436 14464 3464 14495
rect 3694 14492 3700 14504
rect 3752 14532 3758 14544
rect 4338 14532 4344 14544
rect 3752 14504 4344 14532
rect 3752 14492 3758 14504
rect 4338 14492 4344 14504
rect 4396 14492 4402 14544
rect 5813 14535 5871 14541
rect 5813 14501 5825 14535
rect 5859 14532 5871 14535
rect 6270 14532 6276 14544
rect 5859 14504 6276 14532
rect 5859 14501 5871 14504
rect 5813 14495 5871 14501
rect 6270 14492 6276 14504
rect 6328 14532 6334 14544
rect 6365 14535 6423 14541
rect 6365 14532 6377 14535
rect 6328 14504 6377 14532
rect 6328 14492 6334 14504
rect 6365 14501 6377 14504
rect 6411 14532 6423 14535
rect 7484 14532 7512 14572
rect 10965 14569 10977 14572
rect 11011 14600 11023 14603
rect 11146 14600 11152 14612
rect 11011 14572 11152 14600
rect 11011 14569 11023 14572
rect 10965 14563 11023 14569
rect 11146 14560 11152 14572
rect 11204 14560 11210 14612
rect 12158 14600 12164 14612
rect 11256 14572 12164 14600
rect 6411 14504 7512 14532
rect 6411 14501 6423 14504
rect 6365 14495 6423 14501
rect 7558 14492 7564 14544
rect 7616 14532 7622 14544
rect 7806 14535 7864 14541
rect 7806 14532 7818 14535
rect 7616 14504 7818 14532
rect 7616 14492 7622 14504
rect 7806 14501 7818 14504
rect 7852 14501 7864 14535
rect 7806 14495 7864 14501
rect 4246 14464 4252 14476
rect 2363 14436 3464 14464
rect 4207 14436 4252 14464
rect 2363 14433 2375 14436
rect 2317 14427 2375 14433
rect 1596 14396 1624 14427
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 5905 14467 5963 14473
rect 5905 14433 5917 14467
rect 5951 14464 5963 14467
rect 6454 14464 6460 14476
rect 5951 14436 6460 14464
rect 5951 14433 5963 14436
rect 5905 14427 5963 14433
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 6641 14467 6699 14473
rect 6641 14433 6653 14467
rect 6687 14464 6699 14467
rect 7006 14464 7012 14476
rect 6687 14436 7012 14464
rect 6687 14433 6699 14436
rect 6641 14427 6699 14433
rect 7006 14424 7012 14436
rect 7064 14424 7070 14476
rect 7821 14464 7849 14495
rect 8846 14492 8852 14544
rect 8904 14532 8910 14544
rect 9582 14532 9588 14544
rect 8904 14504 9588 14532
rect 8904 14492 8910 14504
rect 9582 14492 9588 14504
rect 9640 14532 9646 14544
rect 10260 14535 10318 14541
rect 10260 14532 10272 14535
rect 9640 14504 10272 14532
rect 9640 14492 9646 14504
rect 10260 14501 10272 14504
rect 10306 14532 10318 14535
rect 11054 14532 11060 14544
rect 10306 14504 11060 14532
rect 10306 14501 10318 14504
rect 10260 14495 10318 14501
rect 11054 14492 11060 14504
rect 11112 14532 11118 14544
rect 11256 14532 11284 14572
rect 12158 14560 12164 14572
rect 12216 14560 12222 14612
rect 12526 14560 12532 14612
rect 12584 14600 12590 14612
rect 12897 14603 12955 14609
rect 12897 14600 12909 14603
rect 12584 14572 12909 14600
rect 12584 14560 12590 14572
rect 12897 14569 12909 14572
rect 12943 14600 12955 14603
rect 13998 14600 14004 14612
rect 12943 14572 14004 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 18966 14600 18972 14612
rect 15663 14572 18972 14600
rect 12345 14535 12403 14541
rect 12345 14532 12357 14535
rect 11112 14504 11284 14532
rect 11716 14504 12357 14532
rect 11112 14492 11118 14504
rect 11422 14464 11428 14476
rect 7821 14436 10640 14464
rect 2406 14396 2412 14408
rect 1596 14368 2412 14396
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 3234 14396 3240 14408
rect 3195 14368 3240 14396
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3697 14399 3755 14405
rect 3697 14365 3709 14399
rect 3743 14396 3755 14399
rect 3970 14396 3976 14408
rect 3743 14368 3976 14396
rect 3743 14365 3755 14368
rect 3697 14359 3755 14365
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4338 14396 4344 14408
rect 4299 14368 4344 14396
rect 4338 14356 4344 14368
rect 4396 14356 4402 14408
rect 4525 14399 4583 14405
rect 4525 14365 4537 14399
rect 4571 14396 4583 14399
rect 5718 14396 5724 14408
rect 4571 14368 5724 14396
rect 4571 14365 4583 14368
rect 4525 14359 4583 14365
rect 5718 14356 5724 14368
rect 5776 14356 5782 14408
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14396 6147 14399
rect 6178 14396 6184 14408
rect 6135 14368 6184 14396
rect 6135 14365 6147 14368
rect 6089 14359 6147 14365
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 7190 14396 7196 14408
rect 7151 14368 7196 14396
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 7285 14399 7343 14405
rect 7285 14365 7297 14399
rect 7331 14365 7343 14399
rect 7285 14359 7343 14365
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14365 10563 14399
rect 10612 14396 10640 14436
rect 11072 14436 11428 14464
rect 10686 14396 10692 14408
rect 10612 14368 10692 14396
rect 10505 14359 10563 14365
rect 2866 14288 2872 14340
rect 2924 14328 2930 14340
rect 3881 14331 3939 14337
rect 3881 14328 3893 14331
rect 2924 14300 3893 14328
rect 2924 14288 2930 14300
rect 3881 14297 3893 14300
rect 3927 14297 3939 14331
rect 3881 14291 3939 14297
rect 4430 14288 4436 14340
rect 4488 14288 4494 14340
rect 5445 14331 5503 14337
rect 5445 14297 5457 14331
rect 5491 14328 5503 14331
rect 5534 14328 5540 14340
rect 5491 14300 5540 14328
rect 5491 14297 5503 14300
rect 5445 14291 5503 14297
rect 5534 14288 5540 14300
rect 5592 14288 5598 14340
rect 6730 14288 6736 14340
rect 6788 14328 6794 14340
rect 7300 14328 7328 14359
rect 7466 14328 7472 14340
rect 6788 14300 7472 14328
rect 6788 14288 6794 14300
rect 7466 14288 7472 14300
rect 7524 14288 7530 14340
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2498 14260 2504 14272
rect 2459 14232 2504 14260
rect 2498 14220 2504 14232
rect 2556 14220 2562 14272
rect 4448 14260 4476 14288
rect 4982 14260 4988 14272
rect 4448 14232 4988 14260
rect 4982 14220 4988 14232
rect 5040 14220 5046 14272
rect 5166 14260 5172 14272
rect 5127 14232 5172 14260
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 7576 14260 7604 14359
rect 8846 14288 8852 14340
rect 8904 14328 8910 14340
rect 8941 14331 8999 14337
rect 8941 14328 8953 14331
rect 8904 14300 8953 14328
rect 8904 14288 8910 14300
rect 8941 14297 8953 14300
rect 8987 14297 8999 14331
rect 9398 14328 9404 14340
rect 8941 14291 8999 14297
rect 9028 14300 9404 14328
rect 8570 14260 8576 14272
rect 7576 14232 8576 14260
rect 8570 14220 8576 14232
rect 8628 14260 8634 14272
rect 9028 14260 9056 14300
rect 9398 14288 9404 14300
rect 9456 14328 9462 14340
rect 9456 14300 9628 14328
rect 9456 14288 9462 14300
rect 8628 14232 9056 14260
rect 9125 14263 9183 14269
rect 8628 14220 8634 14232
rect 9125 14229 9137 14263
rect 9171 14260 9183 14263
rect 9490 14260 9496 14272
rect 9171 14232 9496 14260
rect 9171 14229 9183 14232
rect 9125 14223 9183 14229
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 9600 14260 9628 14300
rect 10520 14260 10548 14359
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 11072 14405 11100 14436
rect 11422 14424 11428 14436
rect 11480 14464 11486 14476
rect 11716 14464 11744 14504
rect 12345 14501 12357 14504
rect 12391 14532 12403 14535
rect 12618 14532 12624 14544
rect 12391 14504 12624 14532
rect 12391 14501 12403 14504
rect 12345 14495 12403 14501
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 13630 14492 13636 14544
rect 13688 14532 13694 14544
rect 15470 14532 15476 14544
rect 15528 14541 15534 14544
rect 13688 14504 15476 14532
rect 13688 14492 13694 14504
rect 15470 14492 15476 14504
rect 15528 14532 15540 14541
rect 15528 14504 15573 14532
rect 15528 14495 15540 14504
rect 15528 14492 15534 14495
rect 11480 14436 11744 14464
rect 11793 14467 11851 14473
rect 11480 14424 11486 14436
rect 11793 14433 11805 14467
rect 11839 14433 11851 14467
rect 11793 14427 11851 14433
rect 11885 14467 11943 14473
rect 11885 14433 11897 14467
rect 11931 14464 11943 14467
rect 11974 14464 11980 14476
rect 11931 14436 11980 14464
rect 11931 14433 11943 14436
rect 11885 14427 11943 14433
rect 11057 14399 11115 14405
rect 11057 14365 11069 14399
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 10597 14331 10655 14337
rect 10597 14297 10609 14331
rect 10643 14328 10655 14331
rect 10778 14328 10784 14340
rect 10643 14300 10784 14328
rect 10643 14297 10655 14300
rect 10597 14291 10655 14297
rect 10778 14288 10784 14300
rect 10836 14288 10842 14340
rect 11164 14328 11192 14359
rect 10980 14300 11192 14328
rect 9600 14232 10548 14260
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 10980 14260 11008 14300
rect 11808 14272 11836 14427
rect 11974 14424 11980 14436
rect 12032 14464 12038 14476
rect 13541 14467 13599 14473
rect 12032 14436 13492 14464
rect 12032 14424 12038 14436
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14396 12127 14399
rect 12158 14396 12164 14408
rect 12115 14368 12164 14396
rect 12115 14365 12127 14368
rect 12069 14359 12127 14365
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12621 14399 12679 14405
rect 12621 14396 12633 14399
rect 12492 14368 12633 14396
rect 12492 14356 12498 14368
rect 12621 14365 12633 14368
rect 12667 14365 12679 14399
rect 12802 14396 12808 14408
rect 12763 14368 12808 14396
rect 12621 14359 12679 14365
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 12986 14356 12992 14408
rect 13044 14396 13050 14408
rect 13464 14396 13492 14436
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 14550 14464 14556 14476
rect 13587 14436 14556 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 15663 14464 15691 14572
rect 18966 14560 18972 14572
rect 19024 14560 19030 14612
rect 19610 14600 19616 14612
rect 19571 14572 19616 14600
rect 19610 14560 19616 14572
rect 19668 14560 19674 14612
rect 20809 14603 20867 14609
rect 20809 14569 20821 14603
rect 20855 14600 20867 14603
rect 20855 14572 21036 14600
rect 20855 14569 20867 14572
rect 20809 14563 20867 14569
rect 17252 14535 17310 14541
rect 17252 14501 17264 14535
rect 17298 14532 17310 14535
rect 17954 14532 17960 14544
rect 17298 14504 17960 14532
rect 17298 14501 17310 14504
rect 17252 14495 17310 14501
rect 17954 14492 17960 14504
rect 18012 14492 18018 14544
rect 21008 14541 21036 14572
rect 20993 14535 21051 14541
rect 20993 14501 21005 14535
rect 21039 14501 21051 14535
rect 21174 14532 21180 14544
rect 21135 14504 21180 14532
rect 20993 14495 21051 14501
rect 21174 14492 21180 14504
rect 21232 14492 21238 14544
rect 14651 14436 15691 14464
rect 15749 14467 15807 14473
rect 14651 14396 14679 14436
rect 15749 14433 15761 14467
rect 15795 14464 15807 14467
rect 16850 14464 16856 14476
rect 15795 14436 16856 14464
rect 15795 14433 15807 14436
rect 15749 14427 15807 14433
rect 16850 14424 16856 14436
rect 16908 14464 16914 14476
rect 17402 14464 17408 14476
rect 16908 14436 17408 14464
rect 16908 14424 16914 14436
rect 17402 14424 17408 14436
rect 17460 14464 17466 14476
rect 17497 14467 17555 14473
rect 17497 14464 17509 14467
rect 17460 14436 17509 14464
rect 17460 14424 17466 14436
rect 17497 14433 17509 14436
rect 17543 14464 17555 14467
rect 17589 14467 17647 14473
rect 17589 14464 17601 14467
rect 17543 14436 17601 14464
rect 17543 14433 17555 14436
rect 17497 14427 17555 14433
rect 17589 14433 17601 14436
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 17856 14467 17914 14473
rect 17856 14433 17868 14467
rect 17902 14464 17914 14467
rect 18138 14464 18144 14476
rect 17902 14436 18144 14464
rect 17902 14433 17914 14436
rect 17856 14427 17914 14433
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 19518 14424 19524 14476
rect 19576 14464 19582 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19576 14436 19993 14464
rect 19576 14424 19582 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 20622 14464 20628 14476
rect 20583 14436 20628 14464
rect 19981 14427 20039 14433
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 21358 14464 21364 14476
rect 21319 14436 21364 14464
rect 21358 14424 21364 14436
rect 21416 14424 21422 14476
rect 19058 14396 19064 14408
rect 13044 14368 13308 14396
rect 13464 14368 14679 14396
rect 19019 14368 19064 14396
rect 13044 14356 13050 14368
rect 13280 14337 13308 14368
rect 19058 14356 19064 14368
rect 19116 14356 19122 14408
rect 19150 14356 19156 14408
rect 19208 14396 19214 14408
rect 20073 14399 20131 14405
rect 20073 14396 20085 14399
rect 19208 14368 20085 14396
rect 19208 14356 19214 14368
rect 20073 14365 20085 14368
rect 20119 14365 20131 14399
rect 20073 14359 20131 14365
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14365 20223 14399
rect 20165 14359 20223 14365
rect 13265 14331 13323 14337
rect 13265 14297 13277 14331
rect 13311 14297 13323 14331
rect 20180 14328 20208 14359
rect 21542 14328 21548 14340
rect 13265 14291 13323 14297
rect 18984 14300 20208 14328
rect 21503 14300 21548 14328
rect 10744 14232 11008 14260
rect 10744 14220 10750 14232
rect 11054 14220 11060 14272
rect 11112 14260 11118 14272
rect 11425 14263 11483 14269
rect 11425 14260 11437 14263
rect 11112 14232 11437 14260
rect 11112 14220 11118 14232
rect 11425 14229 11437 14232
rect 11471 14229 11483 14263
rect 11425 14223 11483 14229
rect 11790 14220 11796 14272
rect 11848 14220 11854 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 13354 14260 13360 14272
rect 11940 14232 13360 14260
rect 11940 14220 11946 14232
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 14369 14263 14427 14269
rect 14369 14260 14381 14263
rect 13504 14232 14381 14260
rect 13504 14220 13510 14232
rect 14369 14229 14381 14232
rect 14415 14260 14427 14263
rect 14734 14260 14740 14272
rect 14415 14232 14740 14260
rect 14415 14229 14427 14232
rect 14369 14223 14427 14229
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 16114 14260 16120 14272
rect 16075 14232 16120 14260
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 17218 14220 17224 14272
rect 17276 14260 17282 14272
rect 18984 14269 19012 14300
rect 21542 14288 21548 14300
rect 21600 14288 21606 14340
rect 18969 14263 19027 14269
rect 18969 14260 18981 14263
rect 17276 14232 18981 14260
rect 17276 14220 17282 14232
rect 18969 14229 18981 14232
rect 19015 14229 19027 14263
rect 18969 14223 19027 14229
rect 20533 14263 20591 14269
rect 20533 14229 20545 14263
rect 20579 14260 20591 14263
rect 20622 14260 20628 14272
rect 20579 14232 20628 14260
rect 20579 14229 20591 14232
rect 20533 14223 20591 14229
rect 20622 14220 20628 14232
rect 20680 14220 20686 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 2222 14016 2228 14068
rect 2280 14056 2286 14068
rect 2685 14059 2743 14065
rect 2685 14056 2697 14059
rect 2280 14028 2697 14056
rect 2280 14016 2286 14028
rect 2685 14025 2697 14028
rect 2731 14025 2743 14059
rect 2685 14019 2743 14025
rect 2958 14016 2964 14068
rect 3016 14056 3022 14068
rect 5810 14056 5816 14068
rect 3016 14028 5816 14056
rect 3016 14016 3022 14028
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 7650 14016 7656 14068
rect 7708 14056 7714 14068
rect 8021 14059 8079 14065
rect 8021 14056 8033 14059
rect 7708 14028 8033 14056
rect 7708 14016 7714 14028
rect 8021 14025 8033 14028
rect 8067 14025 8079 14059
rect 8021 14019 8079 14025
rect 9858 14016 9864 14068
rect 9916 14056 9922 14068
rect 10229 14059 10287 14065
rect 10229 14056 10241 14059
rect 9916 14028 10241 14056
rect 9916 14016 9922 14028
rect 10229 14025 10241 14028
rect 10275 14025 10287 14059
rect 12526 14056 12532 14068
rect 10229 14019 10287 14025
rect 10612 14028 12532 14056
rect 2133 13991 2191 13997
rect 2133 13957 2145 13991
rect 2179 13957 2191 13991
rect 2406 13988 2412 14000
rect 2367 13960 2412 13988
rect 2133 13951 2191 13957
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 1762 13852 1768 13864
rect 1723 13824 1768 13852
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 1949 13855 2007 13861
rect 1949 13821 1961 13855
rect 1995 13852 2007 13855
rect 2148 13852 2176 13951
rect 2406 13948 2412 13960
rect 2464 13948 2470 14000
rect 3237 13991 3295 13997
rect 3237 13957 3249 13991
rect 3283 13988 3295 13991
rect 3878 13988 3884 14000
rect 3283 13960 3884 13988
rect 3283 13957 3295 13960
rect 3237 13951 3295 13957
rect 3252 13920 3280 13951
rect 3878 13948 3884 13960
rect 3936 13948 3942 14000
rect 4890 13948 4896 14000
rect 4948 13988 4954 14000
rect 5537 13991 5595 13997
rect 5537 13988 5549 13991
rect 4948 13960 5549 13988
rect 4948 13948 4954 13960
rect 5537 13957 5549 13960
rect 5583 13957 5595 13991
rect 6457 13991 6515 13997
rect 6457 13988 6469 13991
rect 5537 13951 5595 13957
rect 6012 13960 6469 13988
rect 5626 13920 5632 13932
rect 2608 13892 3280 13920
rect 4816 13892 5632 13920
rect 2314 13852 2320 13864
rect 1995 13824 2176 13852
rect 2275 13824 2320 13852
rect 1995 13821 2007 13824
rect 1949 13815 2007 13821
rect 2314 13812 2320 13824
rect 2372 13812 2378 13864
rect 2608 13861 2636 13892
rect 2593 13855 2651 13861
rect 2593 13821 2605 13855
rect 2639 13821 2651 13855
rect 2593 13815 2651 13821
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13852 2927 13855
rect 4816 13852 4844 13892
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 6012 13929 6040 13960
rect 6457 13957 6469 13960
rect 6503 13957 6515 13991
rect 6457 13951 6515 13957
rect 7116 13960 7788 13988
rect 5997 13923 6055 13929
rect 5997 13889 6009 13923
rect 6043 13889 6055 13923
rect 6178 13920 6184 13932
rect 6139 13892 6184 13920
rect 5997 13883 6055 13889
rect 6178 13880 6184 13892
rect 6236 13880 6242 13932
rect 6638 13880 6644 13932
rect 6696 13920 6702 13932
rect 7009 13923 7067 13929
rect 7009 13920 7021 13923
rect 6696 13892 7021 13920
rect 6696 13880 6702 13892
rect 7009 13889 7021 13892
rect 7055 13889 7067 13923
rect 7009 13883 7067 13889
rect 2915 13824 4844 13852
rect 4893 13855 4951 13861
rect 2915 13821 2927 13824
rect 2869 13815 2927 13821
rect 4893 13821 4905 13855
rect 4939 13852 4951 13855
rect 5350 13852 5356 13864
rect 4939 13824 5356 13852
rect 4939 13821 4951 13824
rect 4893 13815 4951 13821
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 5445 13855 5503 13861
rect 5445 13821 5457 13855
rect 5491 13852 5503 13855
rect 5902 13852 5908 13864
rect 5491 13824 5908 13852
rect 5491 13821 5503 13824
rect 5445 13815 5503 13821
rect 5902 13812 5908 13824
rect 5960 13852 5966 13864
rect 6917 13855 6975 13861
rect 6917 13852 6929 13855
rect 5960 13824 6929 13852
rect 5960 13812 5966 13824
rect 6917 13821 6929 13824
rect 6963 13852 6975 13855
rect 7116 13852 7144 13960
rect 7466 13920 7472 13932
rect 7427 13892 7472 13920
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 7760 13864 7788 13960
rect 9214 13948 9220 14000
rect 9272 13988 9278 14000
rect 10612 13988 10640 14028
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 16482 14056 16488 14068
rect 13412 14028 15148 14056
rect 16395 14028 16488 14056
rect 13412 14016 13418 14028
rect 9272 13960 10640 13988
rect 9272 13948 9278 13960
rect 10686 13948 10692 14000
rect 10744 13988 10750 14000
rect 11333 13991 11391 13997
rect 10744 13960 10824 13988
rect 10744 13948 10750 13960
rect 9582 13920 9588 13932
rect 9543 13892 9588 13920
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 10796 13929 10824 13960
rect 11333 13957 11345 13991
rect 11379 13988 11391 13991
rect 11974 13988 11980 14000
rect 11379 13960 11980 13988
rect 11379 13957 11391 13960
rect 11333 13951 11391 13957
rect 11974 13948 11980 13960
rect 12032 13948 12038 14000
rect 13541 13991 13599 13997
rect 13541 13957 13553 13991
rect 13587 13988 13599 13991
rect 13630 13988 13636 14000
rect 13587 13960 13636 13988
rect 13587 13957 13599 13960
rect 13541 13951 13599 13957
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13889 10839 13923
rect 11882 13920 11888 13932
rect 11843 13892 11888 13920
rect 10781 13883 10839 13889
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 12805 13923 12863 13929
rect 12805 13889 12817 13923
rect 12851 13920 12863 13923
rect 13446 13920 13452 13932
rect 12851 13892 13452 13920
rect 12851 13889 12863 13892
rect 12805 13883 12863 13889
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 15120 13929 15148 14028
rect 16482 14016 16488 14028
rect 16540 14056 16546 14068
rect 16942 14056 16948 14068
rect 16540 14028 16620 14056
rect 16903 14028 16948 14056
rect 16540 14016 16546 14028
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13889 15163 13923
rect 16592 13920 16620 14028
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 19150 14056 19156 14068
rect 18739 14028 19156 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 19518 14056 19524 14068
rect 19479 14028 19524 14056
rect 19518 14016 19524 14028
rect 19576 14016 19582 14068
rect 20993 14059 21051 14065
rect 20993 14025 21005 14059
rect 21039 14056 21051 14059
rect 21358 14056 21364 14068
rect 21039 14028 21364 14056
rect 21039 14025 21051 14028
rect 20993 14019 21051 14025
rect 21358 14016 21364 14028
rect 21416 14016 21422 14068
rect 16666 13948 16672 14000
rect 16724 13988 16730 14000
rect 20717 13991 20775 13997
rect 20717 13988 20729 13991
rect 16724 13960 20729 13988
rect 16724 13948 16730 13960
rect 20717 13957 20729 13960
rect 20763 13957 20775 13991
rect 20717 13951 20775 13957
rect 17497 13923 17555 13929
rect 17497 13920 17509 13923
rect 16592 13892 17509 13920
rect 15105 13883 15163 13889
rect 17497 13889 17509 13892
rect 17543 13889 17555 13923
rect 18138 13920 18144 13932
rect 18051 13892 18144 13920
rect 17497 13883 17555 13889
rect 18138 13880 18144 13892
rect 18196 13920 18202 13932
rect 18874 13920 18880 13932
rect 18196 13892 18880 13920
rect 18196 13880 18202 13892
rect 18874 13880 18880 13892
rect 18932 13880 18938 13932
rect 6963 13824 7144 13852
rect 6963 13821 6975 13824
rect 6917 13815 6975 13821
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 7561 13855 7619 13861
rect 7561 13852 7573 13855
rect 7340 13824 7573 13852
rect 7340 13812 7346 13824
rect 7561 13821 7573 13824
rect 7607 13821 7619 13855
rect 7561 13815 7619 13821
rect 7742 13812 7748 13864
rect 7800 13812 7806 13864
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 11330 13852 11336 13864
rect 11195 13824 11336 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 1581 13787 1639 13793
rect 1581 13753 1593 13787
rect 1627 13784 1639 13787
rect 2130 13784 2136 13796
rect 1627 13756 2136 13784
rect 1627 13753 1639 13756
rect 1581 13747 1639 13753
rect 2130 13744 2136 13756
rect 2188 13744 2194 13796
rect 3142 13744 3148 13796
rect 3200 13784 3206 13796
rect 4706 13793 4712 13796
rect 4648 13787 4712 13793
rect 3200 13756 3648 13784
rect 3200 13744 3206 13756
rect 2406 13676 2412 13728
rect 2464 13716 2470 13728
rect 2961 13719 3019 13725
rect 2961 13716 2973 13719
rect 2464 13688 2973 13716
rect 2464 13676 2470 13688
rect 2961 13685 2973 13688
rect 3007 13685 3019 13719
rect 2961 13679 3019 13685
rect 3234 13676 3240 13728
rect 3292 13716 3298 13728
rect 3513 13719 3571 13725
rect 3513 13716 3525 13719
rect 3292 13688 3525 13716
rect 3292 13676 3298 13688
rect 3513 13685 3525 13688
rect 3559 13685 3571 13719
rect 3620 13716 3648 13756
rect 4648 13753 4660 13787
rect 4694 13753 4712 13787
rect 4648 13747 4712 13753
rect 4706 13744 4712 13747
rect 4764 13744 4770 13796
rect 9582 13784 9588 13796
rect 4816 13756 9588 13784
rect 4816 13716 4844 13756
rect 9582 13744 9588 13756
rect 9640 13744 9646 13796
rect 9769 13787 9827 13793
rect 9769 13753 9781 13787
rect 9815 13784 9827 13787
rect 10318 13784 10324 13796
rect 9815 13756 10324 13784
rect 9815 13753 9827 13756
rect 9769 13747 9827 13753
rect 10318 13744 10324 13756
rect 10376 13744 10382 13796
rect 10597 13787 10655 13793
rect 10597 13753 10609 13787
rect 10643 13784 10655 13787
rect 11164 13784 11192 13815
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 13538 13852 13544 13864
rect 13464 13824 13544 13852
rect 13078 13784 13084 13796
rect 10643 13756 11192 13784
rect 13039 13756 13084 13784
rect 10643 13753 10655 13756
rect 10597 13747 10655 13753
rect 13078 13744 13084 13756
rect 13136 13744 13142 13796
rect 5902 13716 5908 13728
rect 3620 13688 4844 13716
rect 5863 13688 5908 13716
rect 3513 13679 3571 13685
rect 5902 13676 5908 13688
rect 5960 13676 5966 13728
rect 6825 13719 6883 13725
rect 6825 13685 6837 13719
rect 6871 13716 6883 13719
rect 7558 13716 7564 13728
rect 6871 13688 7564 13716
rect 6871 13685 6883 13688
rect 6825 13679 6883 13685
rect 7558 13676 7564 13688
rect 7616 13676 7622 13728
rect 7653 13719 7711 13725
rect 7653 13685 7665 13719
rect 7699 13716 7711 13719
rect 8202 13716 8208 13728
rect 7699 13688 8208 13716
rect 7699 13685 7711 13688
rect 7653 13679 7711 13685
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 9309 13719 9367 13725
rect 9309 13685 9321 13719
rect 9355 13716 9367 13719
rect 9677 13719 9735 13725
rect 9677 13716 9689 13719
rect 9355 13688 9689 13716
rect 9355 13685 9367 13688
rect 9309 13679 9367 13685
rect 9677 13685 9689 13688
rect 9723 13716 9735 13719
rect 9858 13716 9864 13728
rect 9723 13688 9864 13716
rect 9723 13685 9735 13688
rect 9677 13679 9735 13685
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 10134 13716 10140 13728
rect 10095 13688 10140 13716
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 10410 13676 10416 13728
rect 10468 13716 10474 13728
rect 10689 13719 10747 13725
rect 10689 13716 10701 13719
rect 10468 13688 10701 13716
rect 10468 13676 10474 13688
rect 10689 13685 10701 13688
rect 10735 13716 10747 13719
rect 11425 13719 11483 13725
rect 11425 13716 11437 13719
rect 10735 13688 11437 13716
rect 10735 13685 10747 13688
rect 10689 13679 10747 13685
rect 11425 13685 11437 13688
rect 11471 13685 11483 13719
rect 11974 13716 11980 13728
rect 11935 13688 11980 13716
rect 11425 13679 11483 13685
rect 11974 13676 11980 13688
rect 12032 13676 12038 13728
rect 12069 13719 12127 13725
rect 12069 13685 12081 13719
rect 12115 13716 12127 13719
rect 12158 13716 12164 13728
rect 12115 13688 12164 13716
rect 12115 13685 12127 13688
rect 12069 13679 12127 13685
rect 12158 13676 12164 13688
rect 12216 13676 12222 13728
rect 12437 13719 12495 13725
rect 12437 13685 12449 13719
rect 12483 13716 12495 13719
rect 12802 13716 12808 13728
rect 12483 13688 12808 13716
rect 12483 13685 12495 13688
rect 12437 13679 12495 13685
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 12986 13716 12992 13728
rect 12947 13688 12992 13716
rect 12986 13676 12992 13688
rect 13044 13676 13050 13728
rect 13464 13725 13492 13824
rect 13538 13812 13544 13824
rect 13596 13812 13602 13864
rect 13814 13812 13820 13864
rect 13872 13852 13878 13864
rect 14366 13852 14372 13864
rect 13872 13824 14372 13852
rect 13872 13812 13878 13824
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 14921 13855 14979 13861
rect 14921 13821 14933 13855
rect 14967 13852 14979 13855
rect 16850 13852 16856 13864
rect 14967 13824 16856 13852
rect 14967 13821 14979 13824
rect 14921 13815 14979 13821
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 17402 13852 17408 13864
rect 17363 13824 17408 13852
rect 17402 13812 17408 13824
rect 17460 13852 17466 13864
rect 17773 13855 17831 13861
rect 17773 13852 17785 13855
rect 17460 13824 17785 13852
rect 17460 13812 17466 13824
rect 17773 13821 17785 13824
rect 17819 13821 17831 13855
rect 17773 13815 17831 13821
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18233 13855 18291 13861
rect 18233 13852 18245 13855
rect 18012 13824 18245 13852
rect 18012 13812 18018 13824
rect 18233 13821 18245 13824
rect 18279 13852 18291 13855
rect 18690 13852 18696 13864
rect 18279 13824 18696 13852
rect 18279 13821 18291 13824
rect 18233 13815 18291 13821
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 19058 13812 19064 13864
rect 19116 13852 19122 13864
rect 19153 13855 19211 13861
rect 19153 13852 19165 13855
rect 19116 13824 19165 13852
rect 19116 13812 19122 13824
rect 19153 13821 19165 13824
rect 19199 13821 19211 13855
rect 19702 13852 19708 13864
rect 19153 13815 19211 13821
rect 19306 13824 19708 13852
rect 14676 13787 14734 13793
rect 14676 13753 14688 13787
rect 14722 13784 14734 13787
rect 15102 13784 15108 13796
rect 14722 13756 15108 13784
rect 14722 13753 14734 13756
rect 14676 13747 14734 13753
rect 15102 13744 15108 13756
rect 15160 13744 15166 13796
rect 15194 13744 15200 13796
rect 15252 13784 15258 13796
rect 15350 13787 15408 13793
rect 15350 13784 15362 13787
rect 15252 13756 15362 13784
rect 15252 13744 15258 13756
rect 15350 13753 15362 13756
rect 15396 13784 15408 13787
rect 16114 13784 16120 13796
rect 15396 13756 16120 13784
rect 15396 13753 15408 13756
rect 15350 13747 15408 13753
rect 16114 13744 16120 13756
rect 16172 13744 16178 13796
rect 16761 13787 16819 13793
rect 16761 13753 16773 13787
rect 16807 13784 16819 13787
rect 17313 13787 17371 13793
rect 17313 13784 17325 13787
rect 16807 13756 17325 13784
rect 16807 13753 16819 13756
rect 16761 13747 16819 13753
rect 17313 13753 17325 13756
rect 17359 13753 17371 13787
rect 18322 13784 18328 13796
rect 17313 13747 17371 13753
rect 18156 13756 18328 13784
rect 13449 13719 13507 13725
rect 13449 13685 13461 13719
rect 13495 13685 13507 13719
rect 13449 13679 13507 13685
rect 13906 13676 13912 13728
rect 13964 13716 13970 13728
rect 15562 13716 15568 13728
rect 13964 13688 15568 13716
rect 13964 13676 13970 13688
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 18156 13716 18184 13756
rect 18322 13744 18328 13756
rect 18380 13744 18386 13796
rect 15712 13688 18184 13716
rect 15712 13676 15718 13688
rect 18782 13676 18788 13728
rect 18840 13716 18846 13728
rect 19061 13719 19119 13725
rect 19061 13716 19073 13719
rect 18840 13688 19073 13716
rect 18840 13676 18846 13688
rect 19061 13685 19073 13688
rect 19107 13716 19119 13719
rect 19306 13716 19334 13824
rect 19702 13812 19708 13824
rect 19760 13812 19766 13864
rect 20732 13852 20760 13951
rect 20809 13855 20867 13861
rect 20809 13852 20821 13855
rect 20732 13824 20821 13852
rect 20809 13821 20821 13824
rect 20855 13821 20867 13855
rect 21542 13852 21548 13864
rect 21503 13824 21548 13852
rect 20809 13815 20867 13821
rect 21542 13812 21548 13824
rect 21600 13812 21606 13864
rect 21358 13784 21364 13796
rect 21319 13756 21364 13784
rect 21358 13744 21364 13756
rect 21416 13744 21422 13796
rect 19107 13688 19334 13716
rect 19107 13685 19119 13688
rect 19061 13679 19119 13685
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 2130 13512 2136 13524
rect 2091 13484 2136 13512
rect 2130 13472 2136 13484
rect 2188 13472 2194 13524
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 2685 13515 2743 13521
rect 2685 13512 2697 13515
rect 2372 13484 2697 13512
rect 2372 13472 2378 13484
rect 2685 13481 2697 13484
rect 2731 13481 2743 13515
rect 3326 13512 3332 13524
rect 3287 13484 3332 13512
rect 2685 13475 2743 13481
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 3697 13515 3755 13521
rect 3697 13481 3709 13515
rect 3743 13512 3755 13515
rect 4338 13512 4344 13524
rect 3743 13484 4344 13512
rect 3743 13481 3755 13484
rect 3697 13475 3755 13481
rect 4338 13472 4344 13484
rect 4396 13472 4402 13524
rect 5258 13512 5264 13524
rect 5219 13484 5264 13512
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5902 13512 5908 13524
rect 5863 13484 5908 13512
rect 5902 13472 5908 13484
rect 5960 13472 5966 13524
rect 6365 13515 6423 13521
rect 6365 13481 6377 13515
rect 6411 13512 6423 13515
rect 6411 13484 7144 13512
rect 6411 13481 6423 13484
rect 6365 13475 6423 13481
rect 1581 13447 1639 13453
rect 1581 13413 1593 13447
rect 1627 13444 1639 13447
rect 3050 13444 3056 13456
rect 1627 13416 3056 13444
rect 1627 13413 1639 13416
rect 1581 13407 1639 13413
rect 3050 13404 3056 13416
rect 3108 13404 3114 13456
rect 3237 13447 3295 13453
rect 3237 13413 3249 13447
rect 3283 13444 3295 13447
rect 4890 13444 4896 13456
rect 3283 13416 4896 13444
rect 3283 13413 3295 13416
rect 3237 13407 3295 13413
rect 4890 13404 4896 13416
rect 4948 13404 4954 13456
rect 4982 13404 4988 13456
rect 5040 13444 5046 13456
rect 5350 13444 5356 13456
rect 5040 13416 5356 13444
rect 5040 13404 5046 13416
rect 5350 13404 5356 13416
rect 5408 13404 5414 13456
rect 6914 13404 6920 13456
rect 6972 13453 6978 13456
rect 6972 13447 7036 13453
rect 6972 13413 6990 13447
rect 7024 13413 7036 13447
rect 7116 13444 7144 13484
rect 7190 13472 7196 13524
rect 7248 13512 7254 13524
rect 8205 13515 8263 13521
rect 8205 13512 8217 13515
rect 7248 13484 8217 13512
rect 7248 13472 7254 13484
rect 8205 13481 8217 13484
rect 8251 13481 8263 13515
rect 8570 13512 8576 13524
rect 8483 13484 8576 13512
rect 8205 13475 8263 13481
rect 8570 13472 8576 13484
rect 8628 13512 8634 13524
rect 9030 13512 9036 13524
rect 8628 13484 9036 13512
rect 8628 13472 8634 13484
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 9309 13515 9367 13521
rect 9309 13481 9321 13515
rect 9355 13481 9367 13515
rect 9309 13475 9367 13481
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 10134 13512 10140 13524
rect 9723 13484 10140 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 7116 13416 7613 13444
rect 6972 13407 7036 13413
rect 6972 13404 6978 13407
rect 1946 13376 1952 13388
rect 1907 13348 1952 13376
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 2317 13379 2375 13385
rect 2317 13345 2329 13379
rect 2363 13376 2375 13379
rect 2406 13376 2412 13388
rect 2363 13348 2412 13376
rect 2363 13345 2375 13348
rect 2317 13339 2375 13345
rect 2406 13336 2412 13348
rect 2464 13336 2470 13388
rect 2590 13376 2596 13388
rect 2551 13348 2596 13376
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 2866 13376 2872 13388
rect 2827 13348 2872 13376
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 2958 13336 2964 13388
rect 3016 13376 3022 13388
rect 3881 13379 3939 13385
rect 3881 13376 3893 13379
rect 3016 13348 3893 13376
rect 3016 13336 3022 13348
rect 3881 13345 3893 13348
rect 3927 13376 3939 13379
rect 3970 13376 3976 13388
rect 3927 13348 3976 13376
rect 3927 13345 3939 13348
rect 3881 13339 3939 13345
rect 3970 13336 3976 13348
rect 4028 13336 4034 13388
rect 4148 13379 4206 13385
rect 4148 13345 4160 13379
rect 4194 13376 4206 13379
rect 4430 13376 4436 13388
rect 4194 13348 4436 13376
rect 4194 13345 4206 13348
rect 4148 13339 4206 13345
rect 4430 13336 4436 13348
rect 4488 13376 4494 13388
rect 4488 13348 5672 13376
rect 4488 13336 4494 13348
rect 2424 13308 2452 13336
rect 3145 13311 3203 13317
rect 2424 13280 2820 13308
rect 1762 13200 1768 13252
rect 1820 13240 1826 13252
rect 2409 13243 2467 13249
rect 2409 13240 2421 13243
rect 1820 13212 2421 13240
rect 1820 13200 1826 13212
rect 2409 13209 2421 13212
rect 2455 13209 2467 13243
rect 2409 13203 2467 13209
rect 1394 13132 1400 13184
rect 1452 13172 1458 13184
rect 1489 13175 1547 13181
rect 1489 13172 1501 13175
rect 1452 13144 1501 13172
rect 1452 13132 1458 13144
rect 1489 13141 1501 13144
rect 1535 13141 1547 13175
rect 1854 13172 1860 13184
rect 1815 13144 1860 13172
rect 1489 13135 1547 13141
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 2792 13172 2820 13280
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 3234 13308 3240 13320
rect 3191 13280 3240 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 5644 13240 5672 13348
rect 5810 13336 5816 13388
rect 5868 13376 5874 13388
rect 6178 13376 6184 13388
rect 5868 13348 6184 13376
rect 5868 13336 5874 13348
rect 6178 13336 6184 13348
rect 6236 13376 6242 13388
rect 6273 13379 6331 13385
rect 6273 13376 6285 13379
rect 6236 13348 6285 13376
rect 6236 13336 6242 13348
rect 6273 13345 6285 13348
rect 6319 13345 6331 13379
rect 6273 13339 6331 13345
rect 6733 13379 6791 13385
rect 6733 13345 6745 13379
rect 6779 13376 6791 13379
rect 6822 13376 6828 13388
rect 6779 13348 6828 13376
rect 6779 13345 6791 13348
rect 6733 13339 6791 13345
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 7585 13376 7613 13416
rect 7650 13404 7656 13456
rect 7708 13444 7714 13456
rect 7708 13416 8800 13444
rect 7708 13404 7714 13416
rect 8386 13376 8392 13388
rect 7585 13348 8392 13376
rect 8386 13336 8392 13348
rect 8444 13336 8450 13388
rect 5721 13311 5779 13317
rect 5721 13277 5733 13311
rect 5767 13308 5779 13311
rect 5902 13308 5908 13320
rect 5767 13280 5908 13308
rect 5767 13277 5779 13280
rect 5721 13271 5779 13277
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 8772 13317 8800 13416
rect 8846 13404 8852 13456
rect 8904 13444 8910 13456
rect 9324 13444 9352 13475
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 10413 13515 10471 13521
rect 10413 13481 10425 13515
rect 10459 13512 10471 13515
rect 11790 13512 11796 13524
rect 10459 13484 11796 13512
rect 10459 13481 10471 13484
rect 10413 13475 10471 13481
rect 11790 13472 11796 13484
rect 11848 13472 11854 13524
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 11977 13515 12035 13521
rect 11977 13512 11989 13515
rect 11940 13484 11989 13512
rect 11940 13472 11946 13484
rect 11977 13481 11989 13484
rect 12023 13481 12035 13515
rect 11977 13475 12035 13481
rect 12069 13515 12127 13521
rect 12069 13481 12081 13515
rect 12115 13512 12127 13515
rect 12158 13512 12164 13524
rect 12115 13484 12164 13512
rect 12115 13481 12127 13484
rect 12069 13475 12127 13481
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 12342 13472 12348 13524
rect 12400 13512 12406 13524
rect 12529 13515 12587 13521
rect 12529 13512 12541 13515
rect 12400 13484 12541 13512
rect 12400 13472 12406 13484
rect 12529 13481 12541 13484
rect 12575 13512 12587 13515
rect 12897 13515 12955 13521
rect 12897 13512 12909 13515
rect 12575 13484 12909 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 12897 13481 12909 13484
rect 12943 13481 12955 13515
rect 12897 13475 12955 13481
rect 12986 13472 12992 13524
rect 13044 13512 13050 13524
rect 13449 13515 13507 13521
rect 13449 13512 13461 13515
rect 13044 13484 13461 13512
rect 13044 13472 13050 13484
rect 13449 13481 13461 13484
rect 13495 13481 13507 13515
rect 13449 13475 13507 13481
rect 13630 13472 13636 13524
rect 13688 13512 13694 13524
rect 13817 13515 13875 13521
rect 13817 13512 13829 13515
rect 13688 13484 13829 13512
rect 13688 13472 13694 13484
rect 13817 13481 13829 13484
rect 13863 13481 13875 13515
rect 14550 13512 14556 13524
rect 14511 13484 14556 13512
rect 13817 13475 13875 13481
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 15289 13515 15347 13521
rect 15289 13512 15301 13515
rect 14651 13484 15301 13512
rect 8904 13416 9352 13444
rect 9769 13447 9827 13453
rect 8904 13404 8910 13416
rect 9769 13413 9781 13447
rect 9815 13444 9827 13447
rect 11054 13444 11060 13456
rect 9815 13416 11060 13444
rect 9815 13413 9827 13416
rect 9769 13407 9827 13413
rect 11054 13404 11060 13416
rect 11112 13404 11118 13456
rect 13538 13404 13544 13456
rect 13596 13444 13602 13456
rect 14651 13444 14679 13484
rect 15289 13481 15301 13484
rect 15335 13481 15347 13515
rect 15289 13475 15347 13481
rect 15749 13515 15807 13521
rect 15749 13481 15761 13515
rect 15795 13481 15807 13515
rect 15749 13475 15807 13481
rect 15841 13515 15899 13521
rect 15841 13481 15853 13515
rect 15887 13512 15899 13515
rect 15930 13512 15936 13524
rect 15887 13484 15936 13512
rect 15887 13481 15899 13484
rect 15841 13475 15899 13481
rect 13596 13416 14136 13444
rect 13596 13404 13602 13416
rect 9217 13379 9275 13385
rect 9217 13345 9229 13379
rect 9263 13376 9275 13379
rect 9306 13376 9312 13388
rect 9263 13348 9312 13376
rect 9263 13345 9275 13348
rect 9217 13339 9275 13345
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13277 8723 13311
rect 8665 13271 8723 13277
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 6472 13240 6500 13271
rect 6638 13240 6644 13252
rect 5644 13212 6644 13240
rect 6638 13200 6644 13212
rect 6696 13200 6702 13252
rect 8570 13240 8576 13252
rect 8036 13212 8576 13240
rect 5534 13172 5540 13184
rect 2792 13144 5540 13172
rect 5534 13132 5540 13144
rect 5592 13172 5598 13184
rect 8036 13172 8064 13212
rect 8570 13200 8576 13212
rect 8628 13200 8634 13252
rect 8680 13240 8708 13271
rect 9232 13240 9260 13339
rect 9306 13336 9312 13348
rect 9364 13336 9370 13388
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 10870 13385 10876 13388
rect 10597 13379 10655 13385
rect 10597 13376 10609 13379
rect 9456 13348 10609 13376
rect 9456 13336 9462 13348
rect 10597 13345 10609 13348
rect 10643 13345 10655 13379
rect 10864 13376 10876 13385
rect 10783 13348 10876 13376
rect 10597 13339 10655 13345
rect 10864 13339 10876 13348
rect 10928 13376 10934 13388
rect 12437 13379 12495 13385
rect 10928 13348 11652 13376
rect 10870 13336 10876 13339
rect 10928 13336 10934 13348
rect 9490 13308 9496 13320
rect 9451 13280 9496 13308
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 11624 13308 11652 13348
rect 12437 13345 12449 13379
rect 12483 13376 12495 13379
rect 12710 13376 12716 13388
rect 12483 13348 12716 13376
rect 12483 13345 12495 13348
rect 12437 13339 12495 13345
rect 12710 13336 12716 13348
rect 12768 13336 12774 13388
rect 14108 13317 14136 13416
rect 14568 13416 14679 13444
rect 14568 13388 14596 13416
rect 15010 13404 15016 13456
rect 15068 13444 15074 13456
rect 15381 13447 15439 13453
rect 15381 13444 15393 13447
rect 15068 13416 15393 13444
rect 15068 13404 15074 13416
rect 15381 13413 15393 13416
rect 15427 13413 15439 13447
rect 15764 13444 15792 13475
rect 15930 13472 15936 13484
rect 15988 13472 15994 13524
rect 16206 13512 16212 13524
rect 16167 13484 16212 13512
rect 16206 13472 16212 13484
rect 16264 13472 16270 13524
rect 16850 13512 16856 13524
rect 16811 13484 16856 13512
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 17313 13515 17371 13521
rect 17313 13481 17325 13515
rect 17359 13512 17371 13515
rect 17865 13515 17923 13521
rect 17865 13512 17877 13515
rect 17359 13484 17877 13512
rect 17359 13481 17371 13484
rect 17313 13475 17371 13481
rect 17865 13481 17877 13484
rect 17911 13481 17923 13515
rect 17865 13475 17923 13481
rect 18322 13472 18328 13524
rect 18380 13512 18386 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 18380 13484 18889 13512
rect 18380 13472 18386 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 16022 13444 16028 13456
rect 15764 13416 16028 13444
rect 15381 13407 15439 13413
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 16114 13404 16120 13456
rect 16172 13444 16178 13456
rect 18782 13444 18788 13456
rect 16172 13416 16712 13444
rect 18743 13416 18788 13444
rect 16172 13404 16178 13416
rect 14366 13376 14372 13388
rect 14327 13348 14372 13376
rect 14366 13336 14372 13348
rect 14424 13336 14430 13388
rect 14550 13336 14556 13388
rect 14608 13336 14614 13388
rect 16684 13385 16712 13416
rect 18782 13404 18788 13416
rect 18840 13404 18846 13456
rect 18892 13444 18920 13475
rect 19426 13472 19432 13524
rect 19484 13512 19490 13524
rect 20349 13515 20407 13521
rect 20349 13512 20361 13515
rect 19484 13484 20361 13512
rect 19484 13472 19490 13484
rect 20349 13481 20361 13484
rect 20395 13481 20407 13515
rect 20349 13475 20407 13481
rect 20993 13515 21051 13521
rect 20993 13481 21005 13515
rect 21039 13512 21051 13515
rect 21039 13484 21404 13512
rect 21039 13481 21051 13484
rect 20993 13475 21051 13481
rect 20438 13444 20444 13456
rect 18892 13416 20444 13444
rect 20438 13404 20444 13416
rect 20496 13404 20502 13456
rect 21376 13453 21404 13484
rect 21361 13447 21419 13453
rect 21361 13413 21373 13447
rect 21407 13413 21419 13447
rect 21361 13407 21419 13413
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 14844 13348 16313 13376
rect 14844 13320 14872 13348
rect 16301 13345 16313 13348
rect 16347 13345 16359 13379
rect 16301 13339 16359 13345
rect 16669 13379 16727 13385
rect 16669 13345 16681 13379
rect 16715 13345 16727 13379
rect 16669 13339 16727 13345
rect 17405 13379 17463 13385
rect 17405 13345 17417 13379
rect 17451 13376 17463 13379
rect 17862 13376 17868 13388
rect 17451 13348 17868 13376
rect 17451 13345 17463 13348
rect 17405 13339 17463 13345
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18138 13336 18144 13388
rect 18196 13376 18202 13388
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 18196 13348 18245 13376
rect 18196 13336 18202 13348
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 18690 13336 18696 13388
rect 18748 13376 18754 13388
rect 19061 13379 19119 13385
rect 19061 13376 19073 13379
rect 18748 13348 19073 13376
rect 18748 13336 18754 13348
rect 19061 13345 19073 13348
rect 19107 13345 19119 13379
rect 19061 13339 19119 13345
rect 20254 13336 20260 13388
rect 20312 13376 20318 13388
rect 20533 13379 20591 13385
rect 20533 13376 20545 13379
rect 20312 13348 20545 13376
rect 20312 13336 20318 13348
rect 20533 13345 20545 13348
rect 20579 13345 20591 13379
rect 20533 13339 20591 13345
rect 20809 13379 20867 13385
rect 20809 13345 20821 13379
rect 20855 13345 20867 13379
rect 21542 13376 21548 13388
rect 21503 13348 21548 13376
rect 20809 13339 20867 13345
rect 12621 13311 12679 13317
rect 12621 13308 12633 13311
rect 11624 13280 12633 13308
rect 12621 13277 12633 13280
rect 12667 13277 12679 13311
rect 12621 13271 12679 13277
rect 13909 13311 13967 13317
rect 13909 13277 13921 13311
rect 13955 13277 13967 13311
rect 13909 13271 13967 13277
rect 14093 13311 14151 13317
rect 14093 13277 14105 13311
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 14737 13311 14795 13317
rect 14737 13277 14749 13311
rect 14783 13308 14795 13311
rect 14826 13308 14832 13320
rect 14783 13280 14832 13308
rect 14783 13277 14795 13280
rect 14737 13271 14795 13277
rect 8680 13212 9260 13240
rect 9309 13243 9367 13249
rect 9309 13209 9321 13243
rect 9355 13240 9367 13243
rect 10137 13243 10195 13249
rect 9355 13212 9674 13240
rect 9355 13209 9367 13212
rect 9309 13203 9367 13209
rect 5592 13144 8064 13172
rect 8113 13175 8171 13181
rect 5592 13132 5598 13144
rect 8113 13141 8125 13175
rect 8159 13172 8171 13175
rect 8294 13172 8300 13184
rect 8159 13144 8300 13172
rect 8159 13141 8171 13144
rect 8113 13135 8171 13141
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 9646 13172 9674 13212
rect 10137 13209 10149 13243
rect 10183 13240 10195 13243
rect 10226 13240 10232 13252
rect 10183 13212 10232 13240
rect 10183 13209 10195 13212
rect 10137 13203 10195 13209
rect 10226 13200 10232 13212
rect 10284 13200 10290 13252
rect 13262 13240 13268 13252
rect 11624 13212 13268 13240
rect 11624 13172 11652 13212
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 13924 13240 13952 13271
rect 14826 13268 14832 13280
rect 14884 13268 14890 13320
rect 15194 13308 15200 13320
rect 15155 13280 15200 13308
rect 15194 13268 15200 13280
rect 15252 13268 15258 13320
rect 16482 13308 16488 13320
rect 16443 13280 16488 13308
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 17218 13308 17224 13320
rect 17179 13280 17224 13308
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 17770 13268 17776 13320
rect 17828 13308 17834 13320
rect 18325 13311 18383 13317
rect 18325 13308 18337 13311
rect 17828 13280 18337 13308
rect 17828 13268 17834 13280
rect 18325 13277 18337 13280
rect 18371 13277 18383 13311
rect 18325 13271 18383 13277
rect 18509 13311 18567 13317
rect 18509 13277 18521 13311
rect 18555 13308 18567 13311
rect 18874 13308 18880 13320
rect 18555 13280 18880 13308
rect 18555 13277 18567 13280
rect 18509 13271 18567 13277
rect 18874 13268 18880 13280
rect 18932 13268 18938 13320
rect 15746 13240 15752 13252
rect 13924 13212 15752 13240
rect 15746 13200 15752 13212
rect 15804 13200 15810 13252
rect 17402 13200 17408 13252
rect 17460 13240 17466 13252
rect 19245 13243 19303 13249
rect 19245 13240 19257 13243
rect 17460 13212 19257 13240
rect 17460 13200 17466 13212
rect 19245 13209 19257 13212
rect 19291 13209 19303 13243
rect 19245 13203 19303 13209
rect 9646 13144 11652 13172
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 12250 13172 12256 13184
rect 11756 13144 12256 13172
rect 11756 13132 11762 13144
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 12618 13132 12624 13184
rect 12676 13172 12682 13184
rect 14921 13175 14979 13181
rect 14921 13172 14933 13175
rect 12676 13144 14933 13172
rect 12676 13132 12682 13144
rect 14921 13141 14933 13144
rect 14967 13172 14979 13175
rect 16206 13172 16212 13184
rect 14967 13144 16212 13172
rect 14967 13141 14979 13144
rect 14921 13135 14979 13141
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 17773 13175 17831 13181
rect 17773 13141 17785 13175
rect 17819 13172 17831 13175
rect 18046 13172 18052 13184
rect 17819 13144 18052 13172
rect 17819 13141 17831 13144
rect 17773 13135 17831 13141
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 20717 13175 20775 13181
rect 20717 13141 20729 13175
rect 20763 13172 20775 13175
rect 20824 13172 20852 13339
rect 21542 13336 21548 13348
rect 21600 13336 21606 13388
rect 20898 13172 20904 13184
rect 20763 13144 20904 13172
rect 20763 13141 20775 13144
rect 20717 13135 20775 13141
rect 20898 13132 20904 13144
rect 20956 13132 20962 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1946 12968 1952 12980
rect 1907 12940 1952 12968
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 3421 12971 3479 12977
rect 3421 12937 3433 12971
rect 3467 12968 3479 12971
rect 4338 12968 4344 12980
rect 3467 12940 4344 12968
rect 3467 12937 3479 12940
rect 3421 12931 3479 12937
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 5813 12971 5871 12977
rect 5813 12968 5825 12971
rect 5776 12940 5825 12968
rect 5776 12928 5782 12940
rect 5813 12937 5825 12940
rect 5859 12937 5871 12971
rect 6454 12968 6460 12980
rect 6415 12940 6460 12968
rect 5813 12931 5871 12937
rect 6454 12928 6460 12940
rect 6512 12928 6518 12980
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 7745 12971 7803 12977
rect 7745 12968 7757 12971
rect 7064 12940 7757 12968
rect 7064 12928 7070 12940
rect 7745 12937 7757 12940
rect 7791 12937 7803 12971
rect 8662 12968 8668 12980
rect 7745 12931 7803 12937
rect 7852 12940 8668 12968
rect 7852 12900 7880 12940
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 9030 12928 9036 12980
rect 9088 12968 9094 12980
rect 9493 12971 9551 12977
rect 9493 12968 9505 12971
rect 9088 12940 9505 12968
rect 9088 12928 9094 12940
rect 9493 12937 9505 12940
rect 9539 12937 9551 12971
rect 9493 12931 9551 12937
rect 9858 12928 9864 12980
rect 9916 12968 9922 12980
rect 10686 12968 10692 12980
rect 9916 12940 10692 12968
rect 9916 12928 9922 12940
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 11517 12971 11575 12977
rect 11517 12937 11529 12971
rect 11563 12968 11575 12971
rect 11974 12968 11980 12980
rect 11563 12940 11980 12968
rect 11563 12937 11575 12940
rect 11517 12931 11575 12937
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 13817 12971 13875 12977
rect 13817 12937 13829 12971
rect 13863 12968 13875 12971
rect 13998 12968 14004 12980
rect 13863 12940 14004 12968
rect 13863 12937 13875 12940
rect 13817 12931 13875 12937
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 14093 12971 14151 12977
rect 14093 12937 14105 12971
rect 14139 12937 14151 12971
rect 15746 12968 15752 12980
rect 15707 12940 15752 12968
rect 14093 12931 14151 12937
rect 5736 12872 7880 12900
rect 5736 12844 5764 12872
rect 9582 12860 9588 12912
rect 9640 12900 9646 12912
rect 9640 12872 11192 12900
rect 9640 12860 9646 12872
rect 3789 12835 3847 12841
rect 3789 12801 3801 12835
rect 3835 12832 3847 12835
rect 4062 12832 4068 12844
rect 3835 12804 4068 12832
rect 3835 12801 3847 12804
rect 3789 12795 3847 12801
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 5718 12792 5724 12844
rect 5776 12792 5782 12844
rect 5810 12792 5816 12844
rect 5868 12832 5874 12844
rect 5997 12835 6055 12841
rect 5997 12832 6009 12835
rect 5868 12804 6009 12832
rect 5868 12792 5874 12804
rect 5997 12801 6009 12804
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6638 12792 6644 12844
rect 6696 12832 6702 12844
rect 7009 12835 7067 12841
rect 7009 12832 7021 12835
rect 6696 12804 7021 12832
rect 6696 12792 6702 12804
rect 7009 12801 7021 12804
rect 7055 12801 7067 12835
rect 7558 12832 7564 12844
rect 7519 12804 7564 12832
rect 7009 12795 7067 12801
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 10192 12804 10609 12832
rect 10192 12792 10198 12804
rect 10597 12801 10609 12804
rect 10643 12801 10655 12835
rect 10870 12832 10876 12844
rect 10831 12804 10876 12832
rect 10597 12795 10655 12801
rect 1762 12764 1768 12776
rect 1723 12736 1768 12764
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 2041 12767 2099 12773
rect 2041 12733 2053 12767
rect 2087 12764 2099 12767
rect 2087 12736 2728 12764
rect 2087 12733 2099 12736
rect 2041 12727 2099 12733
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12665 1639 12699
rect 1581 12659 1639 12665
rect 1486 12628 1492 12640
rect 1447 12600 1492 12628
rect 1486 12588 1492 12600
rect 1544 12588 1550 12640
rect 1596 12628 1624 12659
rect 1946 12656 1952 12708
rect 2004 12696 2010 12708
rect 2286 12699 2344 12705
rect 2286 12696 2298 12699
rect 2004 12668 2298 12696
rect 2004 12656 2010 12668
rect 2286 12665 2298 12668
rect 2332 12665 2344 12699
rect 2700 12696 2728 12736
rect 2774 12724 2780 12776
rect 2832 12764 2838 12776
rect 3881 12767 3939 12773
rect 3881 12764 3893 12767
rect 2832 12736 3893 12764
rect 2832 12724 2838 12736
rect 3881 12733 3893 12736
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 3970 12724 3976 12776
rect 4028 12764 4034 12776
rect 4433 12767 4491 12773
rect 4433 12764 4445 12767
rect 4028 12736 4445 12764
rect 4028 12724 4034 12736
rect 4433 12733 4445 12736
rect 4479 12733 4491 12767
rect 4433 12727 4491 12733
rect 5074 12724 5080 12776
rect 5132 12764 5138 12776
rect 5902 12764 5908 12776
rect 5132 12736 5908 12764
rect 5132 12724 5138 12736
rect 5902 12724 5908 12736
rect 5960 12764 5966 12776
rect 6089 12767 6147 12773
rect 6089 12764 6101 12767
rect 5960 12736 6101 12764
rect 5960 12724 5966 12736
rect 6089 12733 6101 12736
rect 6135 12733 6147 12767
rect 6089 12727 6147 12733
rect 6178 12724 6184 12776
rect 6236 12764 6242 12776
rect 7576 12764 7604 12792
rect 6236 12736 7604 12764
rect 6236 12724 6242 12736
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 7929 12767 7987 12773
rect 7929 12764 7941 12767
rect 7892 12736 7941 12764
rect 7892 12724 7898 12736
rect 7929 12733 7941 12736
rect 7975 12733 7987 12767
rect 7929 12727 7987 12733
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 9134 12767 9192 12773
rect 9134 12764 9146 12767
rect 8352 12736 9146 12764
rect 8352 12724 8358 12736
rect 9134 12733 9146 12736
rect 9180 12733 9192 12767
rect 9134 12727 9192 12733
rect 9401 12767 9459 12773
rect 9401 12733 9413 12767
rect 9447 12764 9459 12767
rect 9490 12764 9496 12776
rect 9447 12736 9496 12764
rect 9447 12733 9459 12736
rect 9401 12727 9459 12733
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 9582 12724 9588 12776
rect 9640 12764 9646 12776
rect 10321 12767 10379 12773
rect 9640 12736 10180 12764
rect 9640 12724 9646 12736
rect 2866 12696 2872 12708
rect 2700 12668 2872 12696
rect 2286 12659 2344 12665
rect 2866 12656 2872 12668
rect 2924 12656 2930 12708
rect 3234 12656 3240 12708
rect 3292 12696 3298 12708
rect 4700 12699 4758 12705
rect 4700 12696 4712 12699
rect 3292 12668 4712 12696
rect 3292 12656 3298 12668
rect 4700 12665 4712 12668
rect 4746 12696 4758 12699
rect 4982 12696 4988 12708
rect 4746 12668 4988 12696
rect 4746 12665 4758 12668
rect 4700 12659 4758 12665
rect 4982 12656 4988 12668
rect 5040 12656 5046 12708
rect 6825 12699 6883 12705
rect 6825 12665 6837 12699
rect 6871 12696 6883 12699
rect 7098 12696 7104 12708
rect 6871 12668 7104 12696
rect 6871 12665 6883 12668
rect 6825 12659 6883 12665
rect 7098 12656 7104 12668
rect 7156 12656 7162 12708
rect 7742 12656 7748 12708
rect 7800 12696 7806 12708
rect 9306 12696 9312 12708
rect 7800 12668 9312 12696
rect 7800 12656 7806 12668
rect 9306 12656 9312 12668
rect 9364 12696 9370 12708
rect 10152 12705 10180 12736
rect 10321 12733 10333 12767
rect 10367 12764 10379 12767
rect 10502 12764 10508 12776
rect 10367 12736 10508 12764
rect 10367 12733 10379 12736
rect 10321 12727 10379 12733
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 10612 12764 10640 12795
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11164 12773 11192 12872
rect 11238 12792 11244 12844
rect 11296 12832 11302 12844
rect 11698 12832 11704 12844
rect 11296 12804 11704 12832
rect 11296 12792 11302 12804
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 12768 12804 13185 12832
rect 12768 12792 12774 12804
rect 13173 12801 13185 12804
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 14108 12832 14136 12931
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 17770 12968 17776 12980
rect 17731 12940 17776 12968
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 17862 12928 17868 12980
rect 17920 12968 17926 12980
rect 19337 12971 19395 12977
rect 19337 12968 19349 12971
rect 17920 12940 19349 12968
rect 17920 12928 17926 12940
rect 19337 12937 19349 12940
rect 19383 12937 19395 12971
rect 19337 12931 19395 12937
rect 20993 12971 21051 12977
rect 20993 12937 21005 12971
rect 21039 12968 21051 12971
rect 21358 12968 21364 12980
rect 21039 12940 21364 12968
rect 21039 12937 21051 12940
rect 20993 12931 21051 12937
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 15194 12860 15200 12912
rect 15252 12900 15258 12912
rect 16482 12900 16488 12912
rect 15252 12872 16488 12900
rect 15252 12860 15258 12872
rect 13688 12804 14136 12832
rect 14737 12835 14795 12841
rect 13688 12792 13694 12804
rect 14737 12801 14749 12835
rect 14783 12832 14795 12835
rect 14826 12832 14832 12844
rect 14783 12804 14832 12832
rect 14783 12801 14795 12804
rect 14737 12795 14795 12801
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 15580 12841 15608 12872
rect 16482 12860 16488 12872
rect 16540 12860 16546 12912
rect 18874 12860 18880 12912
rect 18932 12900 18938 12912
rect 19245 12903 19303 12909
rect 19245 12900 19257 12903
rect 18932 12872 19257 12900
rect 18932 12860 18938 12872
rect 19245 12869 19257 12872
rect 19291 12869 19303 12903
rect 19245 12863 19303 12869
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12801 15623 12835
rect 15565 12795 15623 12801
rect 16022 12792 16028 12844
rect 16080 12832 16086 12844
rect 16209 12835 16267 12841
rect 16209 12832 16221 12835
rect 16080 12804 16221 12832
rect 16080 12792 16086 12804
rect 16209 12801 16221 12804
rect 16255 12801 16267 12835
rect 16390 12832 16396 12844
rect 16351 12804 16396 12832
rect 16209 12795 16267 12801
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 19260 12832 19288 12863
rect 19889 12835 19947 12841
rect 19889 12832 19901 12835
rect 17267 12804 18000 12832
rect 19260 12804 19901 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 11057 12767 11115 12773
rect 11057 12764 11069 12767
rect 10612 12736 11069 12764
rect 11057 12733 11069 12736
rect 11103 12733 11115 12767
rect 11057 12727 11115 12733
rect 11149 12767 11207 12773
rect 11149 12733 11161 12767
rect 11195 12733 11207 12767
rect 11149 12727 11207 12733
rect 11808 12736 16804 12764
rect 9861 12699 9919 12705
rect 9861 12696 9873 12699
rect 9364 12668 9873 12696
rect 9364 12656 9370 12668
rect 9861 12665 9873 12668
rect 9907 12665 9919 12699
rect 9861 12659 9919 12665
rect 10137 12699 10195 12705
rect 10137 12665 10149 12699
rect 10183 12696 10195 12699
rect 11808 12696 11836 12736
rect 10183 12668 11836 12696
rect 10183 12665 10195 12668
rect 10137 12659 10195 12665
rect 11882 12656 11888 12708
rect 11940 12705 11946 12708
rect 11940 12699 12004 12705
rect 11940 12665 11958 12699
rect 11992 12665 12004 12699
rect 15289 12699 15347 12705
rect 15289 12696 15301 12699
rect 11940 12659 12004 12665
rect 13924 12668 15301 12696
rect 11940 12656 11946 12659
rect 13924 12640 13952 12668
rect 15289 12665 15301 12668
rect 15335 12665 15347 12699
rect 15289 12659 15347 12665
rect 15381 12699 15439 12705
rect 15381 12665 15393 12699
rect 15427 12696 15439 12699
rect 16022 12696 16028 12708
rect 15427 12668 16028 12696
rect 15427 12665 15439 12668
rect 15381 12659 15439 12665
rect 16022 12656 16028 12668
rect 16080 12656 16086 12708
rect 16117 12699 16175 12705
rect 16117 12665 16129 12699
rect 16163 12696 16175 12699
rect 16390 12696 16396 12708
rect 16163 12668 16396 12696
rect 16163 12665 16175 12668
rect 16117 12659 16175 12665
rect 16390 12656 16396 12668
rect 16448 12656 16454 12708
rect 2958 12628 2964 12640
rect 1596 12600 2964 12628
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 3970 12588 3976 12640
rect 4028 12628 4034 12640
rect 4338 12628 4344 12640
rect 4028 12600 4073 12628
rect 4299 12600 4344 12628
rect 4028 12588 4034 12600
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 4890 12588 4896 12640
rect 4948 12628 4954 12640
rect 5258 12628 5264 12640
rect 4948 12600 5264 12628
rect 4948 12588 4954 12600
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5534 12588 5540 12640
rect 5592 12628 5598 12640
rect 6178 12628 6184 12640
rect 5592 12600 6184 12628
rect 5592 12588 5598 12600
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 6638 12588 6644 12640
rect 6696 12628 6702 12640
rect 6917 12631 6975 12637
rect 6917 12628 6929 12631
rect 6696 12600 6929 12628
rect 6696 12588 6702 12600
rect 6917 12597 6929 12600
rect 6963 12628 6975 12631
rect 7285 12631 7343 12637
rect 7285 12628 7297 12631
rect 6963 12600 7297 12628
rect 6963 12597 6975 12600
rect 6917 12591 6975 12597
rect 7285 12597 7297 12600
rect 7331 12597 7343 12631
rect 7285 12591 7343 12597
rect 8021 12631 8079 12637
rect 8021 12597 8033 12631
rect 8067 12628 8079 12631
rect 8202 12628 8208 12640
rect 8067 12600 8208 12628
rect 8067 12597 8079 12600
rect 8021 12591 8079 12597
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 8570 12588 8576 12640
rect 8628 12628 8634 12640
rect 9677 12631 9735 12637
rect 9677 12628 9689 12631
rect 8628 12600 9689 12628
rect 8628 12588 8634 12600
rect 9677 12597 9689 12600
rect 9723 12628 9735 12631
rect 10962 12628 10968 12640
rect 9723 12600 10968 12628
rect 9723 12597 9735 12600
rect 9677 12591 9735 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 13078 12628 13084 12640
rect 13039 12600 13084 12628
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 13262 12588 13268 12640
rect 13320 12628 13326 12640
rect 13630 12628 13636 12640
rect 13320 12600 13636 12628
rect 13320 12588 13326 12600
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 13906 12628 13912 12640
rect 13867 12600 13912 12628
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 16776 12637 16804 12736
rect 16942 12724 16948 12776
rect 17000 12764 17006 12776
rect 17402 12764 17408 12776
rect 17000 12736 17408 12764
rect 17000 12724 17006 12736
rect 17402 12724 17408 12736
rect 17460 12724 17466 12776
rect 17865 12767 17923 12773
rect 17865 12733 17877 12767
rect 17911 12733 17923 12767
rect 17972 12764 18000 12804
rect 19889 12801 19901 12804
rect 19935 12801 19947 12835
rect 21542 12832 21548 12844
rect 21503 12804 21548 12832
rect 19889 12795 19947 12801
rect 21542 12792 21548 12804
rect 21600 12792 21606 12844
rect 18121 12767 18179 12773
rect 18121 12764 18133 12767
rect 17972 12736 18133 12764
rect 17865 12727 17923 12733
rect 18121 12733 18133 12736
rect 18167 12764 18179 12767
rect 18874 12764 18880 12776
rect 18167 12736 18880 12764
rect 18167 12733 18179 12736
rect 18121 12727 18179 12733
rect 16850 12656 16856 12708
rect 16908 12696 16914 12708
rect 17494 12696 17500 12708
rect 16908 12668 17500 12696
rect 16908 12656 16914 12668
rect 17494 12656 17500 12668
rect 17552 12696 17558 12708
rect 17880 12696 17908 12727
rect 18874 12724 18880 12736
rect 18932 12764 18938 12776
rect 19058 12764 19064 12776
rect 18932 12736 19064 12764
rect 18932 12724 18938 12736
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 20162 12724 20168 12776
rect 20220 12764 20226 12776
rect 20809 12767 20867 12773
rect 20809 12764 20821 12767
rect 20220 12736 20821 12764
rect 20220 12724 20226 12736
rect 20809 12733 20821 12736
rect 20855 12733 20867 12767
rect 20809 12727 20867 12733
rect 17552 12668 17908 12696
rect 17552 12656 17558 12668
rect 19426 12656 19432 12708
rect 19484 12696 19490 12708
rect 19797 12699 19855 12705
rect 19797 12696 19809 12699
rect 19484 12668 19809 12696
rect 19484 12656 19490 12668
rect 19797 12665 19809 12668
rect 19843 12665 19855 12699
rect 19797 12659 19855 12665
rect 20714 12656 20720 12708
rect 20772 12696 20778 12708
rect 21361 12699 21419 12705
rect 21361 12696 21373 12699
rect 20772 12668 21373 12696
rect 20772 12656 20778 12668
rect 21361 12665 21373 12668
rect 21407 12665 21419 12699
rect 21361 12659 21419 12665
rect 14461 12631 14519 12637
rect 14461 12628 14473 12631
rect 14056 12600 14473 12628
rect 14056 12588 14062 12600
rect 14461 12597 14473 12600
rect 14507 12597 14519 12631
rect 14461 12591 14519 12597
rect 14553 12631 14611 12637
rect 14553 12597 14565 12631
rect 14599 12628 14611 12631
rect 14921 12631 14979 12637
rect 14921 12628 14933 12631
rect 14599 12600 14933 12628
rect 14599 12597 14611 12600
rect 14553 12591 14611 12597
rect 14921 12597 14933 12600
rect 14967 12597 14979 12631
rect 14921 12591 14979 12597
rect 16761 12631 16819 12637
rect 16761 12597 16773 12631
rect 16807 12628 16819 12631
rect 17313 12631 17371 12637
rect 17313 12628 17325 12631
rect 16807 12600 17325 12628
rect 16807 12597 16819 12600
rect 16761 12591 16819 12597
rect 17313 12597 17325 12600
rect 17359 12597 17371 12631
rect 17313 12591 17371 12597
rect 19242 12588 19248 12640
rect 19300 12628 19306 12640
rect 19705 12631 19763 12637
rect 19705 12628 19717 12631
rect 19300 12600 19717 12628
rect 19300 12588 19306 12600
rect 19705 12597 19717 12600
rect 19751 12597 19763 12631
rect 19705 12591 19763 12597
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 2590 12424 2596 12436
rect 2551 12396 2596 12424
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 2685 12427 2743 12433
rect 2685 12393 2697 12427
rect 2731 12424 2743 12427
rect 3605 12427 3663 12433
rect 3605 12424 3617 12427
rect 2731 12396 3617 12424
rect 2731 12393 2743 12396
rect 2685 12387 2743 12393
rect 3605 12393 3617 12396
rect 3651 12393 3663 12427
rect 3970 12424 3976 12436
rect 3931 12396 3976 12424
rect 3605 12387 3663 12393
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4341 12427 4399 12433
rect 4341 12393 4353 12427
rect 4387 12424 4399 12427
rect 5718 12424 5724 12436
rect 4387 12396 5724 12424
rect 4387 12393 4399 12396
rect 4341 12387 4399 12393
rect 1673 12359 1731 12365
rect 1673 12325 1685 12359
rect 1719 12356 1731 12359
rect 1719 12328 4016 12356
rect 1719 12325 1731 12328
rect 1673 12319 1731 12325
rect 1394 12248 1400 12300
rect 1452 12288 1458 12300
rect 1489 12291 1547 12297
rect 1489 12288 1501 12291
rect 1452 12260 1501 12288
rect 1452 12248 1458 12260
rect 1489 12257 1501 12260
rect 1535 12257 1547 12291
rect 2222 12288 2228 12300
rect 2183 12260 2228 12288
rect 1489 12251 1547 12257
rect 1504 12152 1532 12251
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 3145 12291 3203 12297
rect 3145 12257 3157 12291
rect 3191 12288 3203 12291
rect 3602 12288 3608 12300
rect 3191 12260 3608 12288
rect 3191 12257 3203 12260
rect 3145 12251 3203 12257
rect 3602 12248 3608 12260
rect 3660 12248 3666 12300
rect 3988 12288 4016 12328
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 4890 12356 4896 12368
rect 4120 12328 4896 12356
rect 4120 12316 4126 12328
rect 4154 12288 4160 12300
rect 3988 12260 4160 12288
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 4663 12288 4691 12328
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 5074 12316 5080 12368
rect 5132 12356 5138 12368
rect 5350 12356 5356 12368
rect 5132 12328 5356 12356
rect 5132 12316 5138 12328
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 5460 12300 5488 12396
rect 5718 12384 5724 12396
rect 5776 12384 5782 12436
rect 7653 12427 7711 12433
rect 7653 12393 7665 12427
rect 7699 12424 7711 12427
rect 8205 12427 8263 12433
rect 8205 12424 8217 12427
rect 7699 12396 8217 12424
rect 7699 12393 7711 12396
rect 7653 12387 7711 12393
rect 8205 12393 8217 12396
rect 8251 12393 8263 12427
rect 8205 12387 8263 12393
rect 8665 12427 8723 12433
rect 8665 12393 8677 12427
rect 8711 12424 8723 12427
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 8711 12396 9137 12424
rect 8711 12393 8723 12396
rect 8665 12387 8723 12393
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 9125 12387 9183 12393
rect 9214 12384 9220 12436
rect 9272 12424 9278 12436
rect 9582 12424 9588 12436
rect 9272 12396 9588 12424
rect 9272 12384 9278 12396
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 10042 12424 10048 12436
rect 10003 12396 10048 12424
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10321 12427 10379 12433
rect 10321 12424 10333 12427
rect 10192 12396 10333 12424
rect 10192 12384 10198 12396
rect 10321 12393 10333 12396
rect 10367 12424 10379 12427
rect 10870 12424 10876 12436
rect 10367 12396 10876 12424
rect 10367 12393 10379 12396
rect 10321 12387 10379 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 12066 12424 12072 12436
rect 11848 12396 12072 12424
rect 11848 12384 11854 12396
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 12618 12424 12624 12436
rect 12579 12396 12624 12424
rect 12618 12384 12624 12396
rect 12676 12424 12682 12436
rect 12894 12424 12900 12436
rect 12676 12396 12900 12424
rect 12676 12384 12682 12396
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 13354 12384 13360 12436
rect 13412 12384 13418 12436
rect 13446 12384 13452 12436
rect 13504 12424 13510 12436
rect 15194 12424 15200 12436
rect 13504 12396 15200 12424
rect 13504 12384 13510 12396
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 16209 12427 16267 12433
rect 16209 12393 16221 12427
rect 16255 12424 16267 12427
rect 16390 12424 16396 12436
rect 16255 12396 16396 12424
rect 16255 12393 16267 12396
rect 16209 12387 16267 12393
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 16577 12427 16635 12433
rect 16577 12393 16589 12427
rect 16623 12424 16635 12427
rect 16850 12424 16856 12436
rect 16623 12396 16856 12424
rect 16623 12393 16635 12396
rect 16577 12387 16635 12393
rect 16850 12384 16856 12396
rect 16908 12384 16914 12436
rect 17586 12384 17592 12436
rect 17644 12424 17650 12436
rect 19242 12424 19248 12436
rect 17644 12396 19248 12424
rect 17644 12384 17650 12396
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 19978 12384 19984 12436
rect 20036 12384 20042 12436
rect 20162 12424 20168 12436
rect 20123 12396 20168 12424
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 6454 12316 6460 12368
rect 6512 12356 6518 12368
rect 6672 12359 6730 12365
rect 6672 12356 6684 12359
rect 6512 12328 6684 12356
rect 6512 12316 6518 12328
rect 6672 12325 6684 12328
rect 6718 12356 6730 12359
rect 6718 12328 7880 12356
rect 6718 12325 6730 12328
rect 6672 12319 6730 12325
rect 4632 12260 4691 12288
rect 4801 12291 4859 12297
rect 1946 12220 1952 12232
rect 1907 12192 1952 12220
rect 1946 12180 1952 12192
rect 2004 12180 2010 12232
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 3234 12220 3240 12232
rect 2179 12192 2820 12220
rect 3195 12192 3240 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2792 12161 2820 12192
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 4632 12229 4660 12260
rect 4801 12257 4813 12291
rect 4847 12288 4859 12291
rect 5258 12288 5264 12300
rect 4847 12260 5264 12288
rect 4847 12257 4859 12260
rect 4801 12251 4859 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 5442 12248 5448 12300
rect 5500 12248 5506 12300
rect 6822 12248 6828 12300
rect 6880 12288 6886 12300
rect 6917 12291 6975 12297
rect 6917 12288 6929 12291
rect 6880 12260 6929 12288
rect 6880 12248 6886 12260
rect 6917 12257 6929 12260
rect 6963 12257 6975 12291
rect 6917 12251 6975 12257
rect 7101 12291 7159 12297
rect 7101 12257 7113 12291
rect 7147 12288 7159 12291
rect 7374 12288 7380 12300
rect 7147 12260 7380 12288
rect 7147 12257 7159 12260
rect 7101 12251 7159 12257
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7558 12288 7564 12300
rect 7519 12260 7564 12288
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 7852 12229 7880 12328
rect 8018 12316 8024 12368
rect 8076 12356 8082 12368
rect 8573 12359 8631 12365
rect 8573 12356 8585 12359
rect 8076 12328 8585 12356
rect 8076 12316 8082 12328
rect 8573 12325 8585 12328
rect 8619 12325 8631 12359
rect 8573 12319 8631 12325
rect 9493 12359 9551 12365
rect 9493 12325 9505 12359
rect 9539 12356 9551 12359
rect 10502 12356 10508 12368
rect 9539 12328 10508 12356
rect 9539 12325 9551 12328
rect 9493 12319 9551 12325
rect 10502 12316 10508 12328
rect 10560 12316 10566 12368
rect 11330 12316 11336 12368
rect 11388 12356 11394 12368
rect 11434 12359 11492 12365
rect 11434 12356 11446 12359
rect 11388 12328 11446 12356
rect 11388 12316 11394 12328
rect 11434 12325 11446 12328
rect 11480 12325 11492 12359
rect 11434 12319 11492 12325
rect 11716 12328 12664 12356
rect 11716 12300 11744 12328
rect 8294 12248 8300 12300
rect 8352 12288 8358 12300
rect 8352 12260 8892 12288
rect 8352 12248 8358 12260
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 7837 12223 7895 12229
rect 4755 12192 5396 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 2685 12155 2743 12161
rect 2685 12152 2697 12155
rect 1504 12124 2697 12152
rect 2685 12121 2697 12124
rect 2731 12121 2743 12155
rect 2685 12115 2743 12121
rect 2777 12155 2835 12161
rect 2777 12121 2789 12155
rect 2823 12121 2835 12155
rect 2777 12115 2835 12121
rect 2590 12044 2596 12096
rect 2648 12084 2654 12096
rect 3344 12084 3372 12183
rect 5368 12164 5396 12192
rect 7837 12189 7849 12223
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 8018 12180 8024 12232
rect 8076 12220 8082 12232
rect 8202 12220 8208 12232
rect 8076 12192 8208 12220
rect 8076 12180 8082 12192
rect 8202 12180 8208 12192
rect 8260 12220 8266 12232
rect 8757 12223 8815 12229
rect 8757 12220 8769 12223
rect 8260 12192 8769 12220
rect 8260 12180 8266 12192
rect 8757 12189 8769 12192
rect 8803 12189 8815 12223
rect 8864 12220 8892 12260
rect 9030 12248 9036 12300
rect 9088 12288 9094 12300
rect 10870 12288 10876 12300
rect 9088 12260 10876 12288
rect 9088 12248 9094 12260
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 12158 12288 12164 12300
rect 11756 12260 11801 12288
rect 12119 12260 12164 12288
rect 11756 12248 11762 12260
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12636 12288 12664 12328
rect 12710 12316 12716 12368
rect 12768 12356 12774 12368
rect 13078 12365 13084 12368
rect 13050 12359 13084 12365
rect 13050 12356 13062 12359
rect 12768 12328 13062 12356
rect 12768 12316 12774 12328
rect 13050 12325 13062 12328
rect 13136 12356 13142 12368
rect 13136 12328 13198 12356
rect 13050 12319 13084 12325
rect 13078 12316 13084 12319
rect 13136 12316 13142 12328
rect 13262 12316 13268 12368
rect 13320 12356 13326 12368
rect 13372 12356 13400 12384
rect 13320 12328 13400 12356
rect 13320 12316 13326 12328
rect 13630 12316 13636 12368
rect 13688 12356 13694 12368
rect 13998 12356 14004 12368
rect 13688 12328 14004 12356
rect 13688 12316 13694 12328
rect 13998 12316 14004 12328
rect 14056 12356 14062 12368
rect 14369 12359 14427 12365
rect 14369 12356 14381 12359
rect 14056 12328 14381 12356
rect 14056 12316 14062 12328
rect 14369 12325 14381 12328
rect 14415 12356 14427 12359
rect 14550 12356 14556 12368
rect 14415 12328 14556 12356
rect 14415 12325 14427 12328
rect 14369 12319 14427 12325
rect 14550 12316 14556 12328
rect 14608 12316 14614 12368
rect 14734 12316 14740 12368
rect 14792 12356 14798 12368
rect 14982 12359 15040 12365
rect 14982 12356 14994 12359
rect 14792 12328 14994 12356
rect 14792 12316 14798 12328
rect 14982 12325 14994 12328
rect 15028 12325 15040 12359
rect 14982 12319 15040 12325
rect 16482 12316 16488 12368
rect 16540 12356 16546 12368
rect 16758 12356 16764 12368
rect 16540 12328 16764 12356
rect 16540 12316 16546 12328
rect 16758 12316 16764 12328
rect 16816 12316 16822 12368
rect 17052 12328 18184 12356
rect 17052 12297 17080 12328
rect 12805 12291 12863 12297
rect 12805 12288 12817 12291
rect 12636 12260 12817 12288
rect 12805 12257 12817 12260
rect 12851 12257 12863 12291
rect 17037 12291 17095 12297
rect 17037 12288 17049 12291
rect 12805 12251 12863 12257
rect 16684 12260 17049 12288
rect 9677 12223 9735 12229
rect 9677 12220 9689 12223
rect 8864 12192 9689 12220
rect 8757 12183 8815 12189
rect 9677 12189 9689 12192
rect 9723 12189 9735 12223
rect 9677 12183 9735 12189
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 10042 12220 10048 12232
rect 9824 12192 10048 12220
rect 9824 12180 9830 12192
rect 10042 12180 10048 12192
rect 10100 12220 10106 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10100 12192 10149 12220
rect 10100 12180 10106 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 5350 12152 5356 12164
rect 5311 12124 5356 12152
rect 5350 12112 5356 12124
rect 5408 12112 5414 12164
rect 7098 12112 7104 12164
rect 7156 12152 7162 12164
rect 9858 12152 9864 12164
rect 7156 12124 7788 12152
rect 7156 12112 7162 12124
rect 7760 12096 7788 12124
rect 8772 12124 9864 12152
rect 8772 12096 8800 12124
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 2648 12056 3372 12084
rect 2648 12044 2654 12056
rect 4890 12044 4896 12096
rect 4948 12084 4954 12096
rect 5169 12087 5227 12093
rect 5169 12084 5181 12087
rect 4948 12056 5181 12084
rect 4948 12044 4954 12056
rect 5169 12053 5181 12056
rect 5215 12053 5227 12087
rect 5534 12084 5540 12096
rect 5495 12056 5540 12084
rect 5169 12047 5227 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 7190 12084 7196 12096
rect 7151 12056 7196 12084
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 8021 12087 8079 12093
rect 8021 12084 8033 12087
rect 7800 12056 8033 12084
rect 7800 12044 7806 12056
rect 8021 12053 8033 12056
rect 8067 12053 8079 12087
rect 8021 12047 8079 12053
rect 8754 12044 8760 12096
rect 8812 12044 8818 12096
rect 10152 12084 10180 12183
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10410 12220 10416 12232
rect 10284 12192 10416 12220
rect 10284 12180 10290 12192
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 11974 12220 11980 12232
rect 11935 12192 11980 12220
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 14734 12220 14740 12232
rect 12124 12192 12169 12220
rect 14695 12192 14740 12220
rect 12124 12180 12130 12192
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 16574 12180 16580 12232
rect 16632 12220 16638 12232
rect 16684 12229 16712 12260
rect 17037 12257 17049 12260
rect 17083 12257 17095 12291
rect 17494 12288 17500 12300
rect 17455 12260 17500 12288
rect 17037 12251 17095 12257
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 17764 12291 17822 12297
rect 17764 12257 17776 12291
rect 17810 12288 17822 12291
rect 18046 12288 18052 12300
rect 17810 12260 18052 12288
rect 17810 12257 17822 12260
rect 17764 12251 17822 12257
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 18156 12288 18184 12328
rect 18782 12316 18788 12368
rect 18840 12356 18846 12368
rect 19996 12356 20024 12384
rect 21174 12356 21180 12368
rect 18840 12328 20024 12356
rect 21135 12328 21180 12356
rect 18840 12316 18846 12328
rect 21174 12316 21180 12328
rect 21232 12316 21238 12368
rect 19702 12288 19708 12300
rect 18156 12260 19708 12288
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 19978 12288 19984 12300
rect 19939 12260 19984 12288
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 20990 12288 20996 12300
rect 20951 12260 20996 12288
rect 20990 12248 20996 12260
rect 21048 12248 21054 12300
rect 21361 12291 21419 12297
rect 21361 12257 21373 12291
rect 21407 12288 21419 12291
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 21407 12260 22017 12288
rect 21407 12257 21419 12260
rect 21361 12251 21419 12257
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 16669 12223 16727 12229
rect 16669 12220 16681 12223
rect 16632 12192 16681 12220
rect 16632 12180 16638 12192
rect 16669 12189 16681 12192
rect 16715 12189 16727 12223
rect 16669 12183 16727 12189
rect 16758 12180 16764 12232
rect 16816 12220 16822 12232
rect 16816 12192 16861 12220
rect 16816 12180 16822 12192
rect 18598 12180 18604 12232
rect 18656 12220 18662 12232
rect 20806 12220 20812 12232
rect 18656 12192 20812 12220
rect 18656 12180 18662 12192
rect 20806 12180 20812 12192
rect 20864 12180 20870 12232
rect 16022 12112 16028 12164
rect 16080 12152 16086 12164
rect 16942 12152 16948 12164
rect 16080 12124 16948 12152
rect 16080 12112 16086 12124
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 18506 12112 18512 12164
rect 18564 12152 18570 12164
rect 20254 12152 20260 12164
rect 18564 12124 20260 12152
rect 18564 12112 18570 12124
rect 20254 12112 20260 12124
rect 20312 12112 20318 12164
rect 21542 12152 21548 12164
rect 21503 12124 21548 12152
rect 21542 12112 21548 12124
rect 21600 12112 21606 12164
rect 11974 12084 11980 12096
rect 10152 12056 11980 12084
rect 11974 12044 11980 12056
rect 12032 12084 12038 12096
rect 12342 12084 12348 12096
rect 12032 12056 12348 12084
rect 12032 12044 12038 12056
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12526 12084 12532 12096
rect 12487 12056 12532 12084
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 14185 12087 14243 12093
rect 14185 12053 14197 12087
rect 14231 12084 14243 12087
rect 14274 12084 14280 12096
rect 14231 12056 14280 12084
rect 14231 12053 14243 12056
rect 14185 12047 14243 12053
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 15838 12044 15844 12096
rect 15896 12084 15902 12096
rect 16117 12087 16175 12093
rect 16117 12084 16129 12087
rect 15896 12056 16129 12084
rect 15896 12044 15902 12056
rect 16117 12053 16129 12056
rect 16163 12053 16175 12087
rect 16117 12047 16175 12053
rect 17126 12044 17132 12096
rect 17184 12084 17190 12096
rect 17313 12087 17371 12093
rect 17313 12084 17325 12087
rect 17184 12056 17325 12084
rect 17184 12044 17190 12056
rect 17313 12053 17325 12056
rect 17359 12053 17371 12087
rect 17313 12047 17371 12053
rect 17678 12044 17684 12096
rect 17736 12084 17742 12096
rect 18598 12084 18604 12096
rect 17736 12056 18604 12084
rect 17736 12044 17742 12056
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 18690 12044 18696 12096
rect 18748 12084 18754 12096
rect 18874 12084 18880 12096
rect 18748 12056 18880 12084
rect 18748 12044 18754 12056
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 19061 12087 19119 12093
rect 19061 12053 19073 12087
rect 19107 12084 19119 12087
rect 19150 12084 19156 12096
rect 19107 12056 19156 12084
rect 19107 12053 19119 12056
rect 19061 12047 19119 12053
rect 19150 12044 19156 12056
rect 19208 12044 19214 12096
rect 20162 12044 20168 12096
rect 20220 12084 20226 12096
rect 20622 12084 20628 12096
rect 20220 12056 20628 12084
rect 20220 12044 20226 12056
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 20809 12087 20867 12093
rect 20809 12053 20821 12087
rect 20855 12084 20867 12087
rect 21450 12084 21456 12096
rect 20855 12056 21456 12084
rect 20855 12053 20867 12056
rect 20809 12047 20867 12053
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 1489 11883 1547 11889
rect 1489 11849 1501 11883
rect 1535 11880 1547 11883
rect 1946 11880 1952 11892
rect 1535 11852 1952 11880
rect 1535 11849 1547 11852
rect 1489 11843 1547 11849
rect 1946 11840 1952 11852
rect 2004 11840 2010 11892
rect 2958 11880 2964 11892
rect 2919 11852 2964 11880
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 3050 11840 3056 11892
rect 3108 11880 3114 11892
rect 3237 11883 3295 11889
rect 3237 11880 3249 11883
rect 3108 11852 3249 11880
rect 3108 11840 3114 11852
rect 3237 11849 3249 11852
rect 3283 11849 3295 11883
rect 3602 11880 3608 11892
rect 3563 11852 3608 11880
rect 3237 11843 3295 11849
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4433 11883 4491 11889
rect 4433 11880 4445 11883
rect 4304 11852 4445 11880
rect 4304 11840 4310 11852
rect 4433 11849 4445 11852
rect 4479 11849 4491 11883
rect 4433 11843 4491 11849
rect 5537 11883 5595 11889
rect 5537 11849 5549 11883
rect 5583 11880 5595 11883
rect 5626 11880 5632 11892
rect 5583 11852 5632 11880
rect 5583 11849 5595 11852
rect 5537 11843 5595 11849
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 6454 11880 6460 11892
rect 6415 11852 6460 11880
rect 6454 11840 6460 11852
rect 6512 11840 6518 11892
rect 7926 11840 7932 11892
rect 7984 11880 7990 11892
rect 8757 11883 8815 11889
rect 8757 11880 8769 11883
rect 7984 11852 8769 11880
rect 7984 11840 7990 11852
rect 8757 11849 8769 11852
rect 8803 11849 8815 11883
rect 8757 11843 8815 11849
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 10594 11880 10600 11892
rect 9272 11852 10600 11880
rect 9272 11840 9278 11852
rect 10594 11840 10600 11852
rect 10652 11840 10658 11892
rect 10689 11883 10747 11889
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 12066 11880 12072 11892
rect 10735 11852 12072 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 13265 11883 13323 11889
rect 13265 11849 13277 11883
rect 13311 11880 13323 11883
rect 14458 11880 14464 11892
rect 13311 11852 14464 11880
rect 13311 11849 13323 11852
rect 13265 11843 13323 11849
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 14734 11840 14740 11892
rect 14792 11880 14798 11892
rect 14792 11852 15148 11880
rect 14792 11840 14798 11852
rect 7834 11772 7840 11824
rect 7892 11812 7898 11824
rect 7892 11784 8800 11812
rect 7892 11772 7898 11784
rect 2866 11744 2872 11756
rect 2827 11716 2872 11744
rect 2866 11704 2872 11716
rect 2924 11704 2930 11756
rect 3694 11704 3700 11756
rect 3752 11744 3758 11756
rect 4157 11747 4215 11753
rect 4157 11744 4169 11747
rect 3752 11716 4169 11744
rect 3752 11704 3758 11716
rect 4157 11713 4169 11716
rect 4203 11713 4215 11747
rect 4982 11744 4988 11756
rect 4943 11716 4988 11744
rect 4157 11707 4215 11713
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 6089 11747 6147 11753
rect 6089 11744 6101 11747
rect 5592 11716 6101 11744
rect 5592 11704 5598 11716
rect 6089 11713 6101 11716
rect 6135 11744 6147 11747
rect 6546 11744 6552 11756
rect 6135 11716 6552 11744
rect 6135 11713 6147 11716
rect 6089 11707 6147 11713
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11744 8171 11747
rect 8294 11744 8300 11756
rect 8159 11716 8300 11744
rect 8159 11713 8171 11716
rect 8113 11707 8171 11713
rect 8294 11704 8300 11716
rect 8352 11744 8358 11756
rect 8772 11744 8800 11784
rect 8846 11772 8852 11824
rect 8904 11812 8910 11824
rect 11701 11815 11759 11821
rect 11701 11812 11713 11815
rect 8904 11784 9904 11812
rect 8904 11772 8910 11784
rect 9030 11744 9036 11756
rect 8352 11716 8708 11744
rect 8772 11716 9036 11744
rect 8352 11704 8358 11716
rect 2590 11636 2596 11688
rect 2648 11685 2654 11688
rect 2648 11676 2660 11685
rect 3145 11679 3203 11685
rect 2648 11648 2693 11676
rect 2648 11639 2660 11648
rect 3145 11645 3157 11679
rect 3191 11645 3203 11679
rect 3145 11639 3203 11645
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11645 3479 11679
rect 4890 11676 4896 11688
rect 4851 11648 4896 11676
rect 3421 11639 3479 11645
rect 2648 11636 2654 11639
rect 2038 11568 2044 11620
rect 2096 11608 2102 11620
rect 3160 11608 3188 11639
rect 2096 11580 3188 11608
rect 2096 11568 2102 11580
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3436 11540 3464 11639
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5997 11679 6055 11685
rect 5997 11645 6009 11679
rect 6043 11676 6055 11679
rect 7190 11676 7196 11688
rect 6043 11648 7196 11676
rect 6043 11645 6055 11648
rect 5997 11639 6055 11645
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11676 7895 11679
rect 8570 11676 8576 11688
rect 7883 11648 8576 11676
rect 7883 11645 7895 11648
rect 7837 11639 7895 11645
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 8680 11676 8708 11716
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 9140 11716 9321 11744
rect 9140 11676 9168 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 9766 11744 9772 11756
rect 9309 11707 9367 11713
rect 9646 11716 9772 11744
rect 8680 11648 9168 11676
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11676 9275 11679
rect 9646 11676 9674 11716
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 9876 11685 9904 11784
rect 10244 11784 11713 11812
rect 10134 11744 10140 11756
rect 10095 11716 10140 11744
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 10244 11753 10272 11784
rect 11701 11781 11713 11784
rect 11747 11781 11759 11815
rect 11701 11775 11759 11781
rect 12526 11772 12532 11824
rect 12584 11812 12590 11824
rect 15120 11812 15148 11852
rect 15562 11840 15568 11892
rect 15620 11880 15626 11892
rect 15620 11852 18000 11880
rect 15620 11840 15626 11852
rect 12584 11784 12848 11812
rect 12584 11772 12590 11784
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 11146 11744 11152 11756
rect 10229 11707 10287 11713
rect 10428 11716 11152 11744
rect 9263 11648 9674 11676
rect 9861 11679 9919 11685
rect 9263 11645 9275 11648
rect 9217 11639 9275 11645
rect 9861 11645 9873 11679
rect 9907 11676 9919 11679
rect 10428 11676 10456 11716
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11333 11747 11391 11753
rect 11333 11744 11345 11747
rect 11296 11716 11345 11744
rect 11296 11704 11302 11716
rect 11333 11713 11345 11716
rect 11379 11744 11391 11747
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 11379 11716 12265 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 12253 11713 12265 11716
rect 12299 11713 12311 11747
rect 12710 11744 12716 11756
rect 12671 11716 12716 11744
rect 12253 11707 12311 11713
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 12820 11753 12848 11784
rect 15120 11784 16988 11812
rect 15120 11753 15148 11784
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 15105 11747 15163 11753
rect 15105 11713 15117 11747
rect 15151 11713 15163 11747
rect 15105 11707 15163 11713
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11744 16267 11747
rect 16255 11716 16896 11744
rect 16255 11713 16267 11716
rect 16209 11707 16267 11713
rect 9907 11648 10456 11676
rect 9907 11645 9919 11648
rect 9861 11639 9919 11645
rect 10502 11636 10508 11688
rect 10560 11676 10566 11688
rect 12161 11679 12219 11685
rect 12161 11676 12173 11679
rect 10560 11648 12173 11676
rect 10560 11636 10566 11648
rect 12161 11645 12173 11648
rect 12207 11645 12219 11679
rect 12161 11639 12219 11645
rect 3973 11611 4031 11617
rect 3973 11577 3985 11611
rect 4019 11608 4031 11611
rect 4019 11580 4292 11608
rect 4019 11577 4031 11580
rect 3973 11571 4031 11577
rect 3016 11512 3464 11540
rect 3016 11500 3022 11512
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 3878 11540 3884 11552
rect 3660 11512 3884 11540
rect 3660 11500 3666 11512
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 4154 11540 4160 11552
rect 4111 11512 4160 11540
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4264 11540 4292 11580
rect 4338 11568 4344 11620
rect 4396 11608 4402 11620
rect 4801 11611 4859 11617
rect 4801 11608 4813 11611
rect 4396 11580 4813 11608
rect 4396 11568 4402 11580
rect 4801 11577 4813 11580
rect 4847 11577 4859 11611
rect 5626 11608 5632 11620
rect 4801 11571 4859 11577
rect 5184 11580 5632 11608
rect 5184 11540 5212 11580
rect 5626 11568 5632 11580
rect 5684 11568 5690 11620
rect 7466 11568 7472 11620
rect 7524 11608 7530 11620
rect 7570 11611 7628 11617
rect 7570 11608 7582 11611
rect 7524 11580 7582 11608
rect 7524 11568 7530 11580
rect 7570 11577 7582 11580
rect 7616 11608 7628 11611
rect 8018 11608 8024 11620
rect 7616 11580 8024 11608
rect 7616 11577 7628 11580
rect 7570 11571 7628 11577
rect 8018 11568 8024 11580
rect 8076 11568 8082 11620
rect 8205 11611 8263 11617
rect 8205 11577 8217 11611
rect 8251 11608 8263 11611
rect 10321 11611 10379 11617
rect 8251 11580 8800 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 8772 11552 8800 11580
rect 10321 11577 10333 11611
rect 10367 11608 10379 11611
rect 10367 11580 10824 11608
rect 10367 11577 10379 11580
rect 10321 11571 10379 11577
rect 4264 11512 5212 11540
rect 5261 11543 5319 11549
rect 5261 11509 5273 11543
rect 5307 11540 5319 11543
rect 5534 11540 5540 11552
rect 5307 11512 5540 11540
rect 5307 11509 5319 11512
rect 5261 11503 5319 11509
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5902 11540 5908 11552
rect 5863 11512 5908 11540
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 6822 11540 6828 11552
rect 6696 11512 6828 11540
rect 6696 11500 6702 11512
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 8294 11540 8300 11552
rect 8255 11512 8300 11540
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 8570 11500 8576 11552
rect 8628 11540 8634 11552
rect 8665 11543 8723 11549
rect 8665 11540 8677 11543
rect 8628 11512 8677 11540
rect 8628 11500 8634 11512
rect 8665 11509 8677 11512
rect 8711 11509 8723 11543
rect 8665 11503 8723 11509
rect 8754 11500 8760 11552
rect 8812 11500 8818 11552
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 8904 11512 9137 11540
rect 8904 11500 8910 11512
rect 9125 11509 9137 11512
rect 9171 11509 9183 11543
rect 9125 11503 9183 11509
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 9548 11512 9597 11540
rect 9548 11500 9554 11512
rect 9585 11509 9597 11512
rect 9631 11540 9643 11543
rect 10686 11540 10692 11552
rect 9631 11512 10692 11540
rect 9631 11509 9643 11512
rect 9585 11503 9643 11509
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 10796 11549 10824 11580
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 11241 11611 11299 11617
rect 11241 11608 11253 11611
rect 11112 11580 11253 11608
rect 11112 11568 11118 11580
rect 11241 11577 11253 11580
rect 11287 11577 11299 11611
rect 11241 11571 11299 11577
rect 11974 11568 11980 11620
rect 12032 11608 12038 11620
rect 12069 11611 12127 11617
rect 12069 11608 12081 11611
rect 12032 11580 12081 11608
rect 12032 11568 12038 11580
rect 12069 11577 12081 11580
rect 12115 11577 12127 11611
rect 12176 11608 12204 11639
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 14838 11679 14896 11685
rect 14838 11676 14850 11679
rect 14332 11648 14850 11676
rect 14332 11636 14338 11648
rect 14838 11645 14850 11648
rect 14884 11645 14896 11679
rect 14838 11639 14896 11645
rect 15381 11679 15439 11685
rect 15381 11645 15393 11679
rect 15427 11676 15439 11679
rect 15841 11679 15899 11685
rect 15841 11676 15853 11679
rect 15427 11648 15853 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 15841 11645 15853 11648
rect 15887 11676 15899 11679
rect 16298 11676 16304 11688
rect 15887 11648 16304 11676
rect 15887 11645 15899 11648
rect 15841 11639 15899 11645
rect 16298 11636 16304 11648
rect 16356 11636 16362 11688
rect 15565 11611 15623 11617
rect 15565 11608 15577 11611
rect 12176 11580 15577 11608
rect 12069 11571 12127 11577
rect 15565 11577 15577 11580
rect 15611 11608 15623 11611
rect 16022 11608 16028 11620
rect 15611 11580 16028 11608
rect 15611 11577 15623 11580
rect 15565 11571 15623 11577
rect 16022 11568 16028 11580
rect 16080 11608 16086 11620
rect 16666 11608 16672 11620
rect 16080 11580 16672 11608
rect 16080 11568 16086 11580
rect 16666 11568 16672 11580
rect 16724 11568 16730 11620
rect 16868 11608 16896 11716
rect 16960 11688 16988 11784
rect 17972 11744 18000 11852
rect 18138 11840 18144 11892
rect 18196 11880 18202 11892
rect 18417 11883 18475 11889
rect 18417 11880 18429 11883
rect 18196 11852 18429 11880
rect 18196 11840 18202 11852
rect 18417 11849 18429 11852
rect 18463 11849 18475 11883
rect 19978 11880 19984 11892
rect 18417 11843 18475 11849
rect 18524 11852 19840 11880
rect 19939 11852 19984 11880
rect 18046 11772 18052 11824
rect 18104 11812 18110 11824
rect 18325 11815 18383 11821
rect 18325 11812 18337 11815
rect 18104 11784 18337 11812
rect 18104 11772 18110 11784
rect 18325 11781 18337 11784
rect 18371 11781 18383 11815
rect 18325 11775 18383 11781
rect 18524 11744 18552 11852
rect 17972 11716 18552 11744
rect 18616 11784 19472 11812
rect 16942 11636 16948 11688
rect 17000 11676 17006 11688
rect 17494 11676 17500 11688
rect 17000 11648 17500 11676
rect 17000 11636 17006 11648
rect 17494 11636 17500 11648
rect 17552 11636 17558 11688
rect 18046 11636 18052 11688
rect 18104 11676 18110 11688
rect 18616 11676 18644 11784
rect 18874 11744 18880 11756
rect 18835 11716 18880 11744
rect 18874 11704 18880 11716
rect 18932 11704 18938 11756
rect 19058 11744 19064 11756
rect 19019 11716 19064 11744
rect 19058 11704 19064 11716
rect 19116 11704 19122 11756
rect 19444 11753 19472 11784
rect 19518 11772 19524 11824
rect 19576 11772 19582 11824
rect 19812 11812 19840 11852
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 20254 11880 20260 11892
rect 20215 11852 20260 11880
rect 20254 11840 20260 11852
rect 20312 11840 20318 11892
rect 20714 11880 20720 11892
rect 20675 11852 20720 11880
rect 20714 11840 20720 11852
rect 20772 11840 20778 11892
rect 20990 11880 20996 11892
rect 20951 11852 20996 11880
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 21269 11815 21327 11821
rect 21269 11812 21281 11815
rect 19812 11784 21281 11812
rect 21269 11781 21281 11784
rect 21315 11781 21327 11815
rect 21269 11775 21327 11781
rect 19429 11747 19487 11753
rect 19429 11713 19441 11747
rect 19475 11713 19487 11747
rect 19429 11707 19487 11713
rect 18104 11648 18644 11676
rect 18785 11679 18843 11685
rect 18104 11636 18110 11648
rect 18785 11645 18797 11679
rect 18831 11676 18843 11679
rect 19536 11676 19564 11772
rect 21177 11747 21235 11753
rect 21177 11713 21189 11747
rect 21223 11744 21235 11747
rect 21450 11744 21456 11756
rect 21223 11716 21456 11744
rect 21223 11713 21235 11716
rect 21177 11707 21235 11713
rect 21450 11704 21456 11716
rect 21508 11704 21514 11756
rect 18831 11648 19564 11676
rect 19613 11679 19671 11685
rect 18831 11645 18843 11648
rect 18785 11639 18843 11645
rect 19613 11645 19625 11679
rect 19659 11676 19671 11679
rect 19794 11676 19800 11688
rect 19659 11648 19800 11676
rect 19659 11645 19671 11648
rect 19613 11639 19671 11645
rect 19794 11636 19800 11648
rect 19852 11636 19858 11688
rect 20165 11679 20223 11685
rect 20165 11645 20177 11679
rect 20211 11676 20223 11679
rect 20438 11676 20444 11688
rect 20211 11648 20444 11676
rect 20211 11645 20223 11648
rect 20165 11639 20223 11645
rect 20438 11636 20444 11648
rect 20496 11636 20502 11688
rect 20533 11679 20591 11685
rect 20533 11645 20545 11679
rect 20579 11676 20591 11679
rect 20714 11676 20720 11688
rect 20579 11648 20720 11676
rect 20579 11645 20591 11648
rect 20533 11639 20591 11645
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 20809 11679 20867 11685
rect 20809 11645 20821 11679
rect 20855 11645 20867 11679
rect 20809 11639 20867 11645
rect 17212 11611 17270 11617
rect 17212 11608 17224 11611
rect 16868 11580 17224 11608
rect 17212 11577 17224 11580
rect 17258 11608 17270 11611
rect 17402 11608 17408 11620
rect 17258 11580 17408 11608
rect 17258 11577 17270 11580
rect 17212 11571 17270 11577
rect 17402 11568 17408 11580
rect 17460 11568 17466 11620
rect 19521 11611 19579 11617
rect 19521 11608 19533 11611
rect 18708 11580 19533 11608
rect 10781 11543 10839 11549
rect 10781 11509 10793 11543
rect 10827 11509 10839 11543
rect 11146 11540 11152 11552
rect 11107 11512 11152 11540
rect 10781 11503 10839 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12860 11512 12909 11540
rect 12860 11500 12866 11512
rect 12897 11509 12909 11512
rect 12943 11509 12955 11543
rect 13538 11540 13544 11552
rect 13499 11512 13544 11540
rect 12897 11503 12955 11509
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 13630 11500 13636 11552
rect 13688 11540 13694 11552
rect 13725 11543 13783 11549
rect 13725 11540 13737 11543
rect 13688 11512 13737 11540
rect 13688 11500 13694 11512
rect 13725 11509 13737 11512
rect 13771 11509 13783 11543
rect 16298 11540 16304 11552
rect 16259 11512 16304 11540
rect 13725 11503 13783 11509
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 16761 11543 16819 11549
rect 16448 11512 16493 11540
rect 16448 11500 16454 11512
rect 16761 11509 16773 11543
rect 16807 11540 16819 11543
rect 18708 11540 18736 11580
rect 19521 11577 19533 11580
rect 19567 11577 19579 11611
rect 19521 11571 19579 11577
rect 20622 11568 20628 11620
rect 20680 11608 20686 11620
rect 20824 11608 20852 11639
rect 20680 11580 20852 11608
rect 21453 11611 21511 11617
rect 20680 11568 20686 11580
rect 21453 11577 21465 11611
rect 21499 11608 21511 11611
rect 21542 11608 21548 11620
rect 21499 11580 21548 11608
rect 21499 11577 21511 11580
rect 21453 11571 21511 11577
rect 21542 11568 21548 11580
rect 21600 11568 21606 11620
rect 16807 11512 18736 11540
rect 16807 11509 16819 11512
rect 16761 11503 16819 11509
rect 19150 11500 19156 11552
rect 19208 11540 19214 11552
rect 20806 11540 20812 11552
rect 19208 11512 20812 11540
rect 19208 11500 19214 11512
rect 20806 11500 20812 11512
rect 20864 11500 20870 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 1765 11339 1823 11345
rect 1765 11336 1777 11339
rect 1728 11308 1777 11336
rect 1728 11296 1734 11308
rect 1765 11305 1777 11308
rect 1811 11336 1823 11339
rect 2590 11336 2596 11348
rect 1811 11308 2596 11336
rect 1811 11305 1823 11308
rect 1765 11299 1823 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 3234 11296 3240 11348
rect 3292 11336 3298 11348
rect 3881 11339 3939 11345
rect 3881 11336 3893 11339
rect 3292 11308 3893 11336
rect 3292 11296 3298 11308
rect 3881 11305 3893 11308
rect 3927 11305 3939 11339
rect 3881 11299 3939 11305
rect 3970 11296 3976 11348
rect 4028 11336 4034 11348
rect 6089 11339 6147 11345
rect 4028 11308 5672 11336
rect 4028 11296 4034 11308
rect 3605 11271 3663 11277
rect 3605 11268 3617 11271
rect 1504 11240 3617 11268
rect 1504 11212 1532 11240
rect 3605 11237 3617 11240
rect 3651 11237 3663 11271
rect 3605 11231 3663 11237
rect 4062 11228 4068 11280
rect 4120 11268 4126 11280
rect 4120 11240 4752 11268
rect 4120 11228 4126 11240
rect 1486 11200 1492 11212
rect 1447 11172 1492 11200
rect 1486 11160 1492 11172
rect 1544 11160 1550 11212
rect 2866 11160 2872 11212
rect 2924 11209 2930 11212
rect 2924 11200 2936 11209
rect 3326 11200 3332 11212
rect 2924 11172 2969 11200
rect 3287 11172 3332 11200
rect 2924 11163 2936 11172
rect 2924 11160 2930 11163
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 4246 11200 4252 11212
rect 4207 11172 4252 11200
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 4724 11209 4752 11240
rect 4890 11228 4896 11280
rect 4948 11268 4954 11280
rect 5261 11271 5319 11277
rect 5261 11268 5273 11271
rect 4948 11240 5273 11268
rect 4948 11228 4954 11240
rect 5261 11237 5273 11240
rect 5307 11237 5319 11271
rect 5261 11231 5319 11237
rect 5353 11271 5411 11277
rect 5353 11237 5365 11271
rect 5399 11268 5411 11271
rect 5534 11268 5540 11280
rect 5399 11240 5540 11268
rect 5399 11237 5411 11240
rect 5353 11231 5411 11237
rect 5534 11228 5540 11240
rect 5592 11228 5598 11280
rect 5644 11268 5672 11308
rect 6089 11305 6101 11339
rect 6135 11336 6147 11339
rect 7374 11336 7380 11348
rect 6135 11308 7380 11336
rect 6135 11305 6147 11308
rect 6089 11299 6147 11305
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 7558 11296 7564 11348
rect 7616 11336 7622 11348
rect 8113 11339 8171 11345
rect 8113 11336 8125 11339
rect 7616 11308 8125 11336
rect 7616 11296 7622 11308
rect 8113 11305 8125 11308
rect 8159 11305 8171 11339
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 8113 11299 8171 11305
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 9088 11308 9137 11336
rect 9088 11296 9094 11308
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 10594 11336 10600 11348
rect 9125 11299 9183 11305
rect 9876 11308 10456 11336
rect 10555 11308 10600 11336
rect 6181 11271 6239 11277
rect 6181 11268 6193 11271
rect 5644 11240 6193 11268
rect 6181 11237 6193 11240
rect 6227 11237 6239 11271
rect 6181 11231 6239 11237
rect 6546 11228 6552 11280
rect 6604 11268 6610 11280
rect 6886 11271 6944 11277
rect 6886 11268 6898 11271
rect 6604 11240 6898 11268
rect 6604 11228 6610 11240
rect 6886 11237 6898 11240
rect 6932 11237 6944 11271
rect 6886 11231 6944 11237
rect 7098 11228 7104 11280
rect 7156 11268 7162 11280
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 7156 11240 8953 11268
rect 7156 11228 7162 11240
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 9876 11268 9904 11308
rect 8941 11231 8999 11237
rect 9324 11240 9904 11268
rect 4709 11203 4767 11209
rect 4709 11169 4721 11203
rect 4755 11200 4767 11203
rect 4982 11200 4988 11212
rect 4755 11172 4988 11200
rect 4755 11169 4767 11172
rect 4709 11163 4767 11169
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 7466 11200 7472 11212
rect 5920 11172 7472 11200
rect 3145 11135 3203 11141
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 3878 11132 3884 11144
rect 3191 11104 3884 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 3878 11092 3884 11104
rect 3936 11092 3942 11144
rect 4338 11132 4344 11144
rect 4299 11104 4344 11132
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 5920 11141 5948 11172
rect 7466 11160 7472 11172
rect 7524 11200 7530 11212
rect 9324 11209 9352 11240
rect 9950 11228 9956 11280
rect 10008 11268 10014 11280
rect 10045 11271 10103 11277
rect 10045 11268 10057 11271
rect 10008 11240 10057 11268
rect 10008 11228 10014 11240
rect 10045 11237 10057 11240
rect 10091 11237 10103 11271
rect 10045 11231 10103 11237
rect 10137 11271 10195 11277
rect 10137 11237 10149 11271
rect 10183 11268 10195 11271
rect 10428 11268 10456 11308
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 10928 11308 13492 11336
rect 10928 11296 10934 11308
rect 11425 11271 11483 11277
rect 11425 11268 11437 11271
rect 10183 11240 10263 11268
rect 10428 11240 11437 11268
rect 10183 11237 10195 11240
rect 10137 11231 10195 11237
rect 8481 11203 8539 11209
rect 7524 11172 7880 11200
rect 7524 11160 7530 11172
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 5215 11104 5917 11132
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 5905 11101 5917 11104
rect 5951 11101 5963 11135
rect 6638 11132 6644 11144
rect 6599 11104 6644 11132
rect 5905 11095 5963 11101
rect 3694 11024 3700 11076
rect 3752 11064 3758 11076
rect 4448 11064 4476 11095
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 7852 11132 7880 11172
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 9309 11203 9367 11209
rect 8527 11172 9260 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 8665 11135 8723 11141
rect 8665 11132 8677 11135
rect 7852 11104 8677 11132
rect 8665 11101 8677 11104
rect 8711 11101 8723 11135
rect 8665 11095 8723 11101
rect 9232 11076 9260 11172
rect 9309 11169 9321 11203
rect 9355 11169 9367 11203
rect 9309 11163 9367 11169
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11132 9735 11135
rect 9858 11132 9864 11144
rect 9723 11104 9864 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 9858 11092 9864 11104
rect 9916 11092 9922 11144
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11132 10011 11135
rect 10042 11132 10048 11144
rect 9999 11104 10048 11132
rect 9999 11101 10011 11104
rect 9953 11095 10011 11101
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 10134 11092 10140 11144
rect 10192 11132 10198 11144
rect 10235 11132 10263 11240
rect 11425 11237 11437 11240
rect 11471 11268 11483 11271
rect 13170 11268 13176 11280
rect 11471 11240 12848 11268
rect 13131 11240 13176 11268
rect 11471 11237 11483 11240
rect 11425 11231 11483 11237
rect 10502 11160 10508 11212
rect 10560 11200 10566 11212
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 10560 11172 10977 11200
rect 10560 11160 10566 11172
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11057 11203 11115 11209
rect 11057 11169 11069 11203
rect 11103 11200 11115 11203
rect 11974 11200 11980 11212
rect 11103 11172 11980 11200
rect 11103 11169 11115 11172
rect 11057 11163 11115 11169
rect 10192 11104 10263 11132
rect 10192 11092 10198 11104
rect 10686 11092 10692 11144
rect 10744 11132 10750 11144
rect 11072 11132 11100 11163
rect 11974 11160 11980 11172
rect 12032 11200 12038 11212
rect 12434 11200 12440 11212
rect 12032 11172 12440 11200
rect 12032 11160 12038 11172
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 11238 11132 11244 11144
rect 10744 11104 11100 11132
rect 11199 11104 11244 11132
rect 10744 11092 10750 11104
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 11606 11092 11612 11144
rect 11664 11132 11670 11144
rect 11882 11132 11888 11144
rect 11664 11104 11888 11132
rect 11664 11092 11670 11104
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 3752 11036 4476 11064
rect 4893 11067 4951 11073
rect 3752 11024 3758 11036
rect 4893 11033 4905 11067
rect 4939 11064 4951 11067
rect 6086 11064 6092 11076
rect 4939 11036 6092 11064
rect 4939 11033 4951 11036
rect 4893 11027 4951 11033
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 8294 11024 8300 11076
rect 8352 11064 8358 11076
rect 8570 11064 8576 11076
rect 8352 11036 8576 11064
rect 8352 11024 8358 11036
rect 8570 11024 8576 11036
rect 8628 11024 8634 11076
rect 9214 11024 9220 11076
rect 9272 11064 9278 11076
rect 9401 11067 9459 11073
rect 9401 11064 9413 11067
rect 9272 11036 9413 11064
rect 9272 11024 9278 11036
rect 9401 11033 9413 11036
rect 9447 11033 9459 11067
rect 9401 11027 9459 11033
rect 10505 11067 10563 11073
rect 10505 11033 10517 11067
rect 10551 11064 10563 11067
rect 12158 11064 12164 11076
rect 10551 11036 12164 11064
rect 10551 11033 10563 11036
rect 10505 11027 10563 11033
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 12820 11064 12848 11240
rect 13170 11228 13176 11240
rect 13228 11228 13234 11280
rect 13464 11268 13492 11308
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 14737 11339 14795 11345
rect 14737 11336 14749 11339
rect 13596 11308 14749 11336
rect 13596 11296 13602 11308
rect 14737 11305 14749 11308
rect 14783 11305 14795 11339
rect 14737 11299 14795 11305
rect 15105 11339 15163 11345
rect 15105 11305 15117 11339
rect 15151 11336 15163 11339
rect 15565 11339 15623 11345
rect 15565 11336 15577 11339
rect 15151 11308 15577 11336
rect 15151 11305 15163 11308
rect 15105 11299 15163 11305
rect 15565 11305 15577 11308
rect 15611 11305 15623 11339
rect 17589 11339 17647 11345
rect 17589 11336 17601 11339
rect 15565 11299 15623 11305
rect 15663 11308 17601 11336
rect 13722 11268 13728 11280
rect 13464 11240 13728 11268
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 15194 11228 15200 11280
rect 15252 11268 15258 11280
rect 15663 11268 15691 11308
rect 17589 11305 17601 11308
rect 17635 11336 17647 11339
rect 17678 11336 17684 11348
rect 17635 11308 17684 11336
rect 17635 11305 17647 11308
rect 17589 11299 17647 11305
rect 17678 11296 17684 11308
rect 17736 11296 17742 11348
rect 17770 11296 17776 11348
rect 17828 11336 17834 11348
rect 17828 11308 17873 11336
rect 17828 11296 17834 11308
rect 18046 11296 18052 11348
rect 18104 11336 18110 11348
rect 18601 11339 18659 11345
rect 18601 11336 18613 11339
rect 18104 11308 18613 11336
rect 18104 11296 18110 11308
rect 18601 11305 18613 11308
rect 18647 11305 18659 11339
rect 18601 11299 18659 11305
rect 18874 11296 18880 11348
rect 18932 11336 18938 11348
rect 19061 11339 19119 11345
rect 19061 11336 19073 11339
rect 18932 11308 19073 11336
rect 18932 11296 18938 11308
rect 19061 11305 19073 11308
rect 19107 11305 19119 11339
rect 19061 11299 19119 11305
rect 19150 11296 19156 11348
rect 19208 11336 19214 11348
rect 19426 11336 19432 11348
rect 19208 11308 19432 11336
rect 19208 11296 19214 11308
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 19613 11339 19671 11345
rect 19613 11305 19625 11339
rect 19659 11336 19671 11339
rect 19794 11336 19800 11348
rect 19659 11308 19800 11336
rect 19659 11305 19671 11308
rect 19613 11299 19671 11305
rect 19794 11296 19800 11308
rect 19852 11296 19858 11348
rect 20993 11339 21051 11345
rect 20993 11305 21005 11339
rect 21039 11336 21051 11339
rect 22005 11339 22063 11345
rect 22005 11336 22017 11339
rect 21039 11308 22017 11336
rect 21039 11305 21051 11308
rect 20993 11299 21051 11305
rect 22005 11305 22017 11308
rect 22051 11305 22063 11339
rect 22005 11299 22063 11305
rect 16942 11268 16948 11280
rect 15252 11240 15691 11268
rect 16040 11240 16948 11268
rect 15252 11228 15258 11240
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 13633 11203 13691 11209
rect 13633 11200 13645 11203
rect 12952 11172 13645 11200
rect 12952 11160 12958 11172
rect 13633 11169 13645 11172
rect 13679 11169 13691 11203
rect 13633 11163 13691 11169
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11200 14703 11203
rect 14691 11172 14872 11200
rect 14691 11169 14703 11172
rect 14645 11163 14703 11169
rect 14844 11144 14872 11172
rect 14918 11160 14924 11212
rect 14976 11200 14982 11212
rect 16040 11209 16068 11240
rect 16942 11228 16948 11240
rect 17000 11228 17006 11280
rect 21269 11271 21327 11277
rect 21269 11268 21281 11271
rect 17052 11240 21281 11268
rect 16025 11203 16083 11209
rect 14976 11172 15792 11200
rect 14976 11160 14982 11172
rect 13538 11132 13544 11144
rect 13499 11104 13544 11132
rect 13538 11092 13544 11104
rect 13596 11132 13602 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 13596 11104 14473 11132
rect 13596 11092 13602 11104
rect 14461 11101 14473 11104
rect 14507 11132 14519 11135
rect 14550 11132 14556 11144
rect 14507 11104 14556 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 14550 11092 14556 11104
rect 14608 11092 14614 11144
rect 14826 11092 14832 11144
rect 14884 11092 14890 11144
rect 15764 11141 15792 11172
rect 16025 11169 16037 11203
rect 16071 11169 16083 11203
rect 16281 11203 16339 11209
rect 16281 11200 16293 11203
rect 16025 11163 16083 11169
rect 16132 11172 16293 11200
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 15749 11135 15807 11141
rect 15749 11101 15761 11135
rect 15795 11101 15807 11135
rect 16132 11132 16160 11172
rect 16281 11169 16293 11172
rect 16327 11169 16339 11203
rect 16281 11163 16339 11169
rect 15749 11095 15807 11101
rect 16040 11104 16160 11132
rect 13446 11064 13452 11076
rect 12820 11036 13452 11064
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 14093 11067 14151 11073
rect 14093 11033 14105 11067
rect 14139 11064 14151 11067
rect 15672 11064 15700 11095
rect 16040 11076 16068 11104
rect 14139 11036 15700 11064
rect 14139 11033 14151 11036
rect 14093 11027 14151 11033
rect 16022 11024 16028 11076
rect 16080 11024 16086 11076
rect 3421 10999 3479 11005
rect 3421 10965 3433 10999
rect 3467 10996 3479 10999
rect 5258 10996 5264 11008
rect 3467 10968 5264 10996
rect 3467 10965 3479 10968
rect 3421 10959 3479 10965
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 5718 10996 5724 11008
rect 5679 10968 5724 10996
rect 5718 10956 5724 10968
rect 5776 10956 5782 11008
rect 6546 10996 6552 11008
rect 6507 10968 6552 10996
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 8018 10996 8024 11008
rect 7979 10968 8024 10996
rect 8018 10956 8024 10968
rect 8076 10956 8082 11008
rect 8941 10999 8999 11005
rect 8941 10965 8953 10999
rect 8987 10996 8999 10999
rect 13906 10996 13912 11008
rect 8987 10968 13912 10996
rect 8987 10965 8999 10968
rect 8941 10959 8999 10965
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 15194 10996 15200 11008
rect 15155 10968 15200 10996
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 17052 10996 17080 11240
rect 21269 11237 21281 11240
rect 21315 11237 21327 11271
rect 21269 11231 21327 11237
rect 18509 11203 18567 11209
rect 18509 11169 18521 11203
rect 18555 11200 18567 11203
rect 19610 11200 19616 11212
rect 18555 11172 19616 11200
rect 18555 11169 18567 11172
rect 18509 11163 18567 11169
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 19978 11200 19984 11212
rect 19939 11172 19984 11200
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 20438 11160 20444 11212
rect 20496 11200 20502 11212
rect 20809 11203 20867 11209
rect 20809 11200 20821 11203
rect 20496 11172 20821 11200
rect 20496 11160 20502 11172
rect 20809 11169 20821 11172
rect 20855 11169 20867 11203
rect 21450 11200 21456 11212
rect 21411 11172 21456 11200
rect 20809 11163 20867 11169
rect 21450 11160 21456 11172
rect 21508 11160 21514 11212
rect 18046 11132 18052 11144
rect 18007 11104 18052 11132
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18414 11132 18420 11144
rect 18375 11104 18420 11132
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 20073 11135 20131 11141
rect 20073 11132 20085 11135
rect 19392 11104 20085 11132
rect 19392 11092 19398 11104
rect 20073 11101 20085 11104
rect 20119 11101 20131 11135
rect 20073 11095 20131 11101
rect 20165 11135 20223 11141
rect 20165 11101 20177 11135
rect 20211 11101 20223 11135
rect 20165 11095 20223 11101
rect 20717 11135 20775 11141
rect 20717 11101 20729 11135
rect 20763 11132 20775 11135
rect 21082 11132 21088 11144
rect 20763 11104 21088 11132
rect 20763 11101 20775 11104
rect 20717 11095 20775 11101
rect 17402 11064 17408 11076
rect 17315 11036 17408 11064
rect 17402 11024 17408 11036
rect 17460 11064 17466 11076
rect 20180 11064 20208 11095
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 21177 11135 21235 11141
rect 21177 11101 21189 11135
rect 21223 11132 21235 11135
rect 21358 11132 21364 11144
rect 21223 11104 21364 11132
rect 21223 11101 21235 11104
rect 21177 11095 21235 11101
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 17460 11036 20208 11064
rect 17460 11024 17466 11036
rect 20254 11024 20260 11076
rect 20312 11024 20318 11076
rect 15344 10968 17080 10996
rect 18969 10999 19027 11005
rect 15344 10956 15350 10968
rect 18969 10965 18981 10999
rect 19015 10996 19027 10999
rect 19150 10996 19156 11008
rect 19015 10968 19156 10996
rect 19015 10965 19027 10968
rect 18969 10959 19027 10965
rect 19150 10956 19156 10968
rect 19208 10956 19214 11008
rect 19429 10999 19487 11005
rect 19429 10965 19441 10999
rect 19475 10996 19487 10999
rect 19702 10996 19708 11008
rect 19475 10968 19708 10996
rect 19475 10965 19487 10968
rect 19429 10959 19487 10965
rect 19702 10956 19708 10968
rect 19760 10996 19766 11008
rect 20272 10996 20300 11024
rect 19760 10968 20300 10996
rect 20533 10999 20591 11005
rect 19760 10956 19766 10968
rect 20533 10965 20545 10999
rect 20579 10996 20591 10999
rect 20806 10996 20812 11008
rect 20579 10968 20812 10996
rect 20579 10965 20591 10968
rect 20533 10959 20591 10965
rect 20806 10956 20812 10968
rect 20864 10996 20870 11008
rect 22186 10996 22192 11008
rect 20864 10968 22192 10996
rect 20864 10956 20870 10968
rect 22186 10956 22192 10968
rect 22244 10956 22250 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 2222 10792 2228 10804
rect 2183 10764 2228 10792
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 3878 10792 3884 10804
rect 2332 10764 3884 10792
rect 1670 10656 1676 10668
rect 1631 10628 1676 10656
rect 1670 10616 1676 10628
rect 1728 10616 1734 10668
rect 2332 10665 2360 10764
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 4617 10795 4675 10801
rect 4617 10792 4629 10795
rect 4304 10764 4629 10792
rect 4304 10752 4310 10764
rect 4617 10761 4629 10764
rect 4663 10761 4675 10795
rect 5258 10792 5264 10804
rect 4617 10755 4675 10761
rect 4816 10764 5264 10792
rect 4154 10684 4160 10736
rect 4212 10724 4218 10736
rect 4709 10727 4767 10733
rect 4709 10724 4721 10727
rect 4212 10696 4721 10724
rect 4212 10684 4218 10696
rect 4709 10693 4721 10696
rect 4755 10693 4767 10727
rect 4709 10687 4767 10693
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10625 2375 10659
rect 2317 10619 2375 10625
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10656 4031 10659
rect 4816 10656 4844 10764
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5537 10795 5595 10801
rect 5537 10761 5549 10795
rect 5583 10792 5595 10795
rect 5626 10792 5632 10804
rect 5583 10764 5632 10792
rect 5583 10761 5595 10764
rect 5537 10755 5595 10761
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 6457 10795 6515 10801
rect 6457 10792 6469 10795
rect 5960 10764 6469 10792
rect 5960 10752 5966 10764
rect 6457 10761 6469 10764
rect 6503 10761 6515 10795
rect 7374 10792 7380 10804
rect 7335 10764 7380 10792
rect 6457 10755 6515 10761
rect 7374 10752 7380 10764
rect 7432 10752 7438 10804
rect 7484 10764 11008 10792
rect 7098 10724 7104 10736
rect 4019 10628 4844 10656
rect 4908 10696 7104 10724
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 3988 10588 4016 10619
rect 2608 10560 4016 10588
rect 2608 10532 2636 10560
rect 4062 10548 4068 10600
rect 4120 10588 4126 10600
rect 4908 10588 4936 10696
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 5258 10656 5264 10668
rect 5219 10628 5264 10656
rect 5258 10616 5264 10628
rect 5316 10656 5322 10668
rect 6089 10659 6147 10665
rect 6089 10656 6101 10659
rect 5316 10628 6101 10656
rect 5316 10616 5322 10628
rect 6089 10625 6101 10628
rect 6135 10625 6147 10659
rect 6089 10619 6147 10625
rect 6196 10628 6408 10656
rect 4120 10560 4936 10588
rect 5077 10591 5135 10597
rect 4120 10548 4126 10560
rect 5077 10557 5089 10591
rect 5123 10588 5135 10591
rect 5626 10588 5632 10600
rect 5123 10560 5632 10588
rect 5123 10557 5135 10560
rect 5077 10551 5135 10557
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 5718 10548 5724 10600
rect 5776 10588 5782 10600
rect 6196 10588 6224 10628
rect 5776 10560 6224 10588
rect 6380 10588 6408 10628
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 6604 10628 6929 10656
rect 6604 10616 6610 10628
rect 6917 10625 6929 10628
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6380 10560 6837 10588
rect 5776 10548 5782 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 7024 10588 7052 10619
rect 6825 10551 6883 10557
rect 6993 10560 7052 10588
rect 2590 10529 2596 10532
rect 2584 10520 2596 10529
rect 2551 10492 2596 10520
rect 2584 10483 2596 10492
rect 2590 10480 2596 10483
rect 2648 10480 2654 10532
rect 3786 10480 3792 10532
rect 3844 10520 3850 10532
rect 4522 10520 4528 10532
rect 3844 10492 4528 10520
rect 3844 10480 3850 10492
rect 1762 10452 1768 10464
rect 1723 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 1857 10455 1915 10461
rect 1857 10421 1869 10455
rect 1903 10452 1915 10455
rect 2222 10452 2228 10464
rect 1903 10424 2228 10452
rect 1903 10421 1915 10424
rect 1857 10415 1915 10421
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 3694 10452 3700 10464
rect 2924 10424 3700 10452
rect 2924 10412 2930 10424
rect 3694 10412 3700 10424
rect 3752 10412 3758 10464
rect 4172 10461 4200 10492
rect 4522 10480 4528 10492
rect 4580 10480 4586 10532
rect 5169 10523 5227 10529
rect 5169 10489 5181 10523
rect 5215 10520 5227 10523
rect 5534 10520 5540 10532
rect 5215 10492 5540 10520
rect 5215 10489 5227 10492
rect 5169 10483 5227 10489
rect 5534 10480 5540 10492
rect 5592 10480 5598 10532
rect 6454 10480 6460 10532
rect 6512 10520 6518 10532
rect 6993 10520 7021 10560
rect 6512 10492 7021 10520
rect 6512 10480 6518 10492
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10421 4215 10455
rect 4157 10415 4215 10421
rect 4246 10412 4252 10464
rect 4304 10452 4310 10464
rect 4304 10424 4349 10452
rect 4304 10412 4310 10424
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 5905 10455 5963 10461
rect 5905 10452 5917 10455
rect 5408 10424 5917 10452
rect 5408 10412 5414 10424
rect 5905 10421 5917 10424
rect 5951 10421 5963 10455
rect 5905 10415 5963 10421
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 7484 10452 7512 10764
rect 7558 10684 7564 10736
rect 7616 10724 7622 10736
rect 7616 10696 8708 10724
rect 7616 10684 7622 10696
rect 7650 10616 7656 10668
rect 7708 10656 7714 10668
rect 8018 10656 8024 10668
rect 7708 10628 8024 10656
rect 7708 10616 7714 10628
rect 8018 10616 8024 10628
rect 8076 10656 8082 10668
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 8076 10628 8401 10656
rect 8076 10616 8082 10628
rect 8389 10625 8401 10628
rect 8435 10625 8447 10659
rect 8680 10656 8708 10696
rect 8754 10684 8760 10736
rect 8812 10724 8818 10736
rect 9217 10727 9275 10733
rect 9217 10724 9229 10727
rect 8812 10696 9229 10724
rect 8812 10684 8818 10696
rect 9217 10693 9229 10696
rect 9263 10724 9275 10727
rect 9674 10724 9680 10736
rect 9263 10696 9680 10724
rect 9263 10693 9275 10696
rect 9217 10687 9275 10693
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 9125 10659 9183 10665
rect 8680 10628 8984 10656
rect 8389 10619 8447 10625
rect 8297 10591 8355 10597
rect 8297 10557 8309 10591
rect 8343 10588 8355 10591
rect 8757 10591 8815 10597
rect 8757 10588 8769 10591
rect 8343 10560 8769 10588
rect 8343 10557 8355 10560
rect 8297 10551 8355 10557
rect 8757 10557 8769 10560
rect 8803 10588 8815 10591
rect 8846 10588 8852 10600
rect 8803 10560 8852 10588
rect 8803 10557 8815 10560
rect 8757 10551 8815 10557
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 8956 10588 8984 10628
rect 9125 10625 9137 10659
rect 9171 10656 9183 10659
rect 9490 10656 9496 10668
rect 9171 10628 9496 10656
rect 9171 10625 9183 10628
rect 9125 10619 9183 10625
rect 9490 10616 9496 10628
rect 9548 10656 9554 10668
rect 9766 10656 9772 10668
rect 9548 10628 9772 10656
rect 9548 10616 9554 10628
rect 9766 10616 9772 10628
rect 9824 10656 9830 10668
rect 10980 10656 11008 10764
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11333 10795 11391 10801
rect 11333 10792 11345 10795
rect 11296 10764 11345 10792
rect 11296 10752 11302 10764
rect 11333 10761 11345 10764
rect 11379 10761 11391 10795
rect 11333 10755 11391 10761
rect 11517 10795 11575 10801
rect 11517 10761 11529 10795
rect 11563 10792 11575 10795
rect 11974 10792 11980 10804
rect 11563 10764 11980 10792
rect 11563 10761 11575 10764
rect 11517 10755 11575 10761
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 13262 10752 13268 10804
rect 13320 10792 13326 10804
rect 13817 10795 13875 10801
rect 13320 10764 13768 10792
rect 13320 10752 13326 10764
rect 11054 10684 11060 10736
rect 11112 10724 11118 10736
rect 11701 10727 11759 10733
rect 11701 10724 11713 10727
rect 11112 10696 11713 10724
rect 11112 10684 11118 10696
rect 11701 10693 11713 10696
rect 11747 10724 11759 10727
rect 13630 10724 13636 10736
rect 11747 10696 12112 10724
rect 11747 10693 11759 10696
rect 11701 10687 11759 10693
rect 12084 10668 12112 10696
rect 13556 10696 13636 10724
rect 11606 10656 11612 10668
rect 9824 10628 10088 10656
rect 10980 10628 11612 10656
rect 9824 10616 9830 10628
rect 9674 10588 9680 10600
rect 8956 10560 9680 10588
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 9950 10588 9956 10600
rect 9911 10560 9956 10588
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 10060 10588 10088 10628
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12066 10616 12072 10668
rect 12124 10616 12130 10668
rect 13556 10665 13584 10696
rect 13630 10684 13636 10696
rect 13688 10684 13694 10736
rect 13740 10724 13768 10764
rect 13817 10761 13829 10795
rect 13863 10792 13875 10795
rect 14366 10792 14372 10804
rect 13863 10764 14372 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 14734 10752 14740 10804
rect 14792 10792 14798 10804
rect 15013 10795 15071 10801
rect 15013 10792 15025 10795
rect 14792 10764 15025 10792
rect 14792 10752 14798 10764
rect 15013 10761 15025 10764
rect 15059 10761 15071 10795
rect 15013 10755 15071 10761
rect 16025 10795 16083 10801
rect 16025 10761 16037 10795
rect 16071 10792 16083 10795
rect 16298 10792 16304 10804
rect 16071 10764 16304 10792
rect 16071 10761 16083 10764
rect 16025 10755 16083 10761
rect 14918 10724 14924 10736
rect 13740 10696 14924 10724
rect 14918 10684 14924 10696
rect 14976 10684 14982 10736
rect 13541 10659 13599 10665
rect 13541 10625 13553 10659
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 14645 10659 14703 10665
rect 14645 10656 14657 10659
rect 14608 10628 14657 10656
rect 14608 10616 14614 10628
rect 14645 10625 14657 10628
rect 14691 10625 14703 10659
rect 14645 10619 14703 10625
rect 10060 10560 12664 10588
rect 7742 10480 7748 10532
rect 7800 10480 7806 10532
rect 8205 10523 8263 10529
rect 8205 10489 8217 10523
rect 8251 10520 8263 10523
rect 8941 10523 8999 10529
rect 8941 10520 8953 10523
rect 8251 10492 8953 10520
rect 8251 10489 8263 10492
rect 8205 10483 8263 10489
rect 6052 10424 7512 10452
rect 6052 10412 6058 10424
rect 7558 10412 7564 10464
rect 7616 10452 7622 10464
rect 7653 10455 7711 10461
rect 7653 10452 7665 10455
rect 7616 10424 7665 10452
rect 7616 10412 7622 10424
rect 7653 10421 7665 10424
rect 7699 10421 7711 10455
rect 7760 10452 7788 10480
rect 8864 10464 8892 10492
rect 8941 10489 8953 10492
rect 8987 10520 8999 10523
rect 9122 10520 9128 10532
rect 8987 10492 9128 10520
rect 8987 10489 8999 10492
rect 8941 10483 8999 10489
rect 9122 10480 9128 10492
rect 9180 10480 9186 10532
rect 10220 10523 10278 10529
rect 10220 10489 10232 10523
rect 10266 10520 10278 10523
rect 10502 10520 10508 10532
rect 10266 10492 10508 10520
rect 10266 10489 10278 10492
rect 10220 10483 10278 10489
rect 10502 10480 10508 10492
rect 10560 10480 10566 10532
rect 11146 10480 11152 10532
rect 11204 10520 11210 10532
rect 11977 10523 12035 10529
rect 11977 10520 11989 10523
rect 11204 10492 11989 10520
rect 11204 10480 11210 10492
rect 11977 10489 11989 10492
rect 12023 10520 12035 10523
rect 12342 10520 12348 10532
rect 12023 10492 12348 10520
rect 12023 10489 12035 10492
rect 11977 10483 12035 10489
rect 12342 10480 12348 10492
rect 12400 10480 12406 10532
rect 12636 10520 12664 10560
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 13262 10588 13268 10600
rect 13320 10597 13326 10600
rect 12768 10560 13268 10588
rect 12768 10548 12774 10560
rect 13262 10548 13268 10560
rect 13320 10588 13332 10597
rect 13320 10560 13365 10588
rect 13320 10551 13332 10560
rect 13320 10548 13326 10551
rect 13446 10548 13452 10600
rect 13504 10588 13510 10600
rect 13641 10591 13699 10597
rect 13641 10588 13653 10591
rect 13504 10560 13653 10588
rect 13504 10548 13510 10560
rect 13641 10557 13653 10560
rect 13687 10557 13699 10591
rect 13641 10551 13699 10557
rect 13906 10548 13912 10600
rect 13964 10548 13970 10600
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 14734 10588 14740 10600
rect 14148 10560 14740 10588
rect 14148 10548 14154 10560
rect 14734 10548 14740 10560
rect 14792 10548 14798 10600
rect 15028 10588 15056 10755
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 16758 10752 16764 10804
rect 16816 10792 16822 10804
rect 18509 10795 18567 10801
rect 16816 10764 18092 10792
rect 16816 10752 16822 10764
rect 15933 10727 15991 10733
rect 15933 10693 15945 10727
rect 15979 10724 15991 10727
rect 16390 10724 16396 10736
rect 15979 10696 16396 10724
rect 15979 10693 15991 10696
rect 15933 10687 15991 10693
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 18064 10724 18092 10764
rect 18509 10761 18521 10795
rect 18555 10792 18567 10795
rect 19242 10792 19248 10804
rect 18555 10764 19248 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 19337 10795 19395 10801
rect 19337 10761 19349 10795
rect 19383 10792 19395 10795
rect 19978 10792 19984 10804
rect 19383 10764 19984 10792
rect 19383 10761 19395 10764
rect 19337 10755 19395 10761
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 20438 10792 20444 10804
rect 20399 10764 20444 10792
rect 20438 10752 20444 10764
rect 20496 10752 20502 10804
rect 20714 10792 20720 10804
rect 20675 10764 20720 10792
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 20901 10727 20959 10733
rect 20901 10724 20913 10727
rect 16684 10696 18000 10724
rect 18064 10696 20913 10724
rect 15381 10659 15439 10665
rect 15381 10625 15393 10659
rect 15427 10656 15439 10659
rect 16022 10656 16028 10668
rect 15427 10628 16028 10656
rect 15427 10625 15439 10628
rect 15381 10619 15439 10625
rect 16022 10616 16028 10628
rect 16080 10656 16086 10668
rect 16684 10665 16712 10696
rect 17972 10668 18000 10696
rect 20901 10693 20913 10696
rect 20947 10693 20959 10727
rect 20901 10687 20959 10693
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 16080 10628 16681 10656
rect 16080 10616 16086 10628
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 17586 10656 17592 10668
rect 17547 10628 17592 10656
rect 16669 10619 16727 10625
rect 17586 10616 17592 10628
rect 17644 10616 17650 10668
rect 17954 10656 17960 10668
rect 17867 10628 17960 10656
rect 17954 10616 17960 10628
rect 18012 10656 18018 10668
rect 18693 10659 18751 10665
rect 18693 10656 18705 10659
rect 18012 10628 18705 10656
rect 18012 10616 18018 10628
rect 18693 10625 18705 10628
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10656 19671 10659
rect 19886 10656 19892 10668
rect 19659 10628 19892 10656
rect 19659 10625 19671 10628
rect 19613 10619 19671 10625
rect 19886 10616 19892 10628
rect 19944 10616 19950 10668
rect 15565 10591 15623 10597
rect 15565 10588 15577 10591
rect 15028 10560 15577 10588
rect 15565 10557 15577 10560
rect 15611 10557 15623 10591
rect 15565 10551 15623 10557
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10588 16451 10591
rect 16942 10588 16948 10600
rect 16439 10560 16948 10588
rect 16439 10557 16451 10560
rect 16393 10551 16451 10557
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 17310 10588 17316 10600
rect 17271 10560 17316 10588
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 17678 10548 17684 10600
rect 17736 10588 17742 10600
rect 18141 10591 18199 10597
rect 18141 10588 18153 10591
rect 17736 10560 18153 10588
rect 17736 10548 17742 10560
rect 18141 10557 18153 10560
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 18874 10548 18880 10600
rect 18932 10588 18938 10600
rect 18969 10591 19027 10597
rect 18969 10588 18981 10591
rect 18932 10560 18981 10588
rect 18932 10548 18938 10560
rect 18969 10557 18981 10560
rect 19015 10557 19027 10591
rect 18969 10551 19027 10557
rect 19150 10548 19156 10600
rect 19208 10588 19214 10600
rect 20257 10591 20315 10597
rect 20257 10588 20269 10591
rect 19208 10560 20269 10588
rect 19208 10548 19214 10560
rect 20257 10557 20269 10560
rect 20303 10557 20315 10591
rect 20257 10551 20315 10557
rect 20533 10591 20591 10597
rect 20533 10557 20545 10591
rect 20579 10557 20591 10591
rect 20533 10551 20591 10557
rect 13924 10520 13952 10548
rect 12636 10492 13952 10520
rect 14461 10523 14519 10529
rect 14461 10489 14473 10523
rect 14507 10520 14519 10523
rect 15286 10520 15292 10532
rect 14507 10492 15292 10520
rect 14507 10489 14519 10492
rect 14461 10483 14519 10489
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 15473 10523 15531 10529
rect 15473 10489 15485 10523
rect 15519 10520 15531 10523
rect 15519 10492 16988 10520
rect 15519 10489 15531 10492
rect 15473 10483 15531 10489
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7760 10424 7849 10452
rect 7653 10415 7711 10421
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 7837 10415 7895 10421
rect 8846 10412 8852 10464
rect 8904 10412 8910 10464
rect 9306 10412 9312 10464
rect 9364 10452 9370 10464
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9364 10424 9413 10452
rect 9364 10412 9370 10424
rect 9401 10421 9413 10424
rect 9447 10421 9459 10455
rect 9401 10415 9459 10421
rect 9861 10455 9919 10461
rect 9861 10421 9873 10455
rect 9907 10452 9919 10455
rect 10962 10452 10968 10464
rect 9907 10424 10968 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 12161 10455 12219 10461
rect 12161 10421 12173 10455
rect 12207 10452 12219 10455
rect 12802 10452 12808 10464
rect 12207 10424 12808 10452
rect 12207 10421 12219 10424
rect 12161 10415 12219 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 13909 10455 13967 10461
rect 13909 10452 13921 10455
rect 13780 10424 13921 10452
rect 13780 10412 13786 10424
rect 13909 10421 13921 10424
rect 13955 10421 13967 10455
rect 14090 10452 14096 10464
rect 14051 10424 14096 10452
rect 13909 10415 13967 10421
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 14550 10412 14556 10464
rect 14608 10452 14614 10464
rect 14608 10424 14653 10452
rect 14608 10412 14614 10424
rect 16482 10412 16488 10464
rect 16540 10452 16546 10464
rect 16960 10461 16988 10492
rect 17770 10480 17776 10532
rect 17828 10520 17834 10532
rect 18049 10523 18107 10529
rect 18049 10520 18061 10523
rect 17828 10492 18061 10520
rect 17828 10480 17834 10492
rect 18049 10489 18061 10492
rect 18095 10489 18107 10523
rect 20548 10520 20576 10551
rect 21082 10520 21088 10532
rect 18049 10483 18107 10489
rect 20180 10492 20576 10520
rect 21043 10492 21088 10520
rect 16945 10455 17003 10461
rect 16540 10424 16585 10452
rect 16540 10412 16546 10424
rect 16945 10421 16957 10455
rect 16991 10421 17003 10455
rect 16945 10415 17003 10421
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 17405 10455 17463 10461
rect 17405 10452 17417 10455
rect 17276 10424 17417 10452
rect 17276 10412 17282 10424
rect 17405 10421 17417 10424
rect 17451 10421 17463 10455
rect 17405 10415 17463 10421
rect 18877 10455 18935 10461
rect 18877 10421 18889 10455
rect 18923 10452 18935 10455
rect 18966 10452 18972 10464
rect 18923 10424 18972 10452
rect 18923 10421 18935 10424
rect 18877 10415 18935 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 19702 10452 19708 10464
rect 19663 10424 19708 10452
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 19794 10412 19800 10464
rect 19852 10452 19858 10464
rect 20180 10461 20208 10492
rect 21082 10480 21088 10492
rect 21140 10480 21146 10532
rect 21174 10480 21180 10532
rect 21232 10520 21238 10532
rect 21269 10523 21327 10529
rect 21269 10520 21281 10523
rect 21232 10492 21281 10520
rect 21232 10480 21238 10492
rect 21269 10489 21281 10492
rect 21315 10489 21327 10523
rect 21450 10520 21456 10532
rect 21411 10492 21456 10520
rect 21269 10483 21327 10489
rect 21450 10480 21456 10492
rect 21508 10480 21514 10532
rect 20165 10455 20223 10461
rect 19852 10424 19897 10452
rect 19852 10412 19858 10424
rect 20165 10421 20177 10455
rect 20211 10421 20223 10455
rect 20165 10415 20223 10421
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 1857 10251 1915 10257
rect 1857 10217 1869 10251
rect 1903 10248 1915 10251
rect 2317 10251 2375 10257
rect 2317 10248 2329 10251
rect 1903 10220 2329 10248
rect 1903 10217 1915 10220
rect 1857 10211 1915 10217
rect 2317 10217 2329 10220
rect 2363 10217 2375 10251
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 2317 10211 2375 10217
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 3384 10220 3617 10248
rect 3384 10208 3390 10220
rect 3605 10217 3617 10220
rect 3651 10217 3663 10251
rect 3605 10211 3663 10217
rect 3973 10251 4031 10257
rect 3973 10217 3985 10251
rect 4019 10248 4031 10251
rect 4062 10248 4068 10260
rect 4019 10220 4068 10248
rect 4019 10217 4031 10220
rect 3973 10211 4031 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4338 10208 4344 10260
rect 4396 10248 4402 10260
rect 4433 10251 4491 10257
rect 4433 10248 4445 10251
rect 4396 10220 4445 10248
rect 4396 10208 4402 10220
rect 4433 10217 4445 10220
rect 4479 10217 4491 10251
rect 4433 10211 4491 10217
rect 5537 10251 5595 10257
rect 5537 10217 5549 10251
rect 5583 10217 5595 10251
rect 5537 10211 5595 10217
rect 2866 10180 2872 10192
rect 1688 10152 2872 10180
rect 1688 10056 1716 10152
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 3786 10140 3792 10192
rect 3844 10180 3850 10192
rect 4893 10183 4951 10189
rect 4893 10180 4905 10183
rect 3844 10152 4905 10180
rect 3844 10140 3850 10152
rect 4893 10149 4905 10152
rect 4939 10149 4951 10183
rect 4893 10143 4951 10149
rect 4982 10140 4988 10192
rect 5040 10180 5046 10192
rect 5261 10183 5319 10189
rect 5261 10180 5273 10183
rect 5040 10152 5273 10180
rect 5040 10140 5046 10152
rect 5261 10149 5273 10152
rect 5307 10149 5319 10183
rect 5261 10143 5319 10149
rect 5552 10124 5580 10211
rect 6454 10208 6460 10260
rect 6512 10248 6518 10260
rect 6549 10251 6607 10257
rect 6549 10248 6561 10251
rect 6512 10220 6561 10248
rect 6512 10208 6518 10220
rect 6549 10217 6561 10220
rect 6595 10217 6607 10251
rect 6549 10211 6607 10217
rect 7009 10251 7067 10257
rect 7009 10217 7021 10251
rect 7055 10248 7067 10251
rect 7561 10251 7619 10257
rect 7561 10248 7573 10251
rect 7055 10220 7573 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 7561 10217 7573 10220
rect 7607 10217 7619 10251
rect 7561 10211 7619 10217
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10248 7987 10251
rect 8202 10248 8208 10260
rect 7975 10220 8208 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 8389 10251 8447 10257
rect 8389 10248 8401 10251
rect 8352 10220 8401 10248
rect 8352 10208 8358 10220
rect 8389 10217 8401 10220
rect 8435 10248 8447 10251
rect 9582 10248 9588 10260
rect 8435 10220 9588 10248
rect 8435 10217 8447 10220
rect 8389 10211 8447 10217
rect 9582 10208 9588 10220
rect 9640 10208 9646 10260
rect 10962 10248 10968 10260
rect 10923 10220 10968 10248
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11517 10251 11575 10257
rect 11517 10248 11529 10251
rect 11256 10220 11529 10248
rect 5994 10140 6000 10192
rect 6052 10180 6058 10192
rect 6365 10183 6423 10189
rect 6365 10180 6377 10183
rect 6052 10152 6377 10180
rect 6052 10140 6058 10152
rect 6365 10149 6377 10152
rect 6411 10149 6423 10183
rect 6365 10143 6423 10149
rect 6914 10140 6920 10192
rect 6972 10180 6978 10192
rect 8021 10183 8079 10189
rect 8021 10180 8033 10183
rect 6972 10152 8033 10180
rect 6972 10140 6978 10152
rect 8021 10149 8033 10152
rect 8067 10149 8079 10183
rect 8021 10143 8079 10149
rect 10873 10183 10931 10189
rect 10873 10149 10885 10183
rect 10919 10180 10931 10183
rect 11256 10180 11284 10220
rect 11517 10217 11529 10220
rect 11563 10248 11575 10251
rect 11790 10248 11796 10260
rect 11563 10220 11796 10248
rect 11563 10217 11575 10220
rect 11517 10211 11575 10217
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 14090 10248 14096 10260
rect 11931 10220 14096 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 14090 10208 14096 10220
rect 14148 10208 14154 10260
rect 14461 10251 14519 10257
rect 14461 10217 14473 10251
rect 14507 10248 14519 10251
rect 14550 10248 14556 10260
rect 14507 10220 14556 10248
rect 14507 10217 14519 10220
rect 14461 10211 14519 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 15286 10248 15292 10260
rect 15247 10220 15292 10248
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 15654 10248 15660 10260
rect 15615 10220 15660 10248
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 16117 10251 16175 10257
rect 16117 10217 16129 10251
rect 16163 10248 16175 10251
rect 16482 10248 16488 10260
rect 16163 10220 16488 10248
rect 16163 10217 16175 10220
rect 16117 10211 16175 10217
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 17221 10251 17279 10257
rect 17221 10217 17233 10251
rect 17267 10248 17279 10251
rect 17310 10248 17316 10260
rect 17267 10220 17316 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 17405 10251 17463 10257
rect 17405 10217 17417 10251
rect 17451 10248 17463 10251
rect 17954 10248 17960 10260
rect 17451 10220 17960 10248
rect 17451 10217 17463 10220
rect 17405 10211 17463 10217
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 18966 10248 18972 10260
rect 18927 10220 18972 10248
rect 18966 10208 18972 10220
rect 19024 10208 19030 10260
rect 19058 10208 19064 10260
rect 19116 10248 19122 10260
rect 19153 10251 19211 10257
rect 19153 10248 19165 10251
rect 19116 10220 19165 10248
rect 19116 10208 19122 10220
rect 19153 10217 19165 10220
rect 19199 10217 19211 10251
rect 19153 10211 19211 10217
rect 20993 10251 21051 10257
rect 20993 10217 21005 10251
rect 21039 10217 21051 10251
rect 20993 10211 21051 10217
rect 12158 10180 12164 10192
rect 10919 10152 11284 10180
rect 11348 10152 12164 10180
rect 10919 10149 10931 10152
rect 10873 10143 10931 10149
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 3142 10112 3148 10124
rect 2731 10084 3148 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 3142 10072 3148 10084
rect 3200 10072 3206 10124
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 3418 10112 3424 10124
rect 3375 10084 3424 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10112 4859 10115
rect 4847 10084 5396 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10044 1823 10047
rect 2130 10044 2136 10056
rect 1811 10016 2136 10044
rect 1811 10013 1823 10016
rect 1765 10007 1823 10013
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 2498 10004 2504 10056
rect 2556 10044 2562 10056
rect 2777 10047 2835 10053
rect 2777 10044 2789 10047
rect 2556 10016 2789 10044
rect 2556 10004 2562 10016
rect 2777 10013 2789 10016
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10013 2927 10047
rect 4522 10044 4528 10056
rect 2869 10007 2927 10013
rect 4172 10016 4528 10044
rect 2222 9976 2228 9988
rect 2183 9948 2228 9976
rect 2222 9936 2228 9948
rect 2280 9936 2286 9988
rect 2590 9936 2596 9988
rect 2648 9976 2654 9988
rect 2884 9976 2912 10007
rect 2648 9948 2912 9976
rect 2648 9936 2654 9948
rect 3418 9908 3424 9920
rect 3379 9880 3424 9908
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 4172 9917 4200 10016
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10044 5135 10047
rect 5258 10044 5264 10056
rect 5123 10016 5264 10044
rect 5123 10013 5135 10016
rect 5077 10007 5135 10013
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5368 10044 5396 10084
rect 5534 10072 5540 10124
rect 5592 10072 5598 10124
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10112 5963 10115
rect 6270 10112 6276 10124
rect 5951 10084 6276 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 7098 10112 7104 10124
rect 7059 10084 7104 10112
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 8036 10112 8064 10143
rect 8036 10084 9536 10112
rect 5810 10044 5816 10056
rect 5368 10016 5816 10044
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 5994 10044 6000 10056
rect 5955 10016 6000 10044
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6086 10004 6092 10056
rect 6144 10044 6150 10056
rect 6917 10047 6975 10053
rect 6144 10016 6189 10044
rect 6144 10004 6150 10016
rect 6917 10013 6929 10047
rect 6963 10044 6975 10047
rect 7190 10044 7196 10056
rect 6963 10016 7196 10044
rect 6963 10013 6975 10016
rect 6917 10007 6975 10013
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7650 10004 7656 10056
rect 7708 10044 7714 10056
rect 8113 10047 8171 10053
rect 8113 10044 8125 10047
rect 7708 10016 8125 10044
rect 7708 10004 7714 10016
rect 8113 10013 8125 10016
rect 8159 10044 8171 10047
rect 8202 10044 8208 10056
rect 8159 10016 8208 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9214 10044 9220 10056
rect 8312 10016 9220 10044
rect 4246 9936 4252 9988
rect 4304 9976 4310 9988
rect 4341 9979 4399 9985
rect 4341 9976 4353 9979
rect 4304 9948 4353 9976
rect 4304 9936 4310 9948
rect 4341 9945 4353 9948
rect 4387 9976 4399 9979
rect 8312 9976 8340 10016
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 4387 9948 8340 9976
rect 4387 9945 4399 9948
rect 4341 9939 4399 9945
rect 8478 9936 8484 9988
rect 8536 9976 8542 9988
rect 8757 9979 8815 9985
rect 8757 9976 8769 9979
rect 8536 9948 8769 9976
rect 8536 9936 8542 9948
rect 8757 9945 8769 9948
rect 8803 9976 8815 9979
rect 9306 9976 9312 9988
rect 8803 9948 9312 9976
rect 8803 9945 8815 9948
rect 8757 9939 8815 9945
rect 9306 9936 9312 9948
rect 9364 9936 9370 9988
rect 4157 9911 4215 9917
rect 4157 9877 4169 9911
rect 4203 9908 4215 9911
rect 7006 9908 7012 9920
rect 4203 9880 7012 9908
rect 4203 9877 4215 9880
rect 4157 9871 4215 9877
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9908 7527 9911
rect 7558 9908 7564 9920
rect 7515 9880 7564 9908
rect 7515 9877 7527 9880
rect 7469 9871 7527 9877
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 8018 9868 8024 9920
rect 8076 9908 8082 9920
rect 8294 9908 8300 9920
rect 8076 9880 8300 9908
rect 8076 9868 8082 9880
rect 8294 9868 8300 9880
rect 8352 9908 8358 9920
rect 8573 9911 8631 9917
rect 8573 9908 8585 9911
rect 8352 9880 8585 9908
rect 8352 9868 8358 9880
rect 8573 9877 8585 9880
rect 8619 9877 8631 9911
rect 8573 9871 8631 9877
rect 9125 9911 9183 9917
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9214 9908 9220 9920
rect 9171 9880 9220 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 9508 9908 9536 10084
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 10238 10115 10296 10121
rect 10238 10112 10250 10115
rect 9824 10084 10250 10112
rect 9824 10072 9830 10084
rect 10238 10081 10250 10084
rect 10284 10112 10296 10115
rect 10284 10084 10732 10112
rect 10284 10081 10296 10084
rect 10238 10075 10296 10081
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10044 10563 10047
rect 10594 10044 10600 10056
rect 10551 10016 10600 10044
rect 10551 10013 10563 10016
rect 10505 10007 10563 10013
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 10704 10053 10732 10084
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10013 10747 10047
rect 10689 10007 10747 10013
rect 10962 10004 10968 10056
rect 11020 10044 11026 10056
rect 11348 10044 11376 10152
rect 12158 10140 12164 10152
rect 12216 10140 12222 10192
rect 12526 10140 12532 10192
rect 12584 10180 12590 10192
rect 14001 10183 14059 10189
rect 14001 10180 14013 10183
rect 12584 10152 14013 10180
rect 12584 10140 12590 10152
rect 14001 10149 14013 10152
rect 14047 10180 14059 10183
rect 16577 10183 16635 10189
rect 16577 10180 16589 10183
rect 14047 10152 16589 10180
rect 14047 10149 14059 10152
rect 14001 10143 14059 10149
rect 16577 10149 16589 10152
rect 16623 10149 16635 10183
rect 16577 10143 16635 10149
rect 17586 10140 17592 10192
rect 17644 10180 17650 10192
rect 18540 10183 18598 10189
rect 18540 10180 18552 10183
rect 17644 10152 18552 10180
rect 17644 10140 17650 10152
rect 18540 10149 18552 10152
rect 18586 10180 18598 10183
rect 21008 10180 21036 10211
rect 18586 10152 19564 10180
rect 18586 10149 18598 10152
rect 18540 10143 18598 10149
rect 11977 10115 12035 10121
rect 11977 10081 11989 10115
rect 12023 10112 12035 10115
rect 13262 10112 13268 10124
rect 12023 10084 13268 10112
rect 12023 10081 12035 10084
rect 11977 10075 12035 10081
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13538 10072 13544 10124
rect 13596 10121 13602 10124
rect 13596 10112 13608 10121
rect 13596 10084 13641 10112
rect 13596 10075 13608 10084
rect 13596 10072 13602 10075
rect 13722 10072 13728 10124
rect 13780 10112 13786 10124
rect 13817 10115 13875 10121
rect 13817 10112 13829 10115
rect 13780 10084 13829 10112
rect 13780 10072 13786 10084
rect 13817 10081 13829 10084
rect 13863 10081 13875 10115
rect 13817 10075 13875 10081
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 13964 10084 14105 10112
rect 13964 10072 13970 10084
rect 14093 10081 14105 10084
rect 14139 10112 14151 10115
rect 14829 10115 14887 10121
rect 14829 10112 14841 10115
rect 14139 10084 14841 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 14829 10081 14841 10084
rect 14875 10112 14887 10115
rect 15470 10112 15476 10124
rect 14875 10084 15476 10112
rect 14875 10081 14887 10084
rect 14829 10075 14887 10081
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 15746 10112 15752 10124
rect 15659 10084 15752 10112
rect 15746 10072 15752 10084
rect 15804 10112 15810 10124
rect 15804 10084 16252 10112
rect 15804 10072 15810 10084
rect 11020 10016 11376 10044
rect 11793 10047 11851 10053
rect 11020 10004 11026 10016
rect 11793 10013 11805 10047
rect 11839 10044 11851 10047
rect 11839 10016 12296 10044
rect 11839 10013 11851 10016
rect 11793 10007 11851 10013
rect 11238 9976 11244 9988
rect 10888 9948 11244 9976
rect 10888 9908 10916 9948
rect 11238 9936 11244 9948
rect 11296 9936 11302 9988
rect 9508 9880 10916 9908
rect 10962 9868 10968 9920
rect 11020 9908 11026 9920
rect 11333 9911 11391 9917
rect 11333 9908 11345 9911
rect 11020 9880 11345 9908
rect 11020 9868 11026 9880
rect 11333 9877 11345 9880
rect 11379 9877 11391 9911
rect 12268 9908 12296 10016
rect 13998 10004 14004 10056
rect 14056 10044 14062 10056
rect 14734 10044 14740 10056
rect 14056 10016 14740 10044
rect 14056 10004 14062 10016
rect 14734 10004 14740 10016
rect 14792 10044 14798 10056
rect 14921 10047 14979 10053
rect 14921 10044 14933 10047
rect 14792 10016 14933 10044
rect 14792 10004 14798 10016
rect 14921 10013 14933 10016
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 15013 10047 15071 10053
rect 15013 10013 15025 10047
rect 15059 10013 15071 10047
rect 15013 10007 15071 10013
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10013 15899 10047
rect 16224 10044 16252 10084
rect 16298 10072 16304 10124
rect 16356 10112 16362 10124
rect 16485 10115 16543 10121
rect 16485 10112 16497 10115
rect 16356 10084 16497 10112
rect 16356 10072 16362 10084
rect 16485 10081 16497 10084
rect 16531 10081 16543 10115
rect 19334 10112 19340 10124
rect 16485 10075 16543 10081
rect 16684 10084 19340 10112
rect 16684 10044 16712 10084
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 19536 10112 19564 10152
rect 19720 10152 21036 10180
rect 19720 10112 19748 10152
rect 19886 10121 19892 10124
rect 19880 10112 19892 10121
rect 19536 10084 19748 10112
rect 19799 10084 19892 10112
rect 19880 10075 19892 10084
rect 19944 10112 19950 10124
rect 20438 10112 20444 10124
rect 19944 10084 20444 10112
rect 19886 10072 19892 10075
rect 19944 10072 19950 10084
rect 20438 10072 20444 10084
rect 20496 10072 20502 10124
rect 21177 10115 21235 10121
rect 21177 10081 21189 10115
rect 21223 10112 21235 10115
rect 21545 10115 21603 10121
rect 21545 10112 21557 10115
rect 21223 10084 21557 10112
rect 21223 10081 21235 10084
rect 21177 10075 21235 10081
rect 21545 10081 21557 10084
rect 21591 10112 21603 10115
rect 21634 10112 21640 10124
rect 21591 10084 21640 10112
rect 21591 10081 21603 10084
rect 21545 10075 21603 10081
rect 21634 10072 21640 10084
rect 21692 10072 21698 10124
rect 16224 10016 16712 10044
rect 16761 10047 16819 10053
rect 15841 10007 15899 10013
rect 16761 10013 16773 10047
rect 16807 10044 16819 10047
rect 17586 10044 17592 10056
rect 16807 10016 17592 10044
rect 16807 10013 16819 10016
rect 16761 10007 16819 10013
rect 12345 9979 12403 9985
rect 12345 9945 12357 9979
rect 12391 9976 12403 9979
rect 12391 9948 12949 9976
rect 12391 9945 12403 9948
rect 12345 9939 12403 9945
rect 12437 9911 12495 9917
rect 12437 9908 12449 9911
rect 12268 9880 12449 9908
rect 11333 9871 11391 9877
rect 12437 9877 12449 9880
rect 12483 9908 12495 9911
rect 12710 9908 12716 9920
rect 12483 9880 12716 9908
rect 12483 9877 12495 9880
rect 12437 9871 12495 9877
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 12921 9908 12949 9948
rect 14274 9936 14280 9988
rect 14332 9976 14338 9988
rect 15028 9976 15056 10007
rect 15856 9976 15884 10007
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 18785 10047 18843 10053
rect 18785 10013 18797 10047
rect 18831 10044 18843 10047
rect 19058 10044 19064 10056
rect 18831 10016 19064 10044
rect 18831 10013 18843 10016
rect 18785 10007 18843 10013
rect 19058 10004 19064 10016
rect 19116 10044 19122 10056
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 19116 10016 19625 10044
rect 19116 10004 19122 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 19613 10007 19671 10013
rect 21358 9976 21364 9988
rect 14332 9948 15884 9976
rect 21319 9948 21364 9976
rect 14332 9936 14338 9948
rect 21358 9936 21364 9948
rect 21416 9936 21422 9988
rect 14826 9908 14832 9920
rect 12921 9880 14832 9908
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 15654 9868 15660 9920
rect 15712 9908 15718 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 15712 9880 16957 9908
rect 15712 9868 15718 9880
rect 16945 9877 16957 9880
rect 16991 9908 17003 9911
rect 19242 9908 19248 9920
rect 16991 9880 19248 9908
rect 16991 9877 17003 9880
rect 16945 9871 17003 9877
rect 19242 9868 19248 9880
rect 19300 9868 19306 9920
rect 19426 9908 19432 9920
rect 19387 9880 19432 9908
rect 19426 9868 19432 9880
rect 19484 9868 19490 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 1581 9707 1639 9713
rect 1581 9673 1593 9707
rect 1627 9704 1639 9707
rect 1762 9704 1768 9716
rect 1627 9676 1768 9704
rect 1627 9673 1639 9676
rect 1581 9667 1639 9673
rect 1762 9664 1768 9676
rect 1820 9664 1826 9716
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 4709 9707 4767 9713
rect 4709 9704 4721 9707
rect 3844 9676 4721 9704
rect 3844 9664 3850 9676
rect 4709 9673 4721 9676
rect 4755 9673 4767 9707
rect 4709 9667 4767 9673
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 10502 9704 10508 9716
rect 6604 9676 6776 9704
rect 6604 9664 6610 9676
rect 2682 9596 2688 9648
rect 2740 9636 2746 9648
rect 3970 9636 3976 9648
rect 2740 9608 3976 9636
rect 2740 9596 2746 9608
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 6273 9639 6331 9645
rect 6273 9605 6285 9639
rect 6319 9636 6331 9639
rect 6457 9639 6515 9645
rect 6457 9636 6469 9639
rect 6319 9608 6469 9636
rect 6319 9605 6331 9608
rect 6273 9599 6331 9605
rect 6457 9605 6469 9608
rect 6503 9636 6515 9639
rect 6638 9636 6644 9648
rect 6503 9608 6644 9636
rect 6503 9605 6515 9608
rect 6457 9599 6515 9605
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 6748 9636 6776 9676
rect 7576 9676 10088 9704
rect 10463 9676 10508 9704
rect 7576 9636 7604 9676
rect 8938 9636 8944 9648
rect 6748 9608 7604 9636
rect 8899 9608 8944 9636
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 10060 9636 10088 9676
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 12158 9704 12164 9716
rect 11440 9676 12164 9704
rect 10060 9608 10824 9636
rect 1670 9528 1676 9580
rect 1728 9568 1734 9580
rect 2133 9571 2191 9577
rect 2133 9568 2145 9571
rect 1728 9540 2145 9568
rect 1728 9528 1734 9540
rect 2133 9537 2145 9540
rect 2179 9537 2191 9571
rect 2133 9531 2191 9537
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 2961 9571 3019 9577
rect 2961 9568 2973 9571
rect 2648 9540 2973 9568
rect 2648 9528 2654 9540
rect 2961 9537 2973 9540
rect 3007 9537 3019 9571
rect 4154 9568 4160 9580
rect 4115 9540 4160 9568
rect 2961 9531 3019 9537
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9568 4307 9571
rect 5074 9568 5080 9580
rect 4295 9540 5080 9568
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 7466 9568 7472 9580
rect 6104 9540 7472 9568
rect 6104 9512 6132 9540
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9568 8539 9571
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 8527 9540 9137 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9537 10747 9571
rect 10796 9568 10824 9608
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 11440 9645 11468 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12434 9664 12440 9716
rect 12492 9704 12498 9716
rect 12492 9676 13124 9704
rect 12492 9664 12498 9676
rect 11425 9639 11483 9645
rect 11425 9636 11437 9639
rect 11296 9608 11437 9636
rect 11296 9596 11302 9608
rect 11425 9605 11437 9608
rect 11471 9605 11483 9639
rect 13096 9636 13124 9676
rect 13170 9664 13176 9716
rect 13228 9704 13234 9716
rect 13228 9676 14596 9704
rect 13228 9664 13234 9676
rect 14568 9648 14596 9676
rect 16316 9676 17080 9704
rect 13998 9636 14004 9648
rect 13096 9608 14004 9636
rect 11425 9599 11483 9605
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 14274 9636 14280 9648
rect 14108 9608 14280 9636
rect 11974 9568 11980 9580
rect 10796 9540 11980 9568
rect 10689 9531 10747 9537
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 2866 9500 2872 9512
rect 2823 9472 2872 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 3234 9500 3240 9512
rect 3195 9472 3240 9500
rect 3234 9460 3240 9472
rect 3292 9500 3298 9512
rect 3789 9503 3847 9509
rect 3789 9500 3801 9503
rect 3292 9472 3801 9500
rect 3292 9460 3298 9472
rect 3789 9469 3801 9472
rect 3835 9469 3847 9503
rect 3789 9463 3847 9469
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9500 4399 9503
rect 5442 9500 5448 9512
rect 4387 9472 5448 9500
rect 4387 9469 4399 9472
rect 4341 9463 4399 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5925 9503 5983 9509
rect 5925 9469 5937 9503
rect 5971 9500 5983 9503
rect 6086 9500 6092 9512
rect 5971 9472 6092 9500
rect 5971 9469 5983 9472
rect 5925 9463 5983 9469
rect 6086 9460 6092 9472
rect 6144 9460 6150 9512
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 6273 9503 6331 9509
rect 6273 9500 6285 9503
rect 6227 9472 6285 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 6273 9469 6285 9472
rect 6319 9469 6331 9503
rect 6638 9500 6644 9512
rect 6551 9472 6644 9500
rect 6273 9463 6331 9469
rect 1949 9435 2007 9441
rect 1949 9401 1961 9435
rect 1995 9432 2007 9435
rect 3510 9432 3516 9444
rect 1995 9404 2452 9432
rect 1995 9401 2007 9404
rect 1949 9395 2007 9401
rect 1486 9364 1492 9376
rect 1447 9336 1492 9364
rect 1486 9324 1492 9336
rect 1544 9324 1550 9376
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 2314 9364 2320 9376
rect 2087 9336 2320 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 2424 9373 2452 9404
rect 3436 9404 3516 9432
rect 2409 9367 2467 9373
rect 2409 9333 2421 9367
rect 2455 9333 2467 9367
rect 2409 9327 2467 9333
rect 2869 9367 2927 9373
rect 2869 9333 2881 9367
rect 2915 9364 2927 9367
rect 3050 9364 3056 9376
rect 2915 9336 3056 9364
rect 2915 9333 2927 9336
rect 2869 9327 2927 9333
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3436 9373 3464 9404
rect 3510 9392 3516 9404
rect 3568 9432 3574 9444
rect 4062 9432 4068 9444
rect 3568 9404 4068 9432
rect 3568 9392 3574 9404
rect 4062 9392 4068 9404
rect 4120 9392 4126 9444
rect 4890 9392 4896 9444
rect 4948 9432 4954 9444
rect 5258 9432 5264 9444
rect 4948 9404 5264 9432
rect 4948 9392 4954 9404
rect 5258 9392 5264 9404
rect 5316 9392 5322 9444
rect 6196 9432 6224 9463
rect 6638 9460 6644 9472
rect 6696 9500 6702 9512
rect 6696 9472 6960 9500
rect 6696 9460 6702 9472
rect 5940 9404 6224 9432
rect 6932 9432 6960 9472
rect 7006 9460 7012 9512
rect 7064 9500 7070 9512
rect 8757 9503 8815 9509
rect 7064 9472 8708 9500
rect 7064 9460 7070 9472
rect 6932 9404 8064 9432
rect 5940 9376 5968 9404
rect 3421 9367 3479 9373
rect 3421 9333 3433 9367
rect 3467 9333 3479 9367
rect 3602 9364 3608 9376
rect 3563 9336 3608 9364
rect 3421 9327 3479 9333
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 4801 9367 4859 9373
rect 4801 9333 4813 9367
rect 4847 9364 4859 9367
rect 5626 9364 5632 9376
rect 4847 9336 5632 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 5902 9324 5908 9376
rect 5960 9336 5968 9376
rect 5960 9324 5966 9336
rect 6086 9324 6092 9376
rect 6144 9364 6150 9376
rect 6733 9367 6791 9373
rect 6733 9364 6745 9367
rect 6144 9336 6745 9364
rect 6144 9324 6150 9336
rect 6733 9333 6745 9336
rect 6779 9333 6791 9367
rect 7006 9364 7012 9376
rect 6967 9336 7012 9364
rect 6733 9327 6791 9333
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 7101 9367 7159 9373
rect 7101 9333 7113 9367
rect 7147 9364 7159 9367
rect 7190 9364 7196 9376
rect 7147 9336 7196 9364
rect 7147 9333 7159 9336
rect 7101 9327 7159 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 8036 9364 8064 9404
rect 8202 9392 8208 9444
rect 8260 9441 8266 9444
rect 8260 9435 8283 9441
rect 8271 9401 8283 9435
rect 8260 9395 8283 9401
rect 8260 9392 8266 9395
rect 8573 9367 8631 9373
rect 8573 9364 8585 9367
rect 8036 9336 8585 9364
rect 8573 9333 8585 9336
rect 8619 9333 8631 9367
rect 8680 9364 8708 9472
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 9030 9500 9036 9512
rect 8803 9472 9036 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9140 9500 9168 9531
rect 9950 9500 9956 9512
rect 9140 9472 9956 9500
rect 9950 9460 9956 9472
rect 10008 9500 10014 9512
rect 10594 9500 10600 9512
rect 10008 9472 10600 9500
rect 10008 9460 10014 9472
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 9214 9392 9220 9444
rect 9272 9432 9278 9444
rect 9370 9435 9428 9441
rect 9370 9432 9382 9435
rect 9272 9404 9382 9432
rect 9272 9392 9278 9404
rect 9370 9401 9382 9404
rect 9416 9432 9428 9435
rect 10704 9432 10732 9531
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13170 9568 13176 9580
rect 13127 9540 13176 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 13170 9528 13176 9540
rect 13228 9568 13234 9580
rect 13722 9568 13728 9580
rect 13228 9540 13728 9568
rect 13228 9528 13234 9540
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 14108 9577 14136 9608
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 14550 9596 14556 9648
rect 14608 9636 14614 9648
rect 15289 9639 15347 9645
rect 15289 9636 15301 9639
rect 14608 9608 15301 9636
rect 14608 9596 14614 9608
rect 15289 9605 15301 9608
rect 15335 9636 15347 9639
rect 15562 9636 15568 9648
rect 15335 9608 15568 9636
rect 15335 9605 15347 9608
rect 15289 9599 15347 9605
rect 15562 9596 15568 9608
rect 15620 9596 15626 9648
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 16316 9636 16344 9676
rect 15712 9608 16344 9636
rect 16393 9639 16451 9645
rect 15712 9596 15718 9608
rect 16393 9605 16405 9639
rect 16439 9636 16451 9639
rect 16574 9636 16580 9648
rect 16439 9608 16580 9636
rect 16439 9605 16451 9608
rect 16393 9599 16451 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 16942 9636 16948 9648
rect 16903 9608 16948 9636
rect 16942 9596 16948 9608
rect 17000 9596 17006 9648
rect 17052 9636 17080 9676
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18598 9704 18604 9716
rect 18012 9676 18604 9704
rect 18012 9664 18018 9676
rect 18598 9664 18604 9676
rect 18656 9704 18662 9716
rect 18966 9704 18972 9716
rect 18656 9676 18972 9704
rect 18656 9664 18662 9676
rect 18966 9664 18972 9676
rect 19024 9664 19030 9716
rect 19702 9664 19708 9716
rect 19760 9704 19766 9716
rect 20533 9707 20591 9713
rect 20533 9704 20545 9707
rect 19760 9676 20545 9704
rect 19760 9664 19766 9676
rect 20533 9673 20545 9676
rect 20579 9673 20591 9707
rect 20533 9667 20591 9673
rect 18782 9636 18788 9648
rect 17052 9608 18788 9636
rect 18782 9596 18788 9608
rect 18840 9596 18846 9648
rect 20438 9636 20444 9648
rect 20399 9608 20444 9636
rect 20438 9596 20444 9608
rect 20496 9596 20502 9648
rect 14093 9571 14151 9577
rect 14093 9537 14105 9571
rect 14139 9537 14151 9571
rect 14921 9571 14979 9577
rect 14921 9568 14933 9571
rect 14093 9531 14151 9537
rect 14200 9540 14933 9568
rect 10962 9500 10968 9512
rect 10923 9472 10968 9500
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 11606 9460 11612 9512
rect 11664 9500 11670 9512
rect 12986 9500 12992 9512
rect 11664 9472 12992 9500
rect 11664 9460 11670 9472
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 14200 9500 14228 9540
rect 14921 9537 14933 9540
rect 14967 9537 14979 9571
rect 15838 9568 15844 9580
rect 15799 9540 15844 9568
rect 14921 9531 14979 9537
rect 15838 9528 15844 9540
rect 15896 9528 15902 9580
rect 15933 9571 15991 9577
rect 15933 9537 15945 9571
rect 15979 9568 15991 9571
rect 16666 9568 16672 9580
rect 15979 9540 16672 9568
rect 15979 9537 15991 9540
rect 15933 9531 15991 9537
rect 13372 9472 14228 9500
rect 12526 9432 12532 9444
rect 9416 9404 10732 9432
rect 10796 9404 12532 9432
rect 9416 9401 9428 9404
rect 9370 9395 9428 9401
rect 10796 9364 10824 9404
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 12802 9432 12808 9444
rect 12860 9441 12866 9444
rect 12860 9435 12894 9441
rect 12746 9404 12808 9432
rect 12802 9392 12808 9404
rect 12882 9432 12894 9435
rect 13372 9432 13400 9472
rect 14274 9460 14280 9512
rect 14332 9500 14338 9512
rect 14642 9500 14648 9512
rect 14332 9472 14648 9500
rect 14332 9460 14338 9472
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 14737 9503 14795 9509
rect 14737 9469 14749 9503
rect 14783 9500 14795 9503
rect 15194 9500 15200 9512
rect 14783 9472 15200 9500
rect 14783 9469 14795 9472
rect 14737 9463 14795 9469
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 15948 9500 15976 9531
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 17586 9568 17592 9580
rect 17547 9540 17592 9568
rect 17586 9528 17592 9540
rect 17644 9528 17650 9580
rect 18417 9571 18475 9577
rect 18417 9537 18429 9571
rect 18463 9568 18475 9571
rect 21082 9568 21088 9580
rect 18463 9540 19196 9568
rect 18463 9537 18475 9540
rect 18417 9531 18475 9537
rect 15611 9472 15976 9500
rect 16025 9503 16083 9509
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 16025 9469 16037 9503
rect 16071 9500 16083 9503
rect 16114 9500 16120 9512
rect 16071 9472 16120 9500
rect 16071 9469 16083 9472
rect 16025 9463 16083 9469
rect 16114 9460 16120 9472
rect 16172 9500 16178 9512
rect 16485 9503 16543 9509
rect 16485 9500 16497 9503
rect 16172 9472 16497 9500
rect 16172 9460 16178 9472
rect 16485 9469 16497 9472
rect 16531 9469 16543 9503
rect 16758 9500 16764 9512
rect 16671 9472 16764 9500
rect 16485 9463 16543 9469
rect 16758 9460 16764 9472
rect 16816 9500 16822 9512
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 16816 9472 17417 9500
rect 16816 9460 16822 9472
rect 17405 9469 17417 9472
rect 17451 9500 17463 9503
rect 18141 9503 18199 9509
rect 18141 9500 18153 9503
rect 17451 9472 18153 9500
rect 17451 9469 17463 9472
rect 17405 9463 17463 9469
rect 18141 9469 18153 9472
rect 18187 9500 18199 9503
rect 18690 9500 18696 9512
rect 18187 9472 18696 9500
rect 18187 9469 18199 9472
rect 18141 9463 18199 9469
rect 18690 9460 18696 9472
rect 18748 9460 18754 9512
rect 19058 9500 19064 9512
rect 19019 9472 19064 9500
rect 19058 9460 19064 9472
rect 19116 9460 19122 9512
rect 19168 9500 19196 9540
rect 20180 9540 21088 9568
rect 19328 9503 19386 9509
rect 19328 9500 19340 9503
rect 19168 9472 19340 9500
rect 19328 9469 19340 9472
rect 19374 9500 19386 9503
rect 20180 9500 20208 9540
rect 21082 9528 21088 9540
rect 21140 9568 21146 9580
rect 21177 9571 21235 9577
rect 21177 9568 21189 9571
rect 21140 9540 21189 9568
rect 21140 9528 21146 9540
rect 21177 9537 21189 9540
rect 21223 9537 21235 9571
rect 21177 9531 21235 9537
rect 21542 9500 21548 9512
rect 19374 9472 20208 9500
rect 21503 9472 21548 9500
rect 19374 9469 19386 9472
rect 19328 9463 19386 9469
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 13909 9435 13967 9441
rect 13909 9432 13921 9435
rect 12882 9404 13400 9432
rect 13464 9404 13921 9432
rect 12882 9401 12894 9404
rect 12860 9395 12894 9401
rect 12860 9392 12866 9395
rect 8680 9336 10824 9364
rect 10873 9367 10931 9373
rect 8573 9327 8631 9333
rect 10873 9333 10885 9367
rect 10919 9364 10931 9367
rect 10962 9364 10968 9376
rect 10919 9336 10968 9364
rect 10919 9333 10931 9336
rect 10873 9327 10931 9333
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11146 9324 11152 9376
rect 11204 9364 11210 9376
rect 11333 9367 11391 9373
rect 11333 9364 11345 9367
rect 11204 9336 11345 9364
rect 11204 9324 11210 9336
rect 11333 9333 11345 9336
rect 11379 9333 11391 9367
rect 11698 9364 11704 9376
rect 11659 9336 11704 9364
rect 11333 9327 11391 9333
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13173 9367 13231 9373
rect 13173 9364 13185 9367
rect 13136 9336 13185 9364
rect 13136 9324 13142 9336
rect 13173 9333 13185 9336
rect 13219 9333 13231 9367
rect 13354 9364 13360 9376
rect 13315 9336 13360 9364
rect 13173 9327 13231 9333
rect 13354 9324 13360 9336
rect 13412 9364 13418 9376
rect 13464 9364 13492 9404
rect 13909 9401 13921 9404
rect 13955 9401 13967 9435
rect 13909 9395 13967 9401
rect 14001 9435 14059 9441
rect 14001 9401 14013 9435
rect 14047 9432 14059 9435
rect 14550 9432 14556 9444
rect 14047 9404 14556 9432
rect 14047 9401 14059 9404
rect 14001 9395 14059 9401
rect 14550 9392 14556 9404
rect 14608 9392 14614 9444
rect 14826 9432 14832 9444
rect 14787 9404 14832 9432
rect 14826 9392 14832 9404
rect 14884 9392 14890 9444
rect 17954 9432 17960 9444
rect 17144 9404 17960 9432
rect 13412 9336 13492 9364
rect 13541 9367 13599 9373
rect 13412 9324 13418 9336
rect 13541 9333 13553 9367
rect 13587 9364 13599 9367
rect 13722 9364 13728 9376
rect 13587 9336 13728 9364
rect 13587 9333 13599 9336
rect 13541 9327 13599 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 14369 9367 14427 9373
rect 14369 9333 14381 9367
rect 14415 9364 14427 9367
rect 14642 9364 14648 9376
rect 14415 9336 14648 9364
rect 14415 9333 14427 9336
rect 14369 9327 14427 9333
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 17144 9364 17172 9404
rect 17954 9392 17960 9404
rect 18012 9392 18018 9444
rect 18601 9435 18659 9441
rect 18601 9401 18613 9435
rect 18647 9432 18659 9435
rect 20254 9432 20260 9444
rect 18647 9404 20260 9432
rect 18647 9401 18659 9404
rect 18601 9395 18659 9401
rect 20254 9392 20260 9404
rect 20312 9392 20318 9444
rect 17310 9364 17316 9376
rect 15528 9336 17172 9364
rect 17271 9336 17316 9364
rect 15528 9324 15534 9336
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 18506 9364 18512 9376
rect 18467 9336 18512 9364
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 18969 9367 19027 9373
rect 18969 9333 18981 9367
rect 19015 9364 19027 9367
rect 19794 9364 19800 9376
rect 19015 9336 19800 9364
rect 19015 9333 19027 9336
rect 18969 9327 19027 9333
rect 19794 9324 19800 9336
rect 19852 9324 19858 9376
rect 20898 9364 20904 9376
rect 20859 9336 20904 9364
rect 20898 9324 20904 9336
rect 20956 9324 20962 9376
rect 20990 9324 20996 9376
rect 21048 9364 21054 9376
rect 21358 9364 21364 9376
rect 21048 9336 21093 9364
rect 21319 9336 21364 9364
rect 21048 9324 21054 9336
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 2832 9132 2877 9160
rect 2832 9120 2838 9132
rect 3142 9120 3148 9172
rect 3200 9160 3206 9172
rect 3513 9163 3571 9169
rect 3513 9160 3525 9163
rect 3200 9132 3525 9160
rect 3200 9120 3206 9132
rect 3513 9129 3525 9132
rect 3559 9129 3571 9163
rect 5445 9163 5503 9169
rect 5445 9160 5457 9163
rect 3513 9123 3571 9129
rect 3804 9132 5457 9160
rect 1857 9095 1915 9101
rect 1857 9061 1869 9095
rect 1903 9092 1915 9095
rect 3694 9092 3700 9104
rect 1903 9064 3700 9092
rect 1903 9061 1915 9064
rect 1857 9055 1915 9061
rect 3694 9052 3700 9064
rect 3752 9052 3758 9104
rect 1765 9027 1823 9033
rect 1765 8993 1777 9027
rect 1811 9024 1823 9027
rect 2314 9024 2320 9036
rect 1811 8996 2320 9024
rect 1811 8993 1823 8996
rect 1765 8987 1823 8993
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 2682 9024 2688 9036
rect 2643 8996 2688 9024
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 3142 9024 3148 9036
rect 3055 8996 3148 9024
rect 3142 8984 3148 8996
rect 3200 9024 3206 9036
rect 3602 9024 3608 9036
rect 3200 8996 3608 9024
rect 3200 8984 3206 8996
rect 3602 8984 3608 8996
rect 3660 8984 3666 9036
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 2590 8956 2596 8968
rect 1719 8928 2596 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 2590 8916 2596 8928
rect 2648 8956 2654 8968
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2648 8928 2881 8956
rect 2648 8916 2654 8928
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3804 8956 3832 9132
rect 5445 9129 5457 9132
rect 5491 9129 5503 9163
rect 5445 9123 5503 9129
rect 5718 9120 5724 9172
rect 5776 9160 5782 9172
rect 5776 9132 6316 9160
rect 5776 9120 5782 9132
rect 3896 9064 5948 9092
rect 3896 9036 3924 9064
rect 5920 9036 5948 9064
rect 3878 8984 3884 9036
rect 3936 9024 3942 9036
rect 4154 9033 4160 9036
rect 4148 9024 4160 9033
rect 3936 8996 4029 9024
rect 4115 8996 4160 9024
rect 3936 8984 3942 8996
rect 4148 8987 4160 8996
rect 4154 8984 4160 8987
rect 4212 8984 4218 9036
rect 5902 9024 5908 9036
rect 5863 8996 5908 9024
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 6178 9033 6184 9036
rect 6172 9024 6184 9033
rect 6139 8996 6184 9024
rect 6172 8987 6184 8996
rect 6178 8984 6184 8987
rect 6236 8984 6242 9036
rect 6288 9024 6316 9132
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7929 9163 7987 9169
rect 7929 9160 7941 9163
rect 7156 9132 7941 9160
rect 7156 9120 7162 9132
rect 7929 9129 7941 9132
rect 7975 9129 7987 9163
rect 7929 9123 7987 9129
rect 8297 9163 8355 9169
rect 8297 9129 8309 9163
rect 8343 9160 8355 9163
rect 8938 9160 8944 9172
rect 8343 9132 8944 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 10134 9160 10140 9172
rect 9508 9132 10140 9160
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 7745 9095 7803 9101
rect 7745 9092 7757 9095
rect 6972 9064 7757 9092
rect 6972 9052 6978 9064
rect 7745 9061 7757 9064
rect 7791 9092 7803 9095
rect 8389 9095 8447 9101
rect 7791 9064 8156 9092
rect 7791 9061 7803 9064
rect 7745 9055 7803 9061
rect 8128 9036 8156 9064
rect 8389 9061 8401 9095
rect 8435 9092 8447 9095
rect 8754 9092 8760 9104
rect 8435 9064 8760 9092
rect 8435 9061 8447 9064
rect 8389 9055 8447 9061
rect 8754 9052 8760 9064
rect 8812 9052 8818 9104
rect 9508 9092 9536 9132
rect 10134 9120 10140 9132
rect 10192 9160 10198 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 10192 9132 10241 9160
rect 10192 9120 10198 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 10229 9123 10287 9129
rect 10318 9120 10324 9172
rect 10376 9120 10382 9172
rect 10689 9163 10747 9169
rect 10689 9129 10701 9163
rect 10735 9160 10747 9163
rect 10962 9160 10968 9172
rect 10735 9132 10968 9160
rect 10735 9129 10747 9132
rect 10689 9123 10747 9129
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11146 9160 11152 9172
rect 11107 9132 11152 9160
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 11514 9120 11520 9172
rect 11572 9160 11578 9172
rect 12434 9160 12440 9172
rect 11572 9132 12440 9160
rect 11572 9120 11578 9132
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 12713 9163 12771 9169
rect 12713 9160 12725 9163
rect 12584 9132 12725 9160
rect 12584 9120 12590 9132
rect 12713 9129 12725 9132
rect 12759 9160 12771 9163
rect 12897 9163 12955 9169
rect 12897 9160 12909 9163
rect 12759 9132 12909 9160
rect 12759 9129 12771 9132
rect 12713 9123 12771 9129
rect 12897 9129 12909 9132
rect 12943 9129 12955 9163
rect 12897 9123 12955 9129
rect 8864 9064 9536 9092
rect 9585 9095 9643 9101
rect 7469 9027 7527 9033
rect 7469 9024 7481 9027
rect 6288 8996 7481 9024
rect 7469 8993 7481 8996
rect 7515 9024 7527 9027
rect 7926 9024 7932 9036
rect 7515 8996 7932 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 7926 8984 7932 8996
rect 7984 8984 7990 9036
rect 8110 8984 8116 9036
rect 8168 8984 8174 9036
rect 5810 8956 5816 8968
rect 3292 8928 3832 8956
rect 5771 8928 5816 8956
rect 3292 8916 3298 8928
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 8481 8959 8539 8965
rect 8481 8956 8493 8959
rect 8260 8928 8493 8956
rect 8260 8916 8266 8928
rect 8481 8925 8493 8928
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 8754 8956 8760 8968
rect 8628 8928 8760 8956
rect 8628 8916 8634 8928
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 2130 8848 2136 8900
rect 2188 8888 2194 8900
rect 2225 8891 2283 8897
rect 2225 8888 2237 8891
rect 2188 8860 2237 8888
rect 2188 8848 2194 8860
rect 2225 8857 2237 8860
rect 2271 8857 2283 8891
rect 3326 8888 3332 8900
rect 3287 8860 3332 8888
rect 2225 8851 2283 8857
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 4890 8848 4896 8900
rect 4948 8888 4954 8900
rect 5261 8891 5319 8897
rect 5261 8888 5273 8891
rect 4948 8860 5273 8888
rect 4948 8848 4954 8860
rect 5261 8857 5273 8860
rect 5307 8857 5319 8891
rect 5261 8851 5319 8857
rect 7285 8891 7343 8897
rect 7285 8857 7297 8891
rect 7331 8888 7343 8891
rect 7466 8888 7472 8900
rect 7331 8860 7472 8888
rect 7331 8857 7343 8860
rect 7285 8851 7343 8857
rect 7466 8848 7472 8860
rect 7524 8848 7530 8900
rect 8864 8897 8892 9064
rect 9585 9061 9597 9095
rect 9631 9092 9643 9095
rect 9631 9064 10281 9092
rect 9631 9061 9643 9064
rect 9585 9055 9643 9061
rect 9490 9024 9496 9036
rect 9451 8996 9496 9024
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 9600 8996 10180 9024
rect 8938 8916 8944 8968
rect 8996 8956 9002 8968
rect 9600 8956 9628 8996
rect 9766 8956 9772 8968
rect 8996 8928 9628 8956
rect 9727 8928 9772 8956
rect 8996 8916 9002 8928
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 8849 8891 8907 8897
rect 8849 8888 8861 8891
rect 7585 8860 8861 8888
rect 2682 8780 2688 8832
rect 2740 8820 2746 8832
rect 6822 8820 6828 8832
rect 2740 8792 6828 8820
rect 2740 8780 2746 8792
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7585 8820 7613 8860
rect 8849 8857 8861 8860
rect 8895 8857 8907 8891
rect 8849 8851 8907 8857
rect 6972 8792 7613 8820
rect 7653 8823 7711 8829
rect 6972 8780 6978 8792
rect 7653 8789 7665 8823
rect 7699 8820 7711 8823
rect 8202 8820 8208 8832
rect 7699 8792 8208 8820
rect 7699 8789 7711 8792
rect 7653 8783 7711 8789
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 9180 8792 9225 8820
rect 9180 8780 9186 8792
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10060 8820 10088 8919
rect 10152 8888 10180 8996
rect 10253 8956 10281 9064
rect 10336 9033 10364 9120
rect 10410 9052 10416 9104
rect 10468 9092 10474 9104
rect 11606 9092 11612 9104
rect 10468 9064 11612 9092
rect 10468 9052 10474 9064
rect 11606 9052 11612 9064
rect 11664 9052 11670 9104
rect 11974 9052 11980 9104
rect 12032 9092 12038 9104
rect 12069 9095 12127 9101
rect 12069 9092 12081 9095
rect 12032 9064 12081 9092
rect 12032 9052 12038 9064
rect 12069 9061 12081 9064
rect 12115 9092 12127 9095
rect 12912 9092 12940 9123
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 13044 9132 13093 9160
rect 13044 9120 13050 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13262 9160 13268 9172
rect 13223 9132 13268 9160
rect 13081 9123 13139 9129
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 13722 9160 13728 9172
rect 13683 9132 13728 9160
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 14829 9163 14887 9169
rect 14829 9160 14841 9163
rect 13832 9132 14841 9160
rect 13832 9092 13860 9132
rect 14829 9129 14841 9132
rect 14875 9160 14887 9163
rect 15562 9160 15568 9172
rect 14875 9132 15568 9160
rect 14875 9129 14887 9132
rect 14829 9123 14887 9129
rect 15562 9120 15568 9132
rect 15620 9120 15626 9172
rect 17497 9163 17555 9169
rect 17497 9129 17509 9163
rect 17543 9160 17555 9163
rect 17770 9160 17776 9172
rect 17543 9132 17776 9160
rect 17543 9129 17555 9132
rect 17497 9123 17555 9129
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 17865 9163 17923 9169
rect 17865 9129 17877 9163
rect 17911 9160 17923 9163
rect 17911 9132 18460 9160
rect 17911 9129 17923 9132
rect 17865 9123 17923 9129
rect 15654 9092 15660 9104
rect 12115 9064 12572 9092
rect 12912 9064 13860 9092
rect 13924 9064 15660 9092
rect 12115 9061 12127 9064
rect 12069 9055 12127 9061
rect 10321 9027 10379 9033
rect 10321 8993 10333 9027
rect 10367 9024 10379 9027
rect 10594 9024 10600 9036
rect 10367 8996 10600 9024
rect 10367 8993 10379 8996
rect 10321 8987 10379 8993
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11514 9024 11520 9036
rect 11204 8996 11520 9024
rect 11204 8984 11210 8996
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 11882 8984 11888 9036
rect 11940 9024 11946 9036
rect 12158 9024 12164 9036
rect 11940 8996 12164 9024
rect 11940 8984 11946 8996
rect 12158 8984 12164 8996
rect 12216 8984 12222 9036
rect 10410 8956 10416 8968
rect 10253 8928 10416 8956
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 10560 8928 10885 8956
rect 10560 8916 10566 8928
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8925 11115 8959
rect 11057 8919 11115 8925
rect 11072 8888 11100 8919
rect 10152 8860 11100 8888
rect 11517 8891 11575 8897
rect 11517 8857 11529 8891
rect 11563 8888 11575 8891
rect 11882 8888 11888 8900
rect 11563 8860 11888 8888
rect 11563 8857 11575 8860
rect 11517 8851 11575 8857
rect 11882 8848 11888 8860
rect 11940 8848 11946 8900
rect 12437 8891 12495 8897
rect 12437 8857 12449 8891
rect 12483 8888 12495 8891
rect 12544 8888 12572 9064
rect 12802 8984 12808 9036
rect 12860 9024 12866 9036
rect 13354 9024 13360 9036
rect 12860 8996 13360 9024
rect 12860 8984 12866 8996
rect 13354 8984 13360 8996
rect 13412 8984 13418 9036
rect 13630 9024 13636 9036
rect 13591 8996 13636 9024
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 13722 8984 13728 9036
rect 13780 9024 13786 9036
rect 13924 9024 13952 9064
rect 15654 9052 15660 9064
rect 15712 9052 15718 9104
rect 18432 9092 18460 9132
rect 18506 9120 18512 9172
rect 18564 9160 18570 9172
rect 18693 9163 18751 9169
rect 18693 9160 18705 9163
rect 18564 9132 18705 9160
rect 18564 9120 18570 9132
rect 18693 9129 18705 9132
rect 18739 9129 18751 9163
rect 18693 9123 18751 9129
rect 18782 9120 18788 9172
rect 18840 9160 18846 9172
rect 20993 9163 21051 9169
rect 18840 9132 19012 9160
rect 18840 9120 18846 9132
rect 18601 9095 18659 9101
rect 18601 9092 18613 9095
rect 16684 9064 17080 9092
rect 18432 9064 18613 9092
rect 14366 9024 14372 9036
rect 13780 8996 13952 9024
rect 14327 8996 14372 9024
rect 13780 8984 13786 8996
rect 14366 8984 14372 8996
rect 14424 8984 14430 9036
rect 14550 8984 14556 9036
rect 14608 9024 14614 9036
rect 15381 9027 15439 9033
rect 15381 9024 15393 9027
rect 14608 8996 15393 9024
rect 14608 8984 14614 8996
rect 15381 8993 15393 8996
rect 15427 8993 15439 9027
rect 15746 9024 15752 9036
rect 15381 8987 15439 8993
rect 15488 8996 15752 9024
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 13817 8959 13875 8965
rect 13817 8956 13829 8959
rect 13596 8928 13829 8956
rect 13596 8916 13602 8928
rect 13817 8925 13829 8928
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 15105 8959 15163 8965
rect 15105 8956 15117 8959
rect 14056 8928 15117 8956
rect 14056 8916 14062 8928
rect 15105 8925 15117 8928
rect 15151 8956 15163 8959
rect 15488 8956 15516 8996
rect 15746 8984 15752 8996
rect 15804 8984 15810 9036
rect 16684 9024 16712 9064
rect 16040 8996 16712 9024
rect 15151 8928 15516 8956
rect 15151 8925 15163 8928
rect 15105 8919 15163 8925
rect 12621 8891 12679 8897
rect 12621 8888 12633 8891
rect 12483 8860 12633 8888
rect 12483 8857 12495 8860
rect 12437 8851 12495 8857
rect 12621 8857 12633 8860
rect 12667 8888 12679 8891
rect 13078 8888 13084 8900
rect 12667 8860 13084 8888
rect 12667 8857 12679 8860
rect 12621 8851 12679 8857
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 14185 8891 14243 8897
rect 14185 8857 14197 8891
rect 14231 8888 14243 8891
rect 14231 8860 14780 8888
rect 14231 8857 14243 8860
rect 14185 8851 14243 8857
rect 14752 8832 14780 8860
rect 15470 8848 15476 8900
rect 15528 8888 15534 8900
rect 15565 8891 15623 8897
rect 15565 8888 15577 8891
rect 15528 8860 15577 8888
rect 15528 8848 15534 8860
rect 15565 8857 15577 8860
rect 15611 8888 15623 8891
rect 16040 8888 16068 8996
rect 16758 8984 16764 9036
rect 16816 9033 16822 9036
rect 17052 9033 17080 9064
rect 18601 9061 18613 9064
rect 18647 9061 18659 9095
rect 18984 9092 19012 9132
rect 20993 9129 21005 9163
rect 21039 9160 21051 9163
rect 21082 9160 21088 9172
rect 21039 9132 21088 9160
rect 21039 9129 21051 9132
rect 20993 9123 21051 9129
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 21358 9092 21364 9104
rect 18984 9064 21364 9092
rect 18601 9055 18659 9061
rect 21358 9052 21364 9064
rect 21416 9052 21422 9104
rect 16816 9024 16828 9033
rect 17037 9027 17095 9033
rect 16816 8996 16861 9024
rect 16816 8987 16828 8996
rect 17037 8993 17049 9027
rect 17083 9024 17095 9027
rect 18046 9024 18052 9036
rect 17083 8996 17540 9024
rect 18007 8996 18052 9024
rect 17083 8993 17095 8996
rect 17037 8987 17095 8993
rect 16816 8984 16822 8987
rect 17221 8959 17279 8965
rect 17221 8925 17233 8959
rect 17267 8925 17279 8959
rect 17402 8956 17408 8968
rect 17363 8928 17408 8956
rect 17221 8919 17279 8925
rect 15611 8860 16068 8888
rect 15611 8857 15623 8860
rect 15565 8851 15623 8857
rect 9824 8792 10088 8820
rect 9824 8780 9830 8792
rect 10134 8780 10140 8832
rect 10192 8820 10198 8832
rect 11793 8823 11851 8829
rect 11793 8820 11805 8823
rect 10192 8792 11805 8820
rect 10192 8780 10198 8792
rect 11793 8789 11805 8792
rect 11839 8820 11851 8823
rect 12710 8820 12716 8832
rect 11839 8792 12716 8820
rect 11839 8789 11851 8792
rect 11793 8783 11851 8789
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 14550 8820 14556 8832
rect 14511 8792 14556 8820
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 14734 8820 14740 8832
rect 14695 8792 14740 8820
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 15194 8820 15200 8832
rect 15155 8792 15200 8820
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 15654 8780 15660 8832
rect 15712 8820 15718 8832
rect 17236 8820 17264 8919
rect 17402 8916 17408 8928
rect 17460 8916 17466 8968
rect 17512 8956 17540 8996
rect 18046 8984 18052 8996
rect 18104 9024 18110 9036
rect 18782 9024 18788 9036
rect 18104 8996 18788 9024
rect 18104 8984 18110 8996
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 19058 9024 19064 9036
rect 19019 8996 19064 9024
rect 19058 8984 19064 8996
rect 19116 8984 19122 9036
rect 19153 9027 19211 9033
rect 19153 8993 19165 9027
rect 19199 9024 19211 9027
rect 19426 9024 19432 9036
rect 19199 8996 19432 9024
rect 19199 8993 19211 8996
rect 19153 8987 19211 8993
rect 19426 8984 19432 8996
rect 19484 8984 19490 9036
rect 19886 9033 19892 9036
rect 19880 9024 19892 9033
rect 19536 8996 19892 9024
rect 17954 8956 17960 8968
rect 17512 8928 17960 8956
rect 17954 8916 17960 8928
rect 18012 8956 18018 8968
rect 19337 8959 19395 8965
rect 18012 8928 19012 8956
rect 18012 8916 18018 8928
rect 18984 8900 19012 8928
rect 19337 8925 19349 8959
rect 19383 8956 19395 8959
rect 19536 8956 19564 8996
rect 19880 8987 19892 8996
rect 19886 8984 19892 8987
rect 19944 8984 19950 9036
rect 21177 9027 21235 9033
rect 21177 8993 21189 9027
rect 21223 9024 21235 9027
rect 21542 9024 21548 9036
rect 21223 8996 21548 9024
rect 21223 8993 21235 8996
rect 21177 8987 21235 8993
rect 21542 8984 21548 8996
rect 21600 8984 21606 9036
rect 19383 8928 19564 8956
rect 19613 8959 19671 8965
rect 19383 8925 19395 8928
rect 19337 8919 19395 8925
rect 19613 8925 19625 8959
rect 19659 8925 19671 8959
rect 19613 8919 19671 8925
rect 18230 8888 18236 8900
rect 18191 8860 18236 8888
rect 18230 8848 18236 8860
rect 18288 8848 18294 8900
rect 18966 8848 18972 8900
rect 19024 8888 19030 8900
rect 19628 8888 19656 8919
rect 19024 8860 19656 8888
rect 19024 8848 19030 8860
rect 15712 8792 17264 8820
rect 15712 8780 15718 8792
rect 18138 8780 18144 8832
rect 18196 8820 18202 8832
rect 18417 8823 18475 8829
rect 18417 8820 18429 8823
rect 18196 8792 18429 8820
rect 18196 8780 18202 8792
rect 18417 8789 18429 8792
rect 18463 8789 18475 8823
rect 18417 8783 18475 8789
rect 18601 8823 18659 8829
rect 18601 8789 18613 8823
rect 18647 8820 18659 8823
rect 19334 8820 19340 8832
rect 18647 8792 19340 8820
rect 18647 8789 18659 8792
rect 18601 8783 18659 8789
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 19610 8780 19616 8832
rect 19668 8820 19674 8832
rect 20530 8820 20536 8832
rect 19668 8792 20536 8820
rect 19668 8780 19674 8792
rect 20530 8780 20536 8792
rect 20588 8780 20594 8832
rect 20806 8780 20812 8832
rect 20864 8820 20870 8832
rect 21361 8823 21419 8829
rect 21361 8820 21373 8823
rect 20864 8792 21373 8820
rect 20864 8780 20870 8792
rect 21361 8789 21373 8792
rect 21407 8789 21419 8823
rect 21361 8783 21419 8789
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 1762 8576 1768 8628
rect 1820 8616 1826 8628
rect 1820 8588 3924 8616
rect 1820 8576 1826 8588
rect 1673 8551 1731 8557
rect 1673 8517 1685 8551
rect 1719 8548 1731 8551
rect 1854 8548 1860 8560
rect 1719 8520 1860 8548
rect 1719 8517 1731 8520
rect 1673 8511 1731 8517
rect 1854 8508 1860 8520
rect 1912 8508 1918 8560
rect 1946 8508 1952 8560
rect 2004 8548 2010 8560
rect 3896 8548 3924 8588
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4341 8619 4399 8625
rect 4341 8616 4353 8619
rect 4212 8588 4353 8616
rect 4212 8576 4218 8588
rect 4341 8585 4353 8588
rect 4387 8585 4399 8619
rect 4341 8579 4399 8585
rect 4709 8619 4767 8625
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 4798 8616 4804 8628
rect 4755 8588 4804 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 5626 8576 5632 8628
rect 5684 8576 5690 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6457 8619 6515 8625
rect 6457 8616 6469 8619
rect 6052 8588 6469 8616
rect 6052 8576 6058 8588
rect 6457 8585 6469 8588
rect 6503 8585 6515 8619
rect 6457 8579 6515 8585
rect 8849 8619 8907 8625
rect 8849 8585 8861 8619
rect 8895 8616 8907 8619
rect 8938 8616 8944 8628
rect 8895 8588 8944 8616
rect 8895 8585 8907 8588
rect 8849 8579 8907 8585
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 10594 8616 10600 8628
rect 10192 8588 10600 8616
rect 10192 8576 10198 8588
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 10689 8619 10747 8625
rect 10689 8585 10701 8619
rect 10735 8616 10747 8619
rect 10870 8616 10876 8628
rect 10735 8588 10876 8616
rect 10735 8585 10747 8588
rect 10689 8579 10747 8585
rect 4433 8551 4491 8557
rect 4433 8548 4445 8551
rect 2004 8520 2049 8548
rect 3896 8520 4445 8548
rect 2004 8508 2010 8520
rect 4433 8517 4445 8520
rect 4479 8517 4491 8551
rect 5644 8548 5672 8576
rect 6270 8548 6276 8560
rect 4433 8511 4491 8517
rect 5368 8520 5672 8548
rect 6231 8520 6276 8548
rect 5368 8489 5396 8520
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 9769 8551 9827 8557
rect 7116 8520 7880 8548
rect 7116 8492 7144 8520
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2424 8452 2697 8480
rect 1762 8412 1768 8424
rect 1723 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 1486 8344 1492 8356
rect 1447 8316 1492 8344
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 2424 8344 2452 8452
rect 2685 8449 2697 8452
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 6178 8480 6184 8492
rect 5767 8452 6184 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 6178 8440 6184 8452
rect 6236 8480 6242 8492
rect 7098 8480 7104 8492
rect 6236 8452 7104 8480
rect 6236 8440 6242 8452
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7190 8440 7196 8492
rect 7248 8480 7254 8492
rect 7374 8480 7380 8492
rect 7248 8452 7380 8480
rect 7248 8440 7254 8452
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 7742 8480 7748 8492
rect 7703 8452 7748 8480
rect 7742 8440 7748 8452
rect 7800 8440 7806 8492
rect 7852 8489 7880 8520
rect 8404 8520 9720 8548
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 8294 8480 8300 8492
rect 8255 8452 8300 8480
rect 7837 8443 7895 8449
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8412 2559 8415
rect 2774 8412 2780 8424
rect 2547 8384 2780 8412
rect 2547 8381 2559 8384
rect 2501 8375 2559 8381
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8412 3019 8415
rect 3786 8412 3792 8424
rect 3007 8384 3792 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 3344 8356 3372 8384
rect 3786 8372 3792 8384
rect 3844 8372 3850 8424
rect 5077 8415 5135 8421
rect 5077 8381 5089 8415
rect 5123 8412 5135 8415
rect 5534 8412 5540 8424
rect 5123 8384 5540 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 5810 8372 5816 8424
rect 5868 8412 5874 8424
rect 5905 8415 5963 8421
rect 5905 8412 5917 8415
rect 5868 8384 5917 8412
rect 5868 8372 5874 8384
rect 5905 8381 5917 8384
rect 5951 8381 5963 8415
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 5905 8375 5963 8381
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8412 6975 8415
rect 7006 8412 7012 8424
rect 6963 8384 7012 8412
rect 6963 8381 6975 8384
rect 6917 8375 6975 8381
rect 7006 8372 7012 8384
rect 7064 8412 7070 8424
rect 8404 8412 8432 8520
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 7064 8384 8432 8412
rect 8481 8415 8539 8421
rect 7064 8372 7070 8384
rect 8481 8381 8493 8415
rect 8527 8412 8539 8415
rect 9122 8412 9128 8424
rect 8527 8384 9128 8412
rect 8527 8381 8539 8384
rect 8481 8375 8539 8381
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 9272 8384 9321 8412
rect 9272 8372 9278 8384
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9508 8412 9536 8443
rect 9582 8412 9588 8424
rect 9508 8384 9588 8412
rect 9309 8375 9367 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 9692 8412 9720 8520
rect 9769 8517 9781 8551
rect 9815 8548 9827 8551
rect 10502 8548 10508 8560
rect 9815 8520 10508 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 10410 8480 10416 8492
rect 10371 8452 10416 8480
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10229 8415 10287 8421
rect 9692 8384 10180 8412
rect 2593 8347 2651 8353
rect 2424 8316 2544 8344
rect 2130 8276 2136 8288
rect 2091 8248 2136 8276
rect 2130 8236 2136 8248
rect 2188 8236 2194 8288
rect 2516 8276 2544 8316
rect 2593 8313 2605 8347
rect 2639 8344 2651 8347
rect 2866 8344 2872 8356
rect 2639 8316 2872 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 3050 8304 3056 8356
rect 3108 8344 3114 8356
rect 3206 8347 3264 8353
rect 3206 8344 3218 8347
rect 3108 8316 3218 8344
rect 3108 8304 3114 8316
rect 3206 8313 3218 8316
rect 3252 8313 3264 8347
rect 3206 8307 3264 8313
rect 3326 8304 3332 8356
rect 3384 8304 3390 8356
rect 5169 8347 5227 8353
rect 5169 8313 5181 8347
rect 5215 8344 5227 8347
rect 7098 8344 7104 8356
rect 5215 8316 7104 8344
rect 5215 8313 5227 8316
rect 5169 8307 5227 8313
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 7653 8347 7711 8353
rect 7653 8313 7665 8347
rect 7699 8344 7711 8347
rect 10042 8344 10048 8356
rect 7699 8316 10048 8344
rect 7699 8313 7711 8316
rect 7653 8307 7711 8313
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 10152 8344 10180 8384
rect 10229 8381 10241 8415
rect 10275 8412 10287 8415
rect 10704 8412 10732 8579
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11238 8616 11244 8628
rect 11112 8588 11244 8616
rect 11112 8576 11118 8588
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11517 8619 11575 8625
rect 11517 8585 11529 8619
rect 11563 8616 11575 8619
rect 12526 8616 12532 8628
rect 11563 8588 12532 8616
rect 11563 8585 11575 8588
rect 11517 8579 11575 8585
rect 12526 8576 12532 8588
rect 12584 8576 12590 8628
rect 13262 8616 13268 8628
rect 12636 8588 13268 8616
rect 11701 8551 11759 8557
rect 11701 8548 11713 8551
rect 11072 8520 11713 8548
rect 10962 8480 10968 8492
rect 10923 8452 10968 8480
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 11072 8489 11100 8520
rect 11701 8517 11713 8520
rect 11747 8517 11759 8551
rect 12636 8548 12664 8588
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 15654 8616 15660 8628
rect 15304 8588 15660 8616
rect 11701 8511 11759 8517
rect 11808 8520 12664 8548
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11808 8480 11836 8520
rect 12710 8508 12716 8560
rect 12768 8548 12774 8560
rect 12989 8551 13047 8557
rect 12989 8548 13001 8551
rect 12768 8520 13001 8548
rect 12768 8508 12774 8520
rect 12989 8517 13001 8520
rect 13035 8517 13047 8551
rect 12989 8511 13047 8517
rect 12250 8480 12256 8492
rect 11296 8452 11836 8480
rect 12211 8452 12256 8480
rect 11296 8440 11302 8452
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 13538 8480 13544 8492
rect 13499 8452 13544 8480
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 15304 8480 15332 8588
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 17770 8616 17776 8628
rect 15804 8588 17264 8616
rect 17731 8588 17776 8616
rect 15804 8576 15810 8588
rect 16758 8548 16764 8560
rect 16671 8520 16764 8548
rect 16758 8508 16764 8520
rect 16816 8548 16822 8560
rect 17236 8548 17264 8588
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 20162 8616 20168 8628
rect 19076 8588 20168 8616
rect 18046 8548 18052 8560
rect 16816 8520 17172 8548
rect 17236 8520 18052 8548
rect 16816 8508 16822 8520
rect 15212 8452 15332 8480
rect 17037 8483 17095 8489
rect 12158 8412 12164 8424
rect 10275 8384 10732 8412
rect 12071 8384 12164 8412
rect 10275 8381 10287 8384
rect 10229 8375 10287 8381
rect 12158 8372 12164 8384
rect 12216 8412 12222 8424
rect 12713 8415 12771 8421
rect 12713 8412 12725 8415
rect 12216 8384 12725 8412
rect 12216 8372 12222 8384
rect 12713 8381 12725 8384
rect 12759 8412 12771 8415
rect 13722 8412 13728 8424
rect 12759 8384 13728 8412
rect 12759 8381 12771 8384
rect 12713 8375 12771 8381
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 15033 8415 15091 8421
rect 15033 8381 15045 8415
rect 15079 8412 15091 8415
rect 15212 8412 15240 8452
rect 17037 8449 17049 8483
rect 17083 8449 17095 8483
rect 17144 8480 17172 8520
rect 18046 8508 18052 8520
rect 18104 8508 18110 8560
rect 18325 8483 18383 8489
rect 18325 8480 18337 8483
rect 17144 8452 18337 8480
rect 17037 8443 17095 8449
rect 18325 8449 18337 8452
rect 18371 8449 18383 8483
rect 18325 8443 18383 8449
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8480 18843 8483
rect 18966 8480 18972 8492
rect 18831 8452 18972 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 15079 8384 15240 8412
rect 15289 8415 15347 8421
rect 15079 8381 15091 8384
rect 15033 8375 15091 8381
rect 15289 8381 15301 8415
rect 15335 8412 15347 8415
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 15335 8384 15393 8412
rect 15335 8381 15347 8384
rect 15289 8375 15347 8381
rect 15381 8381 15393 8384
rect 15427 8412 15439 8415
rect 15470 8412 15476 8424
rect 15427 8384 15476 8412
rect 15427 8381 15439 8384
rect 15381 8375 15439 8381
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 17052 8412 17080 8443
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 15856 8384 17080 8412
rect 15856 8356 15884 8384
rect 17678 8372 17684 8424
rect 17736 8412 17742 8424
rect 18877 8415 18935 8421
rect 18877 8412 18889 8415
rect 17736 8384 18889 8412
rect 17736 8372 17742 8384
rect 18877 8381 18889 8384
rect 18923 8381 18935 8415
rect 19076 8412 19104 8588
rect 20162 8576 20168 8588
rect 20220 8576 20226 8628
rect 20441 8619 20499 8625
rect 20441 8585 20453 8619
rect 20487 8616 20499 8619
rect 20898 8616 20904 8628
rect 20487 8588 20904 8616
rect 20487 8585 20499 8588
rect 20441 8579 20499 8585
rect 20898 8576 20904 8588
rect 20956 8576 20962 8628
rect 21361 8551 21419 8557
rect 21361 8548 21373 8551
rect 19306 8520 21373 8548
rect 19306 8480 19334 8520
rect 21361 8517 21373 8520
rect 21407 8517 21419 8551
rect 21361 8511 21419 8517
rect 19886 8480 19892 8492
rect 18877 8375 18935 8381
rect 18984 8384 19104 8412
rect 19168 8452 19334 8480
rect 19847 8452 19892 8480
rect 10870 8344 10876 8356
rect 10152 8316 10876 8344
rect 10870 8304 10876 8316
rect 10928 8304 10934 8356
rect 11149 8347 11207 8353
rect 11149 8313 11161 8347
rect 11195 8344 11207 8347
rect 12434 8344 12440 8356
rect 11195 8316 12440 8344
rect 11195 8313 11207 8316
rect 11149 8307 11207 8313
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 12621 8347 12679 8353
rect 12621 8313 12633 8347
rect 12667 8344 12679 8347
rect 12802 8344 12808 8356
rect 12667 8316 12808 8344
rect 12667 8313 12679 8316
rect 12621 8307 12679 8313
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 12894 8304 12900 8356
rect 12952 8304 12958 8356
rect 14826 8304 14832 8356
rect 14884 8344 14890 8356
rect 15648 8347 15706 8353
rect 14884 8316 14964 8344
rect 14884 8304 14890 8316
rect 3068 8276 3096 8304
rect 2516 8248 3096 8276
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 4890 8276 4896 8288
rect 3476 8248 4896 8276
rect 3476 8236 3482 8248
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 4982 8236 4988 8288
rect 5040 8276 5046 8288
rect 5442 8276 5448 8288
rect 5040 8248 5448 8276
rect 5040 8236 5046 8248
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 5810 8276 5816 8288
rect 5771 8248 5816 8276
rect 5810 8236 5816 8248
rect 5868 8236 5874 8288
rect 7282 8276 7288 8288
rect 7243 8248 7288 8276
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 8386 8276 8392 8288
rect 8347 8248 8392 8276
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 8996 8248 9041 8276
rect 8996 8236 9002 8248
rect 9306 8236 9312 8288
rect 9364 8276 9370 8288
rect 9401 8279 9459 8285
rect 9401 8276 9413 8279
rect 9364 8248 9413 8276
rect 9364 8236 9370 8248
rect 9401 8245 9413 8248
rect 9447 8245 9459 8279
rect 10134 8276 10140 8288
rect 10047 8248 10140 8276
rect 9401 8239 9459 8245
rect 10134 8236 10140 8248
rect 10192 8276 10198 8288
rect 12069 8279 12127 8285
rect 12069 8276 12081 8279
rect 10192 8248 12081 8276
rect 10192 8236 10198 8248
rect 12069 8245 12081 8248
rect 12115 8245 12127 8279
rect 12069 8239 12127 8245
rect 12158 8236 12164 8288
rect 12216 8276 12222 8288
rect 12912 8276 12940 8304
rect 13354 8276 13360 8288
rect 12216 8248 12940 8276
rect 13315 8248 13360 8276
rect 12216 8236 12222 8248
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 13449 8279 13507 8285
rect 13449 8245 13461 8279
rect 13495 8276 13507 8279
rect 13722 8276 13728 8288
rect 13495 8248 13728 8276
rect 13495 8245 13507 8248
rect 13449 8239 13507 8245
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 13909 8279 13967 8285
rect 13909 8245 13921 8279
rect 13955 8276 13967 8279
rect 13998 8276 14004 8288
rect 13955 8248 14004 8276
rect 13955 8245 13967 8248
rect 13909 8239 13967 8245
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 14936 8276 14964 8316
rect 15648 8313 15660 8347
rect 15694 8344 15706 8347
rect 15838 8344 15844 8356
rect 15694 8316 15844 8344
rect 15694 8313 15706 8316
rect 15648 8307 15706 8313
rect 15838 8304 15844 8316
rect 15896 8304 15902 8356
rect 16022 8304 16028 8356
rect 16080 8344 16086 8356
rect 16080 8316 17080 8344
rect 16080 8304 16086 8316
rect 15930 8276 15936 8288
rect 14936 8248 15936 8276
rect 15930 8236 15936 8248
rect 15988 8236 15994 8288
rect 17052 8276 17080 8316
rect 17126 8304 17132 8356
rect 17184 8344 17190 8356
rect 17313 8347 17371 8353
rect 17313 8344 17325 8347
rect 17184 8316 17325 8344
rect 17184 8304 17190 8316
rect 17313 8313 17325 8316
rect 17359 8313 17371 8347
rect 17313 8307 17371 8313
rect 17586 8304 17592 8356
rect 17644 8344 17650 8356
rect 18233 8347 18291 8353
rect 18233 8344 18245 8347
rect 17644 8316 18245 8344
rect 17644 8304 17650 8316
rect 18233 8313 18245 8316
rect 18279 8313 18291 8347
rect 18233 8307 18291 8313
rect 18322 8304 18328 8356
rect 18380 8344 18386 8356
rect 18984 8353 19012 8384
rect 18969 8347 19027 8353
rect 18969 8344 18981 8347
rect 18380 8316 18981 8344
rect 18380 8304 18386 8316
rect 18969 8313 18981 8316
rect 19015 8313 19027 8347
rect 18969 8307 19027 8313
rect 17221 8279 17279 8285
rect 17221 8276 17233 8279
rect 17052 8248 17233 8276
rect 17221 8245 17233 8248
rect 17267 8245 17279 8279
rect 17221 8239 17279 8245
rect 17681 8279 17739 8285
rect 17681 8245 17693 8279
rect 17727 8276 17739 8279
rect 18141 8279 18199 8285
rect 18141 8276 18153 8279
rect 17727 8248 18153 8276
rect 17727 8245 17739 8248
rect 17681 8239 17739 8245
rect 18141 8245 18153 8248
rect 18187 8245 18199 8279
rect 18141 8239 18199 8245
rect 18414 8236 18420 8288
rect 18472 8276 18478 8288
rect 19168 8276 19196 8452
rect 19886 8440 19892 8452
rect 19944 8440 19950 8492
rect 20714 8440 20720 8492
rect 20772 8480 20778 8492
rect 21085 8483 21143 8489
rect 21085 8480 21097 8483
rect 20772 8452 21097 8480
rect 20772 8440 20778 8452
rect 21085 8449 21097 8452
rect 21131 8449 21143 8483
rect 21085 8443 21143 8449
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 19521 8415 19579 8421
rect 19521 8412 19533 8415
rect 19392 8384 19533 8412
rect 19392 8372 19398 8384
rect 19521 8381 19533 8384
rect 19567 8412 19579 8415
rect 19702 8412 19708 8424
rect 19567 8384 19708 8412
rect 19567 8381 19579 8384
rect 19521 8375 19579 8381
rect 19702 8372 19708 8384
rect 19760 8372 19766 8424
rect 20530 8372 20536 8424
rect 20588 8412 20594 8424
rect 20901 8415 20959 8421
rect 20901 8412 20913 8415
rect 20588 8384 20913 8412
rect 20588 8372 20594 8384
rect 20901 8381 20913 8384
rect 20947 8381 20959 8415
rect 20901 8375 20959 8381
rect 20993 8415 21051 8421
rect 20993 8381 21005 8415
rect 21039 8412 21051 8415
rect 21174 8412 21180 8424
rect 21039 8384 21180 8412
rect 21039 8381 21051 8384
rect 20993 8375 21051 8381
rect 21174 8372 21180 8384
rect 21232 8372 21238 8424
rect 21542 8412 21548 8424
rect 21503 8384 21548 8412
rect 21542 8372 21548 8384
rect 21600 8372 21606 8424
rect 21082 8344 21088 8356
rect 19352 8316 21088 8344
rect 19352 8285 19380 8316
rect 21082 8304 21088 8316
rect 21140 8304 21146 8356
rect 18472 8248 19196 8276
rect 19337 8279 19395 8285
rect 18472 8236 18478 8248
rect 19337 8245 19349 8279
rect 19383 8245 19395 8279
rect 19978 8276 19984 8288
rect 19939 8248 19984 8276
rect 19337 8239 19395 8245
rect 19978 8236 19984 8248
rect 20036 8236 20042 8288
rect 20073 8279 20131 8285
rect 20073 8245 20085 8279
rect 20119 8276 20131 8279
rect 20533 8279 20591 8285
rect 20533 8276 20545 8279
rect 20119 8248 20545 8276
rect 20119 8245 20131 8248
rect 20073 8239 20131 8245
rect 20533 8245 20545 8248
rect 20579 8245 20591 8279
rect 20533 8239 20591 8245
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 3050 8072 3056 8084
rect 1627 8044 2912 8072
rect 3011 8044 3056 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 2130 8004 2136 8016
rect 1412 7976 2136 8004
rect 1412 7945 1440 7976
rect 2130 7964 2136 7976
rect 2188 7964 2194 8016
rect 2884 8004 2912 8044
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 3329 8075 3387 8081
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 4709 8075 4767 8081
rect 3375 8044 4660 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 2958 8004 2964 8016
rect 2884 7976 2964 8004
rect 2958 7964 2964 7976
rect 3016 7964 3022 8016
rect 4062 8004 4068 8016
rect 3068 7976 4068 8004
rect 1946 7945 1952 7948
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 1940 7936 1952 7945
rect 1859 7908 1952 7936
rect 1397 7899 1455 7905
rect 1940 7899 1952 7908
rect 2004 7936 2010 7948
rect 3068 7936 3096 7976
rect 4062 7964 4068 7976
rect 4120 8004 4126 8016
rect 4632 8004 4660 8044
rect 4709 8041 4721 8075
rect 4755 8072 4767 8075
rect 5166 8072 5172 8084
rect 4755 8044 5172 8072
rect 4755 8041 4767 8044
rect 4709 8035 4767 8041
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 6822 8032 6828 8084
rect 6880 8032 6886 8084
rect 7098 8072 7104 8084
rect 7059 8044 7104 8072
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 7469 8075 7527 8081
rect 7469 8072 7481 8075
rect 7340 8044 7481 8072
rect 7340 8032 7346 8044
rect 7469 8041 7481 8044
rect 7515 8041 7527 8075
rect 7469 8035 7527 8041
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 8113 8075 8171 8081
rect 7616 8044 7661 8072
rect 7616 8032 7622 8044
rect 8113 8041 8125 8075
rect 8159 8041 8171 8075
rect 8113 8035 8171 8041
rect 8205 8075 8263 8081
rect 8205 8041 8217 8075
rect 8251 8072 8263 8075
rect 8386 8072 8392 8084
rect 8251 8044 8392 8072
rect 8251 8041 8263 8044
rect 8205 8035 8263 8041
rect 4120 7976 4476 8004
rect 4632 7976 5580 8004
rect 4120 7964 4126 7976
rect 3234 7936 3240 7948
rect 2004 7908 3096 7936
rect 3195 7908 3240 7936
rect 1946 7896 1952 7899
rect 2004 7896 2010 7908
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 3510 7936 3516 7948
rect 3471 7908 3516 7936
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 4246 7936 4252 7948
rect 4207 7908 4252 7936
rect 4246 7896 4252 7908
rect 4304 7896 4310 7948
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 1688 7732 1716 7831
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4448 7877 4476 7976
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 5077 7939 5135 7945
rect 5077 7936 5089 7939
rect 4948 7908 5089 7936
rect 4948 7896 4954 7908
rect 5077 7905 5089 7908
rect 5123 7905 5135 7939
rect 5552 7936 5580 7976
rect 5626 7964 5632 8016
rect 5684 8004 5690 8016
rect 6742 8007 6800 8013
rect 6742 8004 6754 8007
rect 5684 7976 6754 8004
rect 5684 7964 5690 7976
rect 6742 7973 6754 7976
rect 6788 7973 6800 8007
rect 6840 8004 6868 8032
rect 6840 7976 7696 8004
rect 6742 7967 6800 7973
rect 7668 7936 7696 7976
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 8128 8004 8156 8035
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8665 8075 8723 8081
rect 8665 8041 8677 8075
rect 8711 8072 8723 8075
rect 8938 8072 8944 8084
rect 8711 8044 8944 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 9950 8072 9956 8084
rect 9140 8044 9956 8072
rect 9140 8004 9168 8044
rect 9950 8032 9956 8044
rect 10008 8072 10014 8084
rect 10778 8072 10784 8084
rect 10008 8044 10784 8072
rect 10008 8032 10014 8044
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 10962 8072 10968 8084
rect 10923 8044 10968 8072
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 12158 8072 12164 8084
rect 11072 8044 12164 8072
rect 7800 7976 9168 8004
rect 7800 7964 7806 7976
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 5552 7908 7420 7936
rect 7668 7908 7941 7936
rect 5077 7899 5135 7905
rect 4341 7871 4399 7877
rect 4341 7868 4353 7871
rect 4212 7840 4353 7868
rect 4212 7828 4218 7840
rect 4341 7837 4353 7840
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 5166 7868 5172 7880
rect 5127 7840 5172 7868
rect 4433 7831 4491 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7055 7840 7328 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 2866 7760 2872 7812
rect 2924 7800 2930 7812
rect 3881 7803 3939 7809
rect 3881 7800 3893 7803
rect 2924 7772 3893 7800
rect 2924 7760 2930 7772
rect 3881 7769 3893 7772
rect 3927 7769 3939 7803
rect 3881 7763 3939 7769
rect 3326 7732 3332 7744
rect 1688 7704 3332 7732
rect 3326 7692 3332 7704
rect 3384 7692 3390 7744
rect 3418 7692 3424 7744
rect 3476 7732 3482 7744
rect 3697 7735 3755 7741
rect 3697 7732 3709 7735
rect 3476 7704 3709 7732
rect 3476 7692 3482 7704
rect 3697 7701 3709 7704
rect 3743 7701 3755 7735
rect 3697 7695 3755 7701
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 5276 7732 5304 7831
rect 4028 7704 5304 7732
rect 5629 7735 5687 7741
rect 4028 7692 4034 7704
rect 5629 7701 5641 7735
rect 5675 7732 5687 7735
rect 6822 7732 6828 7744
rect 5675 7704 6828 7732
rect 5675 7701 5687 7704
rect 5629 7695 5687 7701
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 7300 7732 7328 7840
rect 7392 7800 7420 7908
rect 7929 7905 7941 7908
rect 7975 7905 7987 7939
rect 8570 7936 8576 7948
rect 8531 7908 8576 7936
rect 7929 7899 7987 7905
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 9140 7945 9168 7976
rect 9214 7964 9220 8016
rect 9272 8004 9278 8016
rect 9392 8007 9450 8013
rect 9392 8004 9404 8007
rect 9272 7976 9404 8004
rect 9272 7964 9278 7976
rect 9392 7973 9404 7976
rect 9438 8004 9450 8007
rect 9582 8004 9588 8016
rect 9438 7976 9588 8004
rect 9438 7973 9450 7976
rect 9392 7967 9450 7973
rect 9582 7964 9588 7976
rect 9640 8004 9646 8016
rect 10410 8004 10416 8016
rect 9640 7976 10416 8004
rect 9640 7964 9646 7976
rect 10410 7964 10416 7976
rect 10468 7964 10474 8016
rect 10594 7964 10600 8016
rect 10652 8004 10658 8016
rect 10873 8007 10931 8013
rect 10873 8004 10885 8007
rect 10652 7976 10885 8004
rect 10652 7964 10658 7976
rect 10873 7973 10885 7976
rect 10919 7973 10931 8007
rect 10873 7967 10931 7973
rect 9125 7939 9183 7945
rect 8680 7908 8984 7936
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7524 7840 7665 7868
rect 7524 7828 7530 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 8680 7800 8708 7908
rect 8849 7871 8907 7877
rect 8849 7837 8861 7871
rect 8895 7837 8907 7871
rect 8956 7868 8984 7908
rect 9125 7905 9137 7939
rect 9171 7905 9183 7939
rect 11072 7936 11100 8044
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 12805 8075 12863 8081
rect 12805 8072 12817 8075
rect 12268 8044 12817 8072
rect 12268 8004 12296 8044
rect 12805 8041 12817 8044
rect 12851 8041 12863 8075
rect 12805 8035 12863 8041
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 13412 8044 13461 8072
rect 13412 8032 13418 8044
rect 13449 8041 13461 8044
rect 13495 8041 13507 8075
rect 13449 8035 13507 8041
rect 13722 8032 13728 8084
rect 13780 8072 13786 8084
rect 14369 8075 14427 8081
rect 14369 8072 14381 8075
rect 13780 8044 14381 8072
rect 13780 8032 13786 8044
rect 14369 8041 14381 8044
rect 14415 8041 14427 8075
rect 14369 8035 14427 8041
rect 14829 8075 14887 8081
rect 14829 8041 14841 8075
rect 14875 8072 14887 8075
rect 15562 8072 15568 8084
rect 14875 8044 15568 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 15933 8075 15991 8081
rect 15933 8041 15945 8075
rect 15979 8041 15991 8075
rect 15933 8035 15991 8041
rect 16577 8075 16635 8081
rect 16577 8041 16589 8075
rect 16623 8072 16635 8075
rect 17129 8075 17187 8081
rect 17129 8072 17141 8075
rect 16623 8044 17141 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 17129 8041 17141 8044
rect 17175 8041 17187 8075
rect 17129 8035 17187 8041
rect 17497 8075 17555 8081
rect 17497 8041 17509 8075
rect 17543 8072 17555 8075
rect 19334 8072 19340 8084
rect 17543 8044 19340 8072
rect 17543 8041 17555 8044
rect 17497 8035 17555 8041
rect 9125 7899 9183 7905
rect 9232 7908 11100 7936
rect 11164 7976 12296 8004
rect 12360 7976 12572 8004
rect 9232 7868 9260 7908
rect 8956 7840 9260 7868
rect 8849 7831 8907 7837
rect 7392 7772 8708 7800
rect 7742 7732 7748 7744
rect 7300 7704 7748 7732
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 8864 7732 8892 7831
rect 10410 7828 10416 7880
rect 10468 7868 10474 7880
rect 11164 7868 11192 7976
rect 12089 7939 12147 7945
rect 12089 7905 12101 7939
rect 12135 7936 12147 7939
rect 12250 7936 12256 7948
rect 12135 7908 12256 7936
rect 12135 7905 12147 7908
rect 12089 7899 12147 7905
rect 12250 7896 12256 7908
rect 12308 7896 12314 7948
rect 12360 7945 12388 7976
rect 12345 7939 12403 7945
rect 12345 7905 12357 7939
rect 12391 7905 12403 7939
rect 12544 7936 12572 7976
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 13909 8007 13967 8013
rect 13909 8004 13921 8007
rect 12676 7976 13921 8004
rect 12676 7964 12682 7976
rect 13909 7973 13921 7976
rect 13955 8004 13967 8007
rect 15102 8004 15108 8016
rect 13955 7976 15108 8004
rect 13955 7973 13967 7976
rect 13909 7967 13967 7973
rect 15102 7964 15108 7976
rect 15160 7964 15166 8016
rect 15286 7964 15292 8016
rect 15344 8004 15350 8016
rect 15473 8007 15531 8013
rect 15473 8004 15485 8007
rect 15344 7976 15485 8004
rect 15344 7964 15350 7976
rect 15473 7973 15485 7976
rect 15519 7973 15531 8007
rect 15948 8004 15976 8035
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 19978 8032 19984 8084
rect 20036 8072 20042 8084
rect 20533 8075 20591 8081
rect 20533 8072 20545 8075
rect 20036 8044 20545 8072
rect 20036 8032 20042 8044
rect 20533 8041 20545 8044
rect 20579 8041 20591 8075
rect 21542 8072 21548 8084
rect 21503 8044 21548 8072
rect 20533 8035 20591 8041
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 17586 8004 17592 8016
rect 15948 7976 17592 8004
rect 15473 7967 15531 7973
rect 17586 7964 17592 7976
rect 17644 7964 17650 8016
rect 20901 8007 20959 8013
rect 20901 8004 20913 8007
rect 18156 7976 20913 8004
rect 13170 7936 13176 7948
rect 12544 7908 13176 7936
rect 12345 7899 12403 7905
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 13262 7896 13268 7948
rect 13320 7936 13326 7948
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 13320 7908 13369 7936
rect 13320 7896 13326 7908
rect 13357 7905 13369 7908
rect 13403 7936 13415 7939
rect 13814 7936 13820 7948
rect 13403 7908 13820 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 14734 7936 14740 7948
rect 14647 7908 14740 7936
rect 14734 7896 14740 7908
rect 14792 7936 14798 7948
rect 15565 7939 15623 7945
rect 14792 7908 15516 7936
rect 14792 7896 14798 7908
rect 10468 7840 11192 7868
rect 10468 7828 10474 7840
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12860 7840 12909 7868
rect 12860 7828 12866 7840
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 12434 7760 12440 7812
rect 12492 7800 12498 7812
rect 13004 7800 13032 7831
rect 13078 7828 13084 7880
rect 13136 7868 13142 7880
rect 13722 7868 13728 7880
rect 13136 7840 13728 7868
rect 13136 7828 13142 7840
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 13998 7868 14004 7880
rect 13911 7840 14004 7868
rect 13998 7828 14004 7840
rect 14056 7868 14062 7880
rect 14921 7871 14979 7877
rect 14921 7868 14933 7871
rect 14056 7840 14933 7868
rect 14056 7828 14062 7840
rect 14921 7837 14933 7840
rect 14967 7837 14979 7871
rect 14921 7831 14979 7837
rect 15381 7871 15439 7877
rect 15381 7837 15393 7871
rect 15427 7837 15439 7871
rect 15488 7868 15516 7908
rect 15565 7905 15577 7939
rect 15611 7936 15623 7939
rect 15746 7936 15752 7948
rect 15611 7908 15752 7936
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 15746 7896 15752 7908
rect 15804 7896 15810 7948
rect 16485 7939 16543 7945
rect 16485 7905 16497 7939
rect 16531 7936 16543 7939
rect 16574 7936 16580 7948
rect 16531 7908 16580 7936
rect 16531 7905 16543 7908
rect 16485 7899 16543 7905
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 18156 7936 18184 7976
rect 20548 7948 20576 7976
rect 20901 7973 20913 7976
rect 20947 7973 20959 8007
rect 20901 7967 20959 7973
rect 17604 7908 18184 7936
rect 18224 7939 18282 7945
rect 15654 7868 15660 7880
rect 15488 7840 15660 7868
rect 15381 7831 15439 7837
rect 14016 7800 14044 7828
rect 12492 7772 12537 7800
rect 13004 7772 14044 7800
rect 15396 7800 15424 7831
rect 15654 7828 15660 7840
rect 15712 7828 15718 7880
rect 16022 7868 16028 7880
rect 15983 7840 16028 7868
rect 16022 7828 16028 7840
rect 16080 7828 16086 7880
rect 16393 7871 16451 7877
rect 16393 7837 16405 7871
rect 16439 7868 16451 7871
rect 16758 7868 16764 7880
rect 16439 7840 16764 7868
rect 16439 7837 16451 7840
rect 16393 7831 16451 7837
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 17604 7877 17632 7908
rect 18224 7905 18236 7939
rect 18270 7936 18282 7939
rect 18270 7908 19012 7936
rect 18270 7905 18282 7908
rect 18224 7899 18282 7905
rect 18984 7880 19012 7908
rect 19702 7896 19708 7948
rect 19760 7936 19766 7948
rect 20073 7939 20131 7945
rect 19760 7908 20024 7936
rect 19760 7896 19766 7908
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7837 17647 7871
rect 17589 7831 17647 7837
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7837 17739 7871
rect 17954 7868 17960 7880
rect 17915 7840 17960 7868
rect 17681 7831 17739 7837
rect 15838 7800 15844 7812
rect 15396 7772 15844 7800
rect 12492 7760 12498 7772
rect 9766 7732 9772 7744
rect 8864 7704 9772 7732
rect 9766 7692 9772 7704
rect 9824 7732 9830 7744
rect 10505 7735 10563 7741
rect 10505 7732 10517 7735
rect 9824 7704 10517 7732
rect 9824 7692 9830 7704
rect 10505 7701 10517 7704
rect 10551 7701 10563 7735
rect 10505 7695 10563 7701
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 13004 7732 13032 7772
rect 15838 7760 15844 7772
rect 15896 7800 15902 7812
rect 16945 7803 17003 7809
rect 15896 7772 16896 7800
rect 15896 7760 15902 7772
rect 13078 7732 13084 7744
rect 10652 7704 10697 7732
rect 13004 7704 13084 7732
rect 10652 7692 10658 7704
rect 13078 7692 13084 7704
rect 13136 7692 13142 7744
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 13906 7732 13912 7744
rect 13412 7704 13912 7732
rect 13412 7692 13418 7704
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 16022 7732 16028 7744
rect 15252 7704 16028 7732
rect 15252 7692 15258 7704
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 16390 7692 16396 7744
rect 16448 7732 16454 7744
rect 16758 7732 16764 7744
rect 16448 7704 16764 7732
rect 16448 7692 16454 7704
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 16868 7732 16896 7772
rect 16945 7769 16957 7803
rect 16991 7800 17003 7803
rect 17402 7800 17408 7812
rect 16991 7772 17408 7800
rect 16991 7769 17003 7772
rect 16945 7763 17003 7769
rect 17402 7760 17408 7772
rect 17460 7760 17466 7812
rect 17696 7800 17724 7831
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 18966 7828 18972 7880
rect 19024 7868 19030 7880
rect 19996 7877 20024 7908
rect 20073 7905 20085 7939
rect 20119 7936 20131 7939
rect 20162 7936 20168 7948
rect 20119 7908 20168 7936
rect 20119 7905 20131 7908
rect 20073 7899 20131 7905
rect 20162 7896 20168 7908
rect 20220 7896 20226 7948
rect 20530 7896 20536 7948
rect 20588 7896 20594 7948
rect 21008 7908 21312 7936
rect 19889 7871 19947 7877
rect 19889 7868 19901 7871
rect 19024 7840 19901 7868
rect 19024 7828 19030 7840
rect 19889 7837 19901 7840
rect 19935 7837 19947 7871
rect 19889 7831 19947 7837
rect 19981 7871 20039 7877
rect 19981 7837 19993 7871
rect 20027 7868 20039 7871
rect 20438 7868 20444 7880
rect 20027 7840 20444 7868
rect 20027 7837 20039 7840
rect 19981 7831 20039 7837
rect 17604 7772 17724 7800
rect 19904 7800 19932 7831
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 21008 7877 21036 7908
rect 21284 7880 21312 7908
rect 20993 7871 21051 7877
rect 20993 7868 21005 7871
rect 20864 7840 21005 7868
rect 20864 7828 20870 7840
rect 20993 7837 21005 7840
rect 21039 7837 21051 7871
rect 20993 7831 21051 7837
rect 21085 7871 21143 7877
rect 21085 7837 21097 7871
rect 21131 7837 21143 7871
rect 21085 7831 21143 7837
rect 20714 7800 20720 7812
rect 19904 7772 20720 7800
rect 17604 7732 17632 7772
rect 20714 7760 20720 7772
rect 20772 7800 20778 7812
rect 21100 7800 21128 7831
rect 21266 7828 21272 7880
rect 21324 7828 21330 7880
rect 20772 7772 21128 7800
rect 20772 7760 20778 7772
rect 16868 7704 17632 7732
rect 19337 7735 19395 7741
rect 19337 7701 19349 7735
rect 19383 7732 19395 7735
rect 19886 7732 19892 7744
rect 19383 7704 19892 7732
rect 19383 7701 19395 7704
rect 19337 7695 19395 7701
rect 19886 7692 19892 7704
rect 19944 7692 19950 7744
rect 20438 7732 20444 7744
rect 20399 7704 20444 7732
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 1857 7531 1915 7537
rect 1857 7497 1869 7531
rect 1903 7528 1915 7531
rect 1946 7528 1952 7540
rect 1903 7500 1952 7528
rect 1903 7497 1915 7500
rect 1857 7491 1915 7497
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 3329 7531 3387 7537
rect 3329 7528 3341 7531
rect 2924 7500 3341 7528
rect 2924 7488 2930 7500
rect 3329 7497 3341 7500
rect 3375 7497 3387 7531
rect 3329 7491 3387 7497
rect 3418 7488 3424 7540
rect 3476 7528 3482 7540
rect 3786 7528 3792 7540
rect 3476 7500 3792 7528
rect 3476 7488 3482 7500
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 4154 7528 4160 7540
rect 4115 7500 4160 7528
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4982 7528 4988 7540
rect 4943 7500 4988 7528
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 5074 7488 5080 7540
rect 5132 7528 5138 7540
rect 6457 7531 6515 7537
rect 6457 7528 6469 7531
rect 5132 7500 6469 7528
rect 5132 7488 5138 7500
rect 6457 7497 6469 7500
rect 6503 7497 6515 7531
rect 6457 7491 6515 7497
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 8386 7528 8392 7540
rect 6788 7500 8392 7528
rect 6788 7488 6794 7500
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 8570 7488 8576 7540
rect 8628 7528 8634 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8628 7500 9137 7528
rect 8628 7488 8634 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 10226 7528 10232 7540
rect 9125 7491 9183 7497
rect 9876 7500 10232 7528
rect 6181 7463 6239 7469
rect 6181 7460 6193 7463
rect 3252 7432 6193 7460
rect 3252 7392 3280 7432
rect 6181 7429 6193 7432
rect 6227 7429 6239 7463
rect 9033 7463 9091 7469
rect 6181 7423 6239 7429
rect 6779 7432 7052 7460
rect 3160 7364 3280 7392
rect 3973 7395 4031 7401
rect 1486 7324 1492 7336
rect 1399 7296 1492 7324
rect 1486 7284 1492 7296
rect 1544 7324 1550 7336
rect 3160 7324 3188 7364
rect 3973 7361 3985 7395
rect 4019 7392 4031 7395
rect 4062 7392 4068 7404
rect 4019 7364 4068 7392
rect 4019 7361 4031 7364
rect 3973 7355 4031 7361
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4798 7392 4804 7404
rect 4759 7364 4804 7392
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 5350 7352 5356 7404
rect 5408 7392 5414 7404
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 5408 7364 5549 7392
rect 5408 7352 5414 7364
rect 5537 7361 5549 7364
rect 5583 7392 5595 7395
rect 6779 7392 6807 7432
rect 6914 7392 6920 7404
rect 5583 7364 6807 7392
rect 6875 7364 6920 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7024 7401 7052 7432
rect 9033 7429 9045 7463
rect 9079 7460 9091 7463
rect 9214 7460 9220 7472
rect 9079 7432 9220 7460
rect 9079 7429 9091 7432
rect 9033 7423 9091 7429
rect 9214 7420 9220 7432
rect 9272 7460 9278 7472
rect 9272 7432 9720 7460
rect 9272 7420 9278 7432
rect 7009 7395 7067 7401
rect 7009 7361 7021 7395
rect 7055 7392 7067 7395
rect 7098 7392 7104 7404
rect 7055 7364 7104 7392
rect 7055 7361 7067 7364
rect 7009 7355 7067 7361
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7650 7392 7656 7404
rect 7611 7364 7656 7392
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 9692 7401 9720 7432
rect 9585 7395 9643 7401
rect 9585 7392 9597 7395
rect 9364 7364 9597 7392
rect 9364 7352 9370 7364
rect 1544 7296 3188 7324
rect 3237 7327 3295 7333
rect 1544 7284 1550 7296
rect 3237 7293 3249 7327
rect 3283 7324 3295 7327
rect 3326 7324 3332 7336
rect 3283 7296 3332 7324
rect 3283 7293 3295 7296
rect 3237 7287 3295 7293
rect 3326 7284 3332 7296
rect 3384 7324 3390 7336
rect 4154 7324 4160 7336
rect 3384 7296 4160 7324
rect 3384 7284 3390 7296
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7324 4675 7327
rect 6086 7324 6092 7336
rect 4663 7296 6092 7324
rect 4663 7293 4675 7296
rect 4617 7287 4675 7293
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 2866 7256 2872 7268
rect 1719 7228 2872 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 2866 7216 2872 7228
rect 2924 7216 2930 7268
rect 2981 7259 3039 7265
rect 2981 7225 2993 7259
rect 3027 7225 3039 7259
rect 3789 7259 3847 7265
rect 3789 7256 3801 7259
rect 2981 7219 3039 7225
rect 3344 7228 3801 7256
rect 3007 7188 3035 7219
rect 3344 7200 3372 7228
rect 3789 7225 3801 7228
rect 3835 7225 3847 7259
rect 3789 7219 3847 7225
rect 4062 7216 4068 7268
rect 4120 7256 4126 7268
rect 5813 7259 5871 7265
rect 5813 7256 5825 7259
rect 4120 7228 5825 7256
rect 4120 7216 4126 7228
rect 5813 7225 5825 7228
rect 5859 7225 5871 7259
rect 5813 7219 5871 7225
rect 5902 7216 5908 7268
rect 5960 7256 5966 7268
rect 5960 7228 6960 7256
rect 5960 7216 5966 7228
rect 3234 7188 3240 7200
rect 3007 7160 3240 7188
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 3326 7148 3332 7200
rect 3384 7148 3390 7200
rect 3694 7188 3700 7200
rect 3655 7160 3700 7188
rect 3694 7148 3700 7160
rect 3752 7148 3758 7200
rect 4522 7188 4528 7200
rect 4483 7160 4528 7188
rect 4522 7148 4528 7160
rect 4580 7148 4586 7200
rect 4614 7148 4620 7200
rect 4672 7188 4678 7200
rect 5353 7191 5411 7197
rect 5353 7188 5365 7191
rect 4672 7160 5365 7188
rect 4672 7148 4678 7160
rect 5353 7157 5365 7160
rect 5399 7157 5411 7191
rect 5353 7151 5411 7157
rect 5445 7191 5503 7197
rect 5445 7157 5457 7191
rect 5491 7188 5503 7191
rect 5534 7188 5540 7200
rect 5491 7160 5540 7188
rect 5491 7157 5503 7160
rect 5445 7151 5503 7157
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 5626 7148 5632 7200
rect 5684 7188 5690 7200
rect 5997 7191 6055 7197
rect 5997 7188 6009 7191
rect 5684 7160 6009 7188
rect 5684 7148 5690 7160
rect 5997 7157 6009 7160
rect 6043 7157 6055 7191
rect 5997 7151 6055 7157
rect 6270 7148 6276 7200
rect 6328 7188 6334 7200
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6328 7160 6837 7188
rect 6328 7148 6334 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 6932 7188 6960 7228
rect 7006 7216 7012 7268
rect 7064 7256 7070 7268
rect 7898 7259 7956 7265
rect 7898 7256 7910 7259
rect 7064 7228 7910 7256
rect 7064 7216 7070 7228
rect 7898 7225 7910 7228
rect 7944 7225 7956 7259
rect 9416 7256 9444 7364
rect 9585 7361 9597 7364
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 9493 7327 9551 7333
rect 9493 7293 9505 7327
rect 9539 7324 9551 7327
rect 9876 7324 9904 7500
rect 10226 7488 10232 7500
rect 10284 7528 10290 7540
rect 10873 7531 10931 7537
rect 10873 7528 10885 7531
rect 10284 7500 10885 7528
rect 10284 7488 10290 7500
rect 10873 7497 10885 7500
rect 10919 7528 10931 7531
rect 17957 7531 18015 7537
rect 10919 7500 17908 7528
rect 10919 7497 10931 7500
rect 10873 7491 10931 7497
rect 9950 7420 9956 7472
rect 10008 7460 10014 7472
rect 10045 7463 10103 7469
rect 10045 7460 10057 7463
rect 10008 7432 10057 7460
rect 10008 7420 10014 7432
rect 10045 7429 10057 7432
rect 10091 7460 10103 7463
rect 11238 7460 11244 7472
rect 10091 7432 11244 7460
rect 10091 7429 10103 7432
rect 10045 7423 10103 7429
rect 11238 7420 11244 7432
rect 11296 7420 11302 7472
rect 13265 7463 13323 7469
rect 13265 7429 13277 7463
rect 13311 7460 13323 7463
rect 13354 7460 13360 7472
rect 13311 7432 13360 7460
rect 13311 7429 13323 7432
rect 13265 7423 13323 7429
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 13538 7420 13544 7472
rect 13596 7460 13602 7472
rect 13596 7432 14780 7460
rect 13596 7420 13602 7432
rect 12894 7352 12900 7404
rect 12952 7392 12958 7404
rect 13078 7392 13084 7404
rect 12952 7364 13084 7392
rect 12952 7352 12958 7364
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 13998 7392 14004 7404
rect 13959 7364 14004 7392
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 14752 7401 14780 7432
rect 15102 7420 15108 7472
rect 15160 7460 15166 7472
rect 15289 7463 15347 7469
rect 15289 7460 15301 7463
rect 15160 7432 15301 7460
rect 15160 7420 15166 7432
rect 15289 7429 15301 7432
rect 15335 7460 15347 7463
rect 17770 7460 17776 7472
rect 15335 7432 17776 7460
rect 15335 7429 15347 7432
rect 15289 7423 15347 7429
rect 17770 7420 17776 7432
rect 17828 7420 17834 7472
rect 17880 7460 17908 7500
rect 17957 7497 17969 7531
rect 18003 7528 18015 7531
rect 19058 7528 19064 7540
rect 18003 7500 19064 7528
rect 18003 7497 18015 7500
rect 17957 7491 18015 7497
rect 19058 7488 19064 7500
rect 19116 7488 19122 7540
rect 19242 7488 19248 7540
rect 19300 7528 19306 7540
rect 19337 7531 19395 7537
rect 19337 7528 19349 7531
rect 19300 7500 19349 7528
rect 19300 7488 19306 7500
rect 19337 7497 19349 7500
rect 19383 7497 19395 7531
rect 19337 7491 19395 7497
rect 19426 7488 19432 7540
rect 19484 7528 19490 7540
rect 19613 7531 19671 7537
rect 19613 7528 19625 7531
rect 19484 7500 19625 7528
rect 19484 7488 19490 7500
rect 19613 7497 19625 7500
rect 19659 7497 19671 7531
rect 19613 7491 19671 7497
rect 18506 7460 18512 7472
rect 17880 7432 18512 7460
rect 18506 7420 18512 7432
rect 18564 7420 18570 7472
rect 18785 7463 18843 7469
rect 18785 7429 18797 7463
rect 18831 7460 18843 7463
rect 19978 7460 19984 7472
rect 18831 7432 19984 7460
rect 18831 7429 18843 7432
rect 18785 7423 18843 7429
rect 19978 7420 19984 7432
rect 20036 7420 20042 7472
rect 21818 7460 21824 7472
rect 20088 7432 21824 7460
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 16025 7395 16083 7401
rect 16025 7361 16037 7395
rect 16071 7392 16083 7395
rect 16390 7392 16396 7404
rect 16071 7364 16396 7392
rect 16071 7361 16083 7364
rect 16025 7355 16083 7361
rect 16390 7352 16396 7364
rect 16448 7352 16454 7404
rect 17126 7392 17132 7404
rect 17087 7364 17132 7392
rect 17126 7352 17132 7364
rect 17184 7352 17190 7404
rect 17405 7395 17463 7401
rect 17405 7361 17417 7395
rect 17451 7392 17463 7395
rect 18233 7395 18291 7401
rect 18233 7392 18245 7395
rect 17451 7364 18245 7392
rect 17451 7361 17463 7364
rect 17405 7355 17463 7361
rect 18233 7361 18245 7364
rect 18279 7392 18291 7395
rect 18966 7392 18972 7404
rect 18279 7364 18972 7392
rect 18279 7361 18291 7364
rect 18233 7355 18291 7361
rect 18966 7352 18972 7364
rect 19024 7352 19030 7404
rect 20088 7392 20116 7432
rect 21818 7420 21824 7432
rect 21876 7420 21882 7472
rect 19076 7364 20116 7392
rect 20257 7395 20315 7401
rect 9539 7296 9904 7324
rect 11701 7327 11759 7333
rect 9539 7293 9551 7296
rect 9493 7287 9551 7293
rect 11701 7293 11713 7327
rect 11747 7324 11759 7327
rect 12434 7324 12440 7336
rect 11747 7296 12440 7324
rect 11747 7293 11759 7296
rect 11701 7287 11759 7293
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 13538 7324 13544 7336
rect 12728 7296 13544 7324
rect 10137 7259 10195 7265
rect 10137 7256 10149 7259
rect 9416 7228 10149 7256
rect 7898 7219 7956 7225
rect 10137 7225 10149 7228
rect 10183 7256 10195 7259
rect 10410 7256 10416 7268
rect 10183 7228 10416 7256
rect 10183 7225 10195 7228
rect 10137 7219 10195 7225
rect 10410 7216 10416 7228
rect 10468 7216 10474 7268
rect 10962 7216 10968 7268
rect 11020 7256 11026 7268
rect 11946 7259 12004 7265
rect 11946 7256 11958 7259
rect 11020 7228 11958 7256
rect 11020 7216 11026 7228
rect 11946 7225 11958 7228
rect 11992 7256 12004 7259
rect 12728 7256 12756 7296
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 13906 7324 13912 7336
rect 13771 7296 13912 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 13906 7284 13912 7296
rect 13964 7284 13970 7336
rect 14090 7284 14096 7336
rect 14148 7324 14154 7336
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 14148 7296 14657 7324
rect 14148 7284 14154 7296
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 16666 7324 16672 7336
rect 16627 7296 16672 7324
rect 14645 7287 14703 7293
rect 16666 7284 16672 7296
rect 16724 7324 16730 7336
rect 17497 7327 17555 7333
rect 17497 7324 17509 7327
rect 16724 7296 17509 7324
rect 16724 7284 16730 7296
rect 17497 7293 17509 7296
rect 17543 7293 17555 7327
rect 17497 7287 17555 7293
rect 17586 7284 17592 7336
rect 17644 7324 17650 7336
rect 17644 7296 17689 7324
rect 17644 7284 17650 7296
rect 17770 7284 17776 7336
rect 17828 7324 17834 7336
rect 19076 7324 19104 7364
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20714 7392 20720 7404
rect 20303 7364 20720 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20714 7352 20720 7364
rect 20772 7392 20778 7404
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 20772 7364 21005 7392
rect 20772 7352 20778 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 17828 7296 19104 7324
rect 19153 7327 19211 7333
rect 17828 7284 17834 7296
rect 19153 7293 19165 7327
rect 19199 7324 19211 7327
rect 19242 7324 19248 7336
rect 19199 7296 19248 7324
rect 19199 7293 19211 7296
rect 19153 7287 19211 7293
rect 19242 7284 19248 7296
rect 19300 7324 19306 7336
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 19300 7296 19441 7324
rect 19300 7284 19306 7296
rect 19429 7293 19441 7296
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 19518 7284 19524 7336
rect 19576 7324 19582 7336
rect 19702 7324 19708 7336
rect 19576 7296 19708 7324
rect 19576 7284 19582 7296
rect 19702 7284 19708 7296
rect 19760 7324 19766 7336
rect 20809 7327 20867 7333
rect 20809 7324 20821 7327
rect 19760 7296 20821 7324
rect 19760 7284 19766 7296
rect 20809 7293 20821 7296
rect 20855 7293 20867 7327
rect 21542 7324 21548 7336
rect 21503 7296 21548 7324
rect 20809 7287 20867 7293
rect 21542 7284 21548 7296
rect 21600 7284 21606 7336
rect 13630 7256 13636 7268
rect 11992 7228 12756 7256
rect 12820 7228 13636 7256
rect 11992 7225 12004 7228
rect 11946 7219 12004 7225
rect 7285 7191 7343 7197
rect 7285 7188 7297 7191
rect 6932 7160 7297 7188
rect 6825 7151 6883 7157
rect 7285 7157 7297 7160
rect 7331 7157 7343 7191
rect 7466 7188 7472 7200
rect 7427 7160 7472 7188
rect 7285 7151 7343 7157
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 10318 7188 10324 7200
rect 10279 7160 10324 7188
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 10594 7188 10600 7200
rect 10555 7160 10600 7188
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 11054 7188 11060 7200
rect 11015 7160 11060 7188
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 11422 7188 11428 7200
rect 11204 7160 11249 7188
rect 11383 7160 11428 7188
rect 11204 7148 11210 7160
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 11514 7148 11520 7200
rect 11572 7188 11578 7200
rect 12820 7188 12848 7228
rect 13630 7216 13636 7228
rect 13688 7256 13694 7268
rect 13817 7259 13875 7265
rect 13817 7256 13829 7259
rect 13688 7228 13829 7256
rect 13688 7216 13694 7228
rect 13817 7225 13829 7228
rect 13863 7225 13875 7259
rect 13817 7219 13875 7225
rect 14553 7259 14611 7265
rect 14553 7225 14565 7259
rect 14599 7256 14611 7259
rect 15013 7259 15071 7265
rect 15013 7256 15025 7259
rect 14599 7228 15025 7256
rect 14599 7225 14611 7228
rect 14553 7219 14611 7225
rect 15013 7225 15025 7228
rect 15059 7225 15071 7259
rect 15013 7219 15071 7225
rect 16209 7259 16267 7265
rect 16209 7225 16221 7259
rect 16255 7256 16267 7259
rect 16942 7256 16948 7268
rect 16255 7228 16948 7256
rect 16255 7225 16267 7228
rect 16209 7219 16267 7225
rect 16942 7216 16948 7228
rect 17000 7216 17006 7268
rect 17954 7256 17960 7268
rect 17512 7228 17960 7256
rect 11572 7160 12848 7188
rect 11572 7148 11578 7160
rect 12894 7148 12900 7200
rect 12952 7188 12958 7200
rect 13081 7191 13139 7197
rect 13081 7188 13093 7191
rect 12952 7160 13093 7188
rect 12952 7148 12958 7160
rect 13081 7157 13093 7160
rect 13127 7157 13139 7191
rect 13354 7188 13360 7200
rect 13315 7160 13360 7188
rect 13081 7151 13139 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 14182 7188 14188 7200
rect 14143 7160 14188 7188
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 15286 7188 15292 7200
rect 14424 7160 15292 7188
rect 14424 7148 14430 7160
rect 15286 7148 15292 7160
rect 15344 7188 15350 7200
rect 15473 7191 15531 7197
rect 15473 7188 15485 7191
rect 15344 7160 15485 7188
rect 15344 7148 15350 7160
rect 15473 7157 15485 7160
rect 15519 7157 15531 7191
rect 15654 7188 15660 7200
rect 15615 7160 15660 7188
rect 15473 7151 15531 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 16114 7188 16120 7200
rect 16075 7160 16120 7188
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 16577 7191 16635 7197
rect 16577 7157 16589 7191
rect 16623 7188 16635 7191
rect 17512 7188 17540 7228
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 19058 7256 19064 7268
rect 18064 7228 19064 7256
rect 16623 7160 17540 7188
rect 16623 7157 16635 7160
rect 16577 7151 16635 7157
rect 17678 7148 17684 7200
rect 17736 7188 17742 7200
rect 18064 7188 18092 7228
rect 19058 7216 19064 7228
rect 19116 7256 19122 7268
rect 20073 7259 20131 7265
rect 20073 7256 20085 7259
rect 19116 7228 20085 7256
rect 19116 7216 19122 7228
rect 20073 7225 20085 7228
rect 20119 7225 20131 7259
rect 20073 7219 20131 7225
rect 18322 7188 18328 7200
rect 17736 7160 18092 7188
rect 18283 7160 18328 7188
rect 17736 7148 17742 7160
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 18417 7191 18475 7197
rect 18417 7157 18429 7191
rect 18463 7188 18475 7191
rect 18598 7188 18604 7200
rect 18463 7160 18604 7188
rect 18463 7157 18475 7160
rect 18417 7151 18475 7157
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 18782 7148 18788 7200
rect 18840 7188 18846 7200
rect 18877 7191 18935 7197
rect 18877 7188 18889 7191
rect 18840 7160 18889 7188
rect 18840 7148 18846 7160
rect 18877 7157 18889 7160
rect 18923 7157 18935 7191
rect 18877 7151 18935 7157
rect 19518 7148 19524 7200
rect 19576 7188 19582 7200
rect 19981 7191 20039 7197
rect 19981 7188 19993 7191
rect 19576 7160 19993 7188
rect 19576 7148 19582 7160
rect 19981 7157 19993 7160
rect 20027 7157 20039 7191
rect 19981 7151 20039 7157
rect 20162 7148 20168 7200
rect 20220 7188 20226 7200
rect 20441 7191 20499 7197
rect 20441 7188 20453 7191
rect 20220 7160 20453 7188
rect 20220 7148 20226 7160
rect 20441 7157 20453 7160
rect 20487 7157 20499 7191
rect 20898 7188 20904 7200
rect 20859 7160 20904 7188
rect 20441 7151 20499 7157
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 21361 7191 21419 7197
rect 21361 7157 21373 7191
rect 21407 7188 21419 7191
rect 21450 7188 21456 7200
rect 21407 7160 21456 7188
rect 21407 7157 21419 7160
rect 21361 7151 21419 7157
rect 21450 7148 21456 7160
rect 21508 7148 21514 7200
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 2314 6984 2320 6996
rect 2275 6956 2320 6984
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 2685 6987 2743 6993
rect 2685 6953 2697 6987
rect 2731 6984 2743 6987
rect 3142 6984 3148 6996
rect 2731 6956 3035 6984
rect 3103 6956 3148 6984
rect 2731 6953 2743 6956
rect 2685 6947 2743 6953
rect 1670 6916 1676 6928
rect 1631 6888 1676 6916
rect 1670 6876 1676 6888
rect 1728 6876 1734 6928
rect 3007 6916 3035 6956
rect 3142 6944 3148 6956
rect 3200 6984 3206 6996
rect 4338 6984 4344 6996
rect 3200 6956 4344 6984
rect 3200 6944 3206 6956
rect 4338 6944 4344 6956
rect 4396 6944 4402 6996
rect 4522 6944 4528 6996
rect 4580 6984 4586 6996
rect 6086 6984 6092 6996
rect 4580 6956 5764 6984
rect 6047 6956 6092 6984
rect 4580 6944 4586 6956
rect 3326 6916 3332 6928
rect 3007 6888 3332 6916
rect 3326 6876 3332 6888
rect 3384 6876 3390 6928
rect 3510 6876 3516 6928
rect 3568 6916 3574 6928
rect 3605 6919 3663 6925
rect 3605 6916 3617 6919
rect 3568 6888 3617 6916
rect 3568 6876 3574 6888
rect 3605 6885 3617 6888
rect 3651 6885 3663 6919
rect 3605 6879 3663 6885
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 5736 6916 5764 6956
rect 6086 6944 6092 6956
rect 6144 6944 6150 6996
rect 6457 6987 6515 6993
rect 6457 6953 6469 6987
rect 6503 6984 6515 6987
rect 6730 6984 6736 6996
rect 6503 6956 6736 6984
rect 6503 6953 6515 6956
rect 6457 6947 6515 6953
rect 6730 6944 6736 6956
rect 6788 6944 6794 6996
rect 6917 6987 6975 6993
rect 6917 6953 6929 6987
rect 6963 6953 6975 6987
rect 6917 6947 6975 6953
rect 7285 6987 7343 6993
rect 7285 6953 7297 6987
rect 7331 6984 7343 6987
rect 8202 6984 8208 6996
rect 7331 6956 8208 6984
rect 7331 6953 7343 6956
rect 7285 6947 7343 6953
rect 6932 6916 6960 6947
rect 8202 6944 8208 6956
rect 8260 6984 8266 6996
rect 8260 6956 8708 6984
rect 8260 6944 8266 6956
rect 4212 6888 5304 6916
rect 5736 6888 6960 6916
rect 7377 6919 7435 6925
rect 4212 6876 4218 6888
rect 1486 6848 1492 6860
rect 1447 6820 1492 6848
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 4706 6848 4712 6860
rect 3344 6820 4712 6848
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6749 2191 6783
rect 2133 6743 2191 6749
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2271 6752 2820 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 1394 6604 1400 6656
rect 1452 6644 1458 6656
rect 1765 6647 1823 6653
rect 1765 6644 1777 6647
rect 1452 6616 1777 6644
rect 1452 6604 1458 6616
rect 1765 6613 1777 6616
rect 1811 6613 1823 6647
rect 2148 6644 2176 6743
rect 2792 6721 2820 6752
rect 2958 6740 2964 6792
rect 3016 6780 3022 6792
rect 3234 6780 3240 6792
rect 3016 6752 3240 6780
rect 3016 6740 3022 6752
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3344 6789 3372 6820
rect 4706 6808 4712 6820
rect 4764 6848 4770 6860
rect 5276 6857 5304 6888
rect 7377 6885 7389 6919
rect 7423 6916 7435 6919
rect 8570 6916 8576 6928
rect 7423 6888 8576 6916
rect 7423 6885 7435 6888
rect 7377 6879 7435 6885
rect 8570 6876 8576 6888
rect 8628 6876 8634 6928
rect 8680 6916 8708 6956
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 10318 6984 10324 6996
rect 9272 6956 10180 6984
rect 10279 6956 10324 6984
rect 9272 6944 9278 6956
rect 9677 6919 9735 6925
rect 9677 6916 9689 6919
rect 8680 6888 9689 6916
rect 9677 6885 9689 6888
rect 9723 6885 9735 6919
rect 10152 6916 10180 6956
rect 10318 6944 10324 6956
rect 10376 6944 10382 6996
rect 11241 6987 11299 6993
rect 11241 6953 11253 6987
rect 11287 6984 11299 6987
rect 12250 6984 12256 6996
rect 11287 6956 12256 6984
rect 11287 6953 11299 6956
rect 11241 6947 11299 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 13170 6984 13176 6996
rect 12492 6956 13176 6984
rect 12492 6944 12498 6956
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 13354 6944 13360 6996
rect 13412 6984 13418 6996
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 13412 6956 13737 6984
rect 13412 6944 13418 6956
rect 13725 6953 13737 6956
rect 13771 6953 13783 6987
rect 14090 6984 14096 6996
rect 14051 6956 14096 6984
rect 13725 6947 13783 6953
rect 14090 6944 14096 6956
rect 14148 6984 14154 6996
rect 15841 6987 15899 6993
rect 14148 6956 15608 6984
rect 14148 6944 14154 6956
rect 11146 6916 11152 6928
rect 10152 6888 11152 6916
rect 9677 6879 9735 6885
rect 11146 6876 11152 6888
rect 11204 6876 11210 6928
rect 11333 6919 11391 6925
rect 11333 6885 11345 6919
rect 11379 6916 11391 6919
rect 12342 6916 12348 6928
rect 11379 6888 12348 6916
rect 11379 6885 11391 6888
rect 11333 6879 11391 6885
rect 12342 6876 12348 6888
rect 12400 6876 12406 6928
rect 12986 6876 12992 6928
rect 13044 6916 13050 6928
rect 13044 6888 13124 6916
rect 13044 6876 13050 6888
rect 4994 6851 5052 6857
rect 4994 6848 5006 6851
rect 4764 6820 5006 6848
rect 4764 6808 4770 6820
rect 4994 6817 5006 6820
rect 5040 6817 5052 6851
rect 4994 6811 5052 6817
rect 5261 6851 5319 6857
rect 5261 6817 5273 6851
rect 5307 6817 5319 6851
rect 5261 6811 5319 6817
rect 5534 6808 5540 6860
rect 5592 6857 5598 6860
rect 5592 6848 5603 6857
rect 5813 6851 5871 6857
rect 5592 6820 5637 6848
rect 5592 6811 5603 6820
rect 5813 6817 5825 6851
rect 5859 6848 5871 6851
rect 6086 6848 6092 6860
rect 5859 6820 6092 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 5592 6808 5598 6811
rect 6086 6808 6092 6820
rect 6144 6848 6150 6860
rect 8665 6851 8723 6857
rect 8665 6848 8677 6851
rect 6144 6820 8677 6848
rect 6144 6808 6150 6820
rect 8665 6817 8677 6820
rect 8711 6817 8723 6851
rect 8665 6811 8723 6817
rect 9217 6851 9275 6857
rect 9217 6817 9229 6851
rect 9263 6848 9275 6851
rect 9858 6848 9864 6860
rect 9263 6820 9864 6848
rect 9263 6817 9275 6820
rect 9217 6811 9275 6817
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10873 6851 10931 6857
rect 10376 6820 10548 6848
rect 10376 6808 10382 6820
rect 10520 6792 10548 6820
rect 10873 6817 10885 6851
rect 10919 6848 10931 6851
rect 10962 6848 10968 6860
rect 10919 6820 10968 6848
rect 10919 6817 10931 6820
rect 10873 6811 10931 6817
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 12894 6808 12900 6860
rect 12952 6857 12958 6860
rect 12952 6848 12964 6857
rect 13096 6848 13124 6888
rect 13538 6876 13544 6928
rect 13596 6916 13602 6928
rect 15013 6919 15071 6925
rect 15013 6916 15025 6919
rect 13596 6888 13860 6916
rect 13596 6876 13602 6888
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 12952 6820 12997 6848
rect 13096 6820 13645 6848
rect 12952 6811 12964 6820
rect 13633 6817 13645 6820
rect 13679 6848 13691 6851
rect 13679 6820 13768 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 12952 6808 12958 6811
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6749 3387 6783
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 3329 6743 3387 6749
rect 5276 6752 5917 6780
rect 2777 6715 2835 6721
rect 2777 6681 2789 6715
rect 2823 6681 2835 6715
rect 2777 6675 2835 6681
rect 3142 6672 3148 6724
rect 3200 6712 3206 6724
rect 3344 6712 3372 6743
rect 3200 6684 3372 6712
rect 3200 6672 3206 6684
rect 2222 6644 2228 6656
rect 2135 6616 2228 6644
rect 1765 6607 1823 6613
rect 2222 6604 2228 6616
rect 2280 6644 2286 6656
rect 3050 6644 3056 6656
rect 2280 6616 3056 6644
rect 2280 6604 2286 6616
rect 3050 6604 3056 6616
rect 3108 6644 3114 6656
rect 3786 6644 3792 6656
rect 3108 6616 3792 6644
rect 3108 6604 3114 6616
rect 3786 6604 3792 6616
rect 3844 6644 3850 6656
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3844 6616 3893 6644
rect 3844 6604 3850 6616
rect 3881 6613 3893 6616
rect 3927 6613 3939 6647
rect 3881 6607 3939 6613
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 5276 6644 5304 6752
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 6546 6780 6552 6792
rect 6507 6752 6552 6780
rect 5905 6743 5963 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 7098 6780 7104 6792
rect 6687 6752 7104 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 7098 6740 7104 6752
rect 7156 6780 7162 6792
rect 7469 6783 7527 6789
rect 7469 6780 7481 6783
rect 7156 6752 7481 6780
rect 7156 6740 7162 6752
rect 7469 6749 7481 6752
rect 7515 6749 7527 6783
rect 7469 6743 7527 6749
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 7708 6752 8309 6780
rect 7708 6740 7714 6752
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 9306 6780 9312 6792
rect 8444 6752 9312 6780
rect 8444 6740 8450 6752
rect 9306 6740 9312 6752
rect 9364 6780 9370 6792
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 9364 6752 9505 6780
rect 9364 6740 9370 6752
rect 9493 6749 9505 6752
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9732 6752 9781 6780
rect 9732 6740 9738 6752
rect 9769 6749 9781 6752
rect 9815 6780 9827 6783
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 9815 6752 10425 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 10560 6752 10653 6780
rect 10560 6740 10566 6752
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 13170 6780 13176 6792
rect 11204 6752 11249 6780
rect 13131 6752 13176 6780
rect 11204 6740 11210 6752
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 5359 6721 5365 6724
rect 5353 6675 5365 6721
rect 5417 6712 5423 6724
rect 5417 6684 5453 6712
rect 5359 6672 5365 6675
rect 5417 6672 5423 6684
rect 6730 6672 6736 6724
rect 6788 6712 6794 6724
rect 8113 6715 8171 6721
rect 8113 6712 8125 6715
rect 6788 6684 8125 6712
rect 6788 6672 6794 6684
rect 8113 6681 8125 6684
rect 8159 6681 8171 6715
rect 8478 6712 8484 6724
rect 8439 6684 8484 6712
rect 8113 6675 8171 6681
rect 8478 6672 8484 6684
rect 8536 6672 8542 6724
rect 13188 6712 13216 6740
rect 13740 6712 13768 6820
rect 13832 6789 13860 6888
rect 13924 6888 15025 6916
rect 13817 6783 13875 6789
rect 13817 6749 13829 6783
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 13924 6724 13952 6888
rect 15013 6885 15025 6888
rect 15059 6916 15071 6919
rect 15470 6916 15476 6928
rect 15059 6888 15476 6916
rect 15059 6885 15071 6888
rect 15013 6879 15071 6885
rect 15470 6876 15476 6888
rect 15528 6876 15534 6928
rect 15580 6916 15608 6956
rect 15841 6953 15853 6987
rect 15887 6984 15899 6987
rect 16114 6984 16120 6996
rect 15887 6956 16120 6984
rect 15887 6953 15899 6956
rect 15841 6947 15899 6953
rect 16114 6944 16120 6956
rect 16172 6944 16178 6996
rect 16485 6987 16543 6993
rect 16485 6953 16497 6987
rect 16531 6984 16543 6987
rect 16942 6984 16948 6996
rect 16531 6956 16804 6984
rect 16903 6956 16948 6984
rect 16531 6953 16543 6956
rect 16485 6947 16543 6953
rect 15933 6919 15991 6925
rect 15933 6916 15945 6919
rect 15580 6888 15945 6916
rect 15933 6885 15945 6888
rect 15979 6885 15991 6919
rect 16776 6916 16804 6956
rect 16942 6944 16948 6956
rect 17000 6944 17006 6996
rect 17310 6984 17316 6996
rect 17052 6956 17316 6984
rect 17052 6916 17080 6956
rect 17310 6944 17316 6956
rect 17368 6984 17374 6996
rect 17368 6956 18276 6984
rect 17368 6944 17374 6956
rect 17405 6919 17463 6925
rect 17405 6916 17417 6919
rect 16776 6888 17080 6916
rect 17144 6888 17417 6916
rect 15933 6879 15991 6885
rect 14550 6848 14556 6860
rect 14511 6820 14556 6848
rect 14550 6808 14556 6820
rect 14608 6808 14614 6860
rect 15948 6848 15976 6879
rect 17144 6848 17172 6888
rect 17405 6885 17417 6888
rect 17451 6885 17463 6919
rect 18248 6916 18276 6956
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 18785 6987 18843 6993
rect 18785 6984 18797 6987
rect 18380 6956 18797 6984
rect 18380 6944 18386 6956
rect 18785 6953 18797 6956
rect 18831 6953 18843 6987
rect 20162 6984 20168 6996
rect 20123 6956 20168 6984
rect 18785 6947 18843 6953
rect 20162 6944 20168 6956
rect 20220 6944 20226 6996
rect 20438 6944 20444 6996
rect 20496 6984 20502 6996
rect 20993 6987 21051 6993
rect 20993 6984 21005 6987
rect 20496 6956 21005 6984
rect 20496 6944 20502 6956
rect 20993 6953 21005 6956
rect 21039 6953 21051 6987
rect 21542 6984 21548 6996
rect 21503 6956 21548 6984
rect 20993 6947 21051 6953
rect 21542 6944 21548 6956
rect 21600 6944 21606 6996
rect 20806 6916 20812 6928
rect 18248 6888 20812 6916
rect 17405 6879 17463 6885
rect 20806 6876 20812 6888
rect 20864 6876 20870 6928
rect 20916 6888 21220 6916
rect 17310 6848 17316 6860
rect 15304 6820 15792 6848
rect 15948 6820 17172 6848
rect 17271 6820 17316 6848
rect 15304 6789 15332 6820
rect 15764 6792 15792 6820
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 18325 6851 18383 6857
rect 18325 6848 18337 6851
rect 18104 6820 18337 6848
rect 18104 6808 18110 6820
rect 18325 6817 18337 6820
rect 18371 6817 18383 6851
rect 18325 6811 18383 6817
rect 18414 6808 18420 6860
rect 18472 6848 18478 6860
rect 19061 6851 19119 6857
rect 18472 6820 18517 6848
rect 18472 6808 18478 6820
rect 19061 6817 19073 6851
rect 19107 6848 19119 6851
rect 19242 6848 19248 6860
rect 19107 6820 19248 6848
rect 19107 6817 19119 6820
rect 19061 6811 19119 6817
rect 19242 6808 19248 6820
rect 19300 6848 19306 6860
rect 19337 6851 19395 6857
rect 19337 6848 19349 6851
rect 19300 6820 19349 6848
rect 19300 6808 19306 6820
rect 19337 6817 19349 6820
rect 19383 6817 19395 6851
rect 19337 6811 19395 6817
rect 19978 6808 19984 6860
rect 20036 6848 20042 6860
rect 20073 6851 20131 6857
rect 20073 6848 20085 6851
rect 20036 6820 20085 6848
rect 20036 6808 20042 6820
rect 20073 6817 20085 6820
rect 20119 6817 20131 6851
rect 20916 6848 20944 6888
rect 21082 6848 21088 6860
rect 20073 6811 20131 6817
rect 20180 6820 20944 6848
rect 21043 6820 21088 6848
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 15381 6783 15439 6789
rect 15381 6749 15393 6783
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 13906 6712 13912 6724
rect 9416 6684 12132 6712
rect 13188 6684 13676 6712
rect 13740 6684 13912 6712
rect 9416 6656 9444 6684
rect 4120 6616 5304 6644
rect 4120 6604 4126 6616
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 5629 6647 5687 6653
rect 5629 6644 5641 6647
rect 5592 6616 5641 6644
rect 5592 6604 5598 6616
rect 5629 6613 5641 6616
rect 5675 6644 5687 6647
rect 5810 6644 5816 6656
rect 5675 6616 5816 6644
rect 5675 6613 5687 6616
rect 5629 6607 5687 6613
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 7098 6604 7104 6656
rect 7156 6644 7162 6656
rect 7745 6647 7803 6653
rect 7745 6644 7757 6647
rect 7156 6616 7757 6644
rect 7156 6604 7162 6616
rect 7745 6613 7757 6616
rect 7791 6613 7803 6647
rect 7745 6607 7803 6613
rect 7834 6604 7840 6656
rect 7892 6644 7898 6656
rect 7929 6647 7987 6653
rect 7929 6644 7941 6647
rect 7892 6616 7941 6644
rect 7892 6604 7898 6616
rect 7929 6613 7941 6616
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 8202 6604 8208 6656
rect 8260 6644 8266 6656
rect 8849 6647 8907 6653
rect 8849 6644 8861 6647
rect 8260 6616 8861 6644
rect 8260 6604 8266 6616
rect 8849 6613 8861 6616
rect 8895 6613 8907 6647
rect 9398 6644 9404 6656
rect 9359 6616 9404 6644
rect 8849 6607 8907 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 9950 6644 9956 6656
rect 9732 6616 9777 6644
rect 9911 6616 9956 6644
rect 9732 6604 9738 6616
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10318 6604 10324 6656
rect 10376 6644 10382 6656
rect 10686 6644 10692 6656
rect 10376 6616 10692 6644
rect 10376 6604 10382 6616
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 11698 6644 11704 6656
rect 11659 6616 11704 6644
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 12104 6644 12132 6684
rect 12802 6644 12808 6656
rect 11848 6616 11893 6644
rect 12104 6616 12808 6644
rect 11848 6604 11854 6616
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 13265 6647 13323 6653
rect 13265 6613 13277 6647
rect 13311 6644 13323 6647
rect 13538 6644 13544 6656
rect 13311 6616 13544 6644
rect 13311 6613 13323 6616
rect 13265 6607 13323 6613
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 13648 6644 13676 6684
rect 13906 6672 13912 6684
rect 13964 6672 13970 6724
rect 14734 6672 14740 6724
rect 14792 6712 14798 6724
rect 15396 6712 15424 6743
rect 15746 6740 15752 6792
rect 15804 6740 15810 6792
rect 16114 6740 16120 6792
rect 16172 6780 16178 6792
rect 16577 6783 16635 6789
rect 16577 6780 16589 6783
rect 16172 6752 16589 6780
rect 16172 6740 16178 6752
rect 16577 6749 16589 6752
rect 16623 6749 16635 6783
rect 16577 6743 16635 6749
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 17494 6780 17500 6792
rect 16724 6752 16769 6780
rect 17455 6752 17500 6780
rect 16724 6740 16730 6752
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 17773 6783 17831 6789
rect 17773 6780 17785 6783
rect 17644 6752 17785 6780
rect 17644 6740 17650 6752
rect 17773 6749 17785 6752
rect 17819 6749 17831 6783
rect 18138 6780 18144 6792
rect 18099 6752 18144 6780
rect 17773 6743 17831 6749
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 18966 6740 18972 6792
rect 19024 6780 19030 6792
rect 19153 6783 19211 6789
rect 19153 6780 19165 6783
rect 19024 6752 19165 6780
rect 19024 6740 19030 6752
rect 19153 6749 19165 6752
rect 19199 6749 19211 6783
rect 19886 6780 19892 6792
rect 19799 6752 19892 6780
rect 19153 6743 19211 6749
rect 19886 6740 19892 6752
rect 19944 6780 19950 6792
rect 20180 6780 20208 6820
rect 21082 6808 21088 6820
rect 21140 6808 21146 6860
rect 21192 6789 21220 6888
rect 19944 6752 20208 6780
rect 21177 6783 21235 6789
rect 19944 6740 19950 6752
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 14792 6684 15424 6712
rect 14792 6672 14798 6684
rect 18506 6672 18512 6724
rect 18564 6712 18570 6724
rect 19705 6715 19763 6721
rect 18564 6684 19656 6712
rect 18564 6672 18570 6684
rect 14369 6647 14427 6653
rect 14369 6644 14381 6647
rect 13648 6616 14381 6644
rect 14369 6613 14381 6616
rect 14415 6613 14427 6647
rect 14369 6607 14427 6613
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 14608 6616 14657 6644
rect 14608 6604 14614 6616
rect 14645 6613 14657 6616
rect 14691 6613 14703 6647
rect 14645 6607 14703 6613
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 15562 6644 15568 6656
rect 14884 6616 15568 6644
rect 14884 6604 14890 6616
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 16022 6604 16028 6656
rect 16080 6644 16086 6656
rect 16117 6647 16175 6653
rect 16117 6644 16129 6647
rect 16080 6616 16129 6644
rect 16080 6604 16086 6616
rect 16117 6613 16129 6616
rect 16163 6613 16175 6647
rect 16117 6607 16175 6613
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 17678 6644 17684 6656
rect 16264 6616 17684 6644
rect 16264 6604 16270 6616
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 19628 6644 19656 6684
rect 19705 6681 19717 6715
rect 19751 6712 19763 6715
rect 20438 6712 20444 6724
rect 19751 6684 20444 6712
rect 19751 6681 19763 6684
rect 19705 6675 19763 6681
rect 20438 6672 20444 6684
rect 20496 6672 20502 6724
rect 20533 6715 20591 6721
rect 20533 6681 20545 6715
rect 20579 6712 20591 6715
rect 20990 6712 20996 6724
rect 20579 6684 20996 6712
rect 20579 6681 20591 6684
rect 20533 6675 20591 6681
rect 20990 6672 20996 6684
rect 21048 6672 21054 6724
rect 20162 6644 20168 6656
rect 19628 6616 20168 6644
rect 20162 6604 20168 6616
rect 20220 6604 20226 6656
rect 20254 6604 20260 6656
rect 20312 6644 20318 6656
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 20312 6616 20637 6644
rect 20312 6604 20318 6616
rect 20625 6613 20637 6616
rect 20671 6613 20683 6647
rect 20625 6607 20683 6613
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 1946 6440 1952 6452
rect 1907 6412 1952 6440
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 3694 6440 3700 6452
rect 2823 6412 3700 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 3694 6400 3700 6412
rect 3752 6400 3758 6452
rect 4246 6400 4252 6452
rect 4304 6440 4310 6452
rect 4617 6443 4675 6449
rect 4617 6440 4629 6443
rect 4304 6412 4629 6440
rect 4304 6400 4310 6412
rect 4617 6409 4629 6412
rect 4663 6409 4675 6443
rect 4617 6403 4675 6409
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 5224 6412 5457 6440
rect 5224 6400 5230 6412
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 6730 6440 6736 6452
rect 5776 6412 6736 6440
rect 5776 6400 5782 6412
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 6880 6412 7144 6440
rect 6880 6400 6886 6412
rect 1581 6375 1639 6381
rect 1581 6341 1593 6375
rect 1627 6372 1639 6375
rect 2406 6372 2412 6384
rect 1627 6344 2412 6372
rect 1627 6341 1639 6344
rect 1581 6335 1639 6341
rect 2406 6332 2412 6344
rect 2464 6332 2470 6384
rect 2866 6332 2872 6384
rect 2924 6372 2930 6384
rect 3786 6372 3792 6384
rect 2924 6344 3792 6372
rect 2924 6332 2930 6344
rect 3786 6332 3792 6344
rect 3844 6332 3850 6384
rect 4341 6375 4399 6381
rect 4341 6372 4353 6375
rect 3896 6344 4353 6372
rect 2222 6304 2228 6316
rect 2183 6276 2228 6304
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 3896 6304 3924 6344
rect 4341 6341 4353 6344
rect 4387 6372 4399 6375
rect 4430 6372 4436 6384
rect 4387 6344 4436 6372
rect 4387 6341 4399 6344
rect 4341 6335 4399 6341
rect 4430 6332 4436 6344
rect 4488 6332 4494 6384
rect 4798 6332 4804 6384
rect 4856 6372 4862 6384
rect 4856 6344 5212 6372
rect 4856 6332 4862 6344
rect 2740 6276 3924 6304
rect 3973 6307 4031 6313
rect 2740 6264 2746 6276
rect 3973 6273 3985 6307
rect 4019 6304 4031 6307
rect 4019 6276 4568 6304
rect 4019 6273 4031 6276
rect 3973 6267 4031 6273
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 1762 6236 1768 6248
rect 1723 6208 1768 6236
rect 1397 6199 1455 6205
rect 1210 6128 1216 6180
rect 1268 6168 1274 6180
rect 1412 6168 1440 6199
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 4062 6236 4068 6248
rect 1872 6208 4068 6236
rect 1872 6168 1900 6208
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6236 4215 6239
rect 4246 6236 4252 6248
rect 4203 6208 4252 6236
rect 4203 6205 4215 6208
rect 4157 6199 4215 6205
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 1268 6140 1900 6168
rect 2409 6171 2467 6177
rect 1268 6128 1274 6140
rect 2409 6137 2421 6171
rect 2455 6168 2467 6171
rect 2869 6171 2927 6177
rect 2869 6168 2881 6171
rect 2455 6140 2881 6168
rect 2455 6137 2467 6140
rect 2409 6131 2467 6137
rect 2869 6137 2881 6140
rect 2915 6137 2927 6171
rect 2869 6131 2927 6137
rect 3510 6128 3516 6180
rect 3568 6168 3574 6180
rect 4433 6171 4491 6177
rect 4433 6168 4445 6171
rect 3568 6140 4445 6168
rect 3568 6128 3574 6140
rect 4433 6137 4445 6140
rect 4479 6137 4491 6171
rect 4540 6168 4568 6276
rect 4982 6264 4988 6316
rect 5040 6304 5046 6316
rect 5184 6313 5212 6344
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 5040 6276 5089 6304
rect 5040 6264 5046 6276
rect 5077 6273 5089 6276
rect 5123 6273 5135 6307
rect 5077 6267 5135 6273
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 5997 6307 6055 6313
rect 5997 6304 6009 6307
rect 5592 6276 6009 6304
rect 5592 6264 5598 6276
rect 5997 6273 6009 6276
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 7116 6313 7144 6412
rect 7374 6400 7380 6452
rect 7432 6440 7438 6452
rect 8021 6443 8079 6449
rect 8021 6440 8033 6443
rect 7432 6412 8033 6440
rect 7432 6400 7438 6412
rect 8021 6409 8033 6412
rect 8067 6409 8079 6443
rect 9490 6440 9496 6452
rect 8021 6403 8079 6409
rect 8496 6412 9496 6440
rect 7282 6332 7288 6384
rect 7340 6372 7346 6384
rect 7834 6372 7840 6384
rect 7340 6344 7840 6372
rect 7340 6332 7346 6344
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 6917 6307 6975 6313
rect 6917 6304 6929 6307
rect 6696 6276 6929 6304
rect 6696 6264 6702 6276
rect 6917 6273 6929 6276
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6273 7159 6307
rect 7101 6267 7159 6273
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7248 6276 7389 6304
rect 7248 6264 7254 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7466 6264 7472 6316
rect 7524 6304 7530 6316
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 7524 6276 7573 6304
rect 7524 6264 7530 6276
rect 7561 6273 7573 6276
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 7282 6236 7288 6248
rect 5184 6208 7288 6236
rect 5184 6180 5212 6208
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6236 7711 6239
rect 7742 6236 7748 6248
rect 7699 6208 7748 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 7742 6196 7748 6208
rect 7800 6196 7806 6248
rect 4798 6168 4804 6180
rect 4540 6140 4804 6168
rect 4433 6131 4491 6137
rect 4798 6128 4804 6140
rect 4856 6128 4862 6180
rect 4985 6171 5043 6177
rect 4985 6137 4997 6171
rect 5031 6168 5043 6171
rect 5074 6168 5080 6180
rect 5031 6140 5080 6168
rect 5031 6137 5043 6140
rect 4985 6131 5043 6137
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 5166 6128 5172 6180
rect 5224 6128 5230 6180
rect 8113 6171 8171 6177
rect 8113 6168 8125 6171
rect 6564 6140 8125 6168
rect 6564 6112 6592 6140
rect 8113 6137 8125 6140
rect 8159 6137 8171 6171
rect 8496 6168 8524 6412
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 10321 6443 10379 6449
rect 10321 6409 10333 6443
rect 10367 6440 10379 6443
rect 10367 6412 10824 6440
rect 10367 6409 10379 6412
rect 10321 6403 10379 6409
rect 8662 6332 8668 6384
rect 8720 6372 8726 6384
rect 9674 6372 9680 6384
rect 8720 6344 9680 6372
rect 8720 6332 8726 6344
rect 9674 6332 9680 6344
rect 9732 6332 9738 6384
rect 10796 6372 10824 6412
rect 10962 6400 10968 6452
rect 11020 6440 11026 6452
rect 11020 6412 11192 6440
rect 11020 6400 11026 6412
rect 11054 6372 11060 6384
rect 10796 6344 11060 6372
rect 11054 6332 11060 6344
rect 11112 6332 11118 6384
rect 11164 6372 11192 6412
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 12250 6440 12256 6452
rect 11296 6412 11928 6440
rect 12211 6412 12256 6440
rect 11296 6400 11302 6412
rect 11164 6344 11468 6372
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8628 6276 8953 6304
rect 8628 6264 8634 6276
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 9766 6304 9772 6316
rect 9679 6276 9772 6304
rect 8941 6267 8999 6273
rect 9766 6264 9772 6276
rect 9824 6304 9830 6316
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 9824 6276 10517 6304
rect 9824 6264 9830 6276
rect 10505 6273 10517 6276
rect 10551 6273 10563 6307
rect 11330 6304 11336 6316
rect 10505 6267 10563 6273
rect 10704 6276 11336 6304
rect 9950 6236 9956 6248
rect 8956 6208 9674 6236
rect 9911 6208 9956 6236
rect 8956 6180 8984 6208
rect 8113 6131 8171 6137
rect 8240 6140 8524 6168
rect 8849 6171 8907 6177
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 2498 6100 2504 6112
rect 2363 6072 2504 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 2498 6060 2504 6072
rect 2556 6100 2562 6112
rect 2682 6100 2688 6112
rect 2556 6072 2688 6100
rect 2556 6060 2562 6072
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 3145 6103 3203 6109
rect 3145 6100 3157 6103
rect 3016 6072 3157 6100
rect 3016 6060 3022 6072
rect 3145 6069 3157 6072
rect 3191 6069 3203 6103
rect 3326 6100 3332 6112
rect 3287 6072 3332 6100
rect 3145 6063 3203 6069
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 3694 6100 3700 6112
rect 3655 6072 3700 6100
rect 3694 6060 3700 6072
rect 3752 6060 3758 6112
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 5810 6100 5816 6112
rect 3844 6072 3889 6100
rect 5771 6072 5816 6100
rect 3844 6060 3850 6072
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 5905 6103 5963 6109
rect 5905 6069 5917 6103
rect 5951 6100 5963 6103
rect 6457 6103 6515 6109
rect 6457 6100 6469 6103
rect 5951 6072 6469 6100
rect 5951 6069 5963 6072
rect 5905 6063 5963 6069
rect 6457 6069 6469 6072
rect 6503 6069 6515 6103
rect 6457 6063 6515 6069
rect 6546 6060 6552 6112
rect 6604 6060 6610 6112
rect 6825 6103 6883 6109
rect 6825 6069 6837 6103
rect 6871 6100 6883 6103
rect 8240 6100 8268 6140
rect 8849 6137 8861 6171
rect 8895 6168 8907 6171
rect 8938 6168 8944 6180
rect 8895 6140 8944 6168
rect 8895 6137 8907 6140
rect 8849 6131 8907 6137
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 9306 6168 9312 6180
rect 9267 6140 9312 6168
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 9646 6168 9674 6208
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 10704 6245 10732 6276
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6205 10747 6239
rect 11440 6236 11468 6344
rect 11900 6304 11928 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 12342 6400 12348 6452
rect 12400 6440 12406 6452
rect 13081 6443 13139 6449
rect 13081 6440 13093 6443
rect 12400 6412 13093 6440
rect 12400 6400 12406 6412
rect 13081 6409 13093 6412
rect 13127 6409 13139 6443
rect 13081 6403 13139 6409
rect 13170 6400 13176 6452
rect 13228 6440 13234 6452
rect 21361 6443 21419 6449
rect 21361 6440 21373 6443
rect 13228 6412 21373 6440
rect 13228 6400 13234 6412
rect 21361 6409 21373 6412
rect 21407 6409 21419 6443
rect 22002 6440 22008 6452
rect 21963 6412 22008 6440
rect 21361 6403 21419 6409
rect 22002 6400 22008 6412
rect 22060 6400 22066 6452
rect 12894 6372 12900 6384
rect 12807 6344 12900 6372
rect 12250 6304 12256 6316
rect 11900 6276 12256 6304
rect 12250 6264 12256 6276
rect 12308 6264 12314 6316
rect 12710 6304 12716 6316
rect 12671 6276 12716 6304
rect 12710 6264 12716 6276
rect 12768 6264 12774 6316
rect 12820 6313 12848 6344
rect 12894 6332 12900 6344
rect 12952 6372 12958 6384
rect 13906 6372 13912 6384
rect 12952 6344 13676 6372
rect 13867 6344 13912 6372
rect 12952 6332 12958 6344
rect 12805 6307 12863 6313
rect 12805 6273 12817 6307
rect 12851 6273 12863 6307
rect 13538 6304 13544 6316
rect 13499 6276 13544 6304
rect 12805 6267 12863 6273
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 13648 6313 13676 6344
rect 13906 6332 13912 6344
rect 13964 6332 13970 6384
rect 14090 6332 14096 6384
rect 14148 6372 14154 6384
rect 15013 6375 15071 6381
rect 15013 6372 15025 6375
rect 14148 6344 15025 6372
rect 14148 6332 14154 6344
rect 15013 6341 15025 6344
rect 15059 6341 15071 6375
rect 18509 6375 18567 6381
rect 15013 6335 15071 6341
rect 15856 6344 17540 6372
rect 13633 6307 13691 6313
rect 13633 6273 13645 6307
rect 13679 6273 13691 6307
rect 14274 6304 14280 6316
rect 14235 6276 14280 6304
rect 13633 6267 13691 6273
rect 14274 6264 14280 6276
rect 14332 6264 14338 6316
rect 14461 6307 14519 6313
rect 14461 6273 14473 6307
rect 14507 6304 14519 6307
rect 14826 6304 14832 6316
rect 14507 6276 14832 6304
rect 14507 6273 14519 6276
rect 14461 6267 14519 6273
rect 14826 6264 14832 6276
rect 14884 6264 14890 6316
rect 15746 6264 15752 6316
rect 15804 6304 15810 6316
rect 15856 6313 15884 6344
rect 17512 6316 17540 6344
rect 18509 6341 18521 6375
rect 18555 6372 18567 6375
rect 19150 6372 19156 6384
rect 18555 6344 19156 6372
rect 18555 6341 18567 6344
rect 18509 6335 18567 6341
rect 19150 6332 19156 6344
rect 19208 6332 19214 6384
rect 20625 6375 20683 6381
rect 20625 6341 20637 6375
rect 20671 6372 20683 6375
rect 20714 6372 20720 6384
rect 20671 6344 20720 6372
rect 20671 6341 20683 6344
rect 20625 6335 20683 6341
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 15841 6307 15899 6313
rect 15841 6304 15853 6307
rect 15804 6276 15853 6304
rect 15804 6264 15810 6276
rect 15841 6273 15853 6276
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 16761 6307 16819 6313
rect 16761 6273 16773 6307
rect 16807 6304 16819 6307
rect 17310 6304 17316 6316
rect 16807 6276 17316 6304
rect 16807 6273 16819 6276
rect 16761 6267 16819 6273
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17494 6304 17500 6316
rect 17455 6276 17500 6304
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 17862 6304 17868 6316
rect 17823 6276 17868 6304
rect 17862 6264 17868 6276
rect 17920 6264 17926 6316
rect 18046 6264 18052 6316
rect 18104 6304 18110 6316
rect 18874 6304 18880 6316
rect 18104 6276 18880 6304
rect 18104 6264 18110 6276
rect 18874 6264 18880 6276
rect 18932 6304 18938 6316
rect 19242 6304 19248 6316
rect 18932 6276 19248 6304
rect 18932 6264 18938 6276
rect 19242 6264 19248 6276
rect 19300 6264 19306 6316
rect 11514 6236 11520 6248
rect 11427 6208 11520 6236
rect 10689 6199 10747 6205
rect 11514 6196 11520 6208
rect 11572 6236 11578 6248
rect 13354 6236 13360 6248
rect 11572 6208 13360 6236
rect 11572 6196 11578 6208
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 13449 6239 13507 6245
rect 13449 6205 13461 6239
rect 13495 6236 13507 6239
rect 14182 6236 14188 6248
rect 13495 6208 14188 6236
rect 13495 6205 13507 6208
rect 13449 6199 13507 6205
rect 14182 6196 14188 6208
rect 14240 6196 14246 6248
rect 14550 6236 14556 6248
rect 14511 6208 14556 6236
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 15470 6236 15476 6248
rect 14752 6208 15476 6236
rect 9646 6140 9996 6168
rect 8386 6100 8392 6112
rect 6871 6072 8268 6100
rect 8347 6072 8392 6100
rect 6871 6069 6883 6072
rect 6825 6063 6883 6069
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8757 6103 8815 6109
rect 8757 6069 8769 6103
rect 8803 6100 8815 6103
rect 9122 6100 9128 6112
rect 8803 6072 9128 6100
rect 8803 6069 8815 6072
rect 8757 6063 8815 6069
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9398 6100 9404 6112
rect 9359 6072 9404 6100
rect 9398 6060 9404 6072
rect 9456 6060 9462 6112
rect 9858 6100 9864 6112
rect 9819 6072 9864 6100
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 9968 6100 9996 6140
rect 11238 6128 11244 6180
rect 11296 6168 11302 6180
rect 11333 6171 11391 6177
rect 11333 6168 11345 6171
rect 11296 6140 11345 6168
rect 11296 6128 11302 6140
rect 11333 6137 11345 6140
rect 11379 6168 11391 6171
rect 12618 6168 12624 6180
rect 11379 6140 12204 6168
rect 12579 6140 12624 6168
rect 11379 6137 11391 6140
rect 11333 6131 11391 6137
rect 10594 6100 10600 6112
rect 9968 6072 10600 6100
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 10781 6103 10839 6109
rect 10781 6069 10793 6103
rect 10827 6100 10839 6103
rect 10962 6100 10968 6112
rect 10827 6072 10968 6100
rect 10827 6069 10839 6072
rect 10781 6063 10839 6069
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 11146 6100 11152 6112
rect 11107 6072 11152 6100
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 11422 6100 11428 6112
rect 11383 6072 11428 6100
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 11701 6103 11759 6109
rect 11701 6100 11713 6103
rect 11664 6072 11713 6100
rect 11664 6060 11670 6072
rect 11701 6069 11713 6072
rect 11747 6069 11759 6103
rect 11882 6100 11888 6112
rect 11843 6072 11888 6100
rect 11701 6063 11759 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 12176 6109 12204 6140
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 12802 6128 12808 6180
rect 12860 6168 12866 6180
rect 14752 6168 14780 6208
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 16022 6236 16028 6248
rect 15983 6208 16028 6236
rect 16022 6196 16028 6208
rect 16080 6196 16086 6248
rect 18138 6196 18144 6248
rect 18196 6236 18202 6248
rect 18196 6208 18552 6236
rect 18196 6196 18202 6208
rect 12860 6140 14780 6168
rect 12860 6128 12866 6140
rect 14826 6128 14832 6180
rect 14884 6128 14890 6180
rect 15933 6171 15991 6177
rect 15933 6168 15945 6171
rect 14936 6140 15945 6168
rect 12161 6103 12219 6109
rect 12161 6069 12173 6103
rect 12207 6100 12219 6103
rect 13998 6100 14004 6112
rect 12207 6072 14004 6100
rect 12207 6069 12219 6072
rect 12161 6063 12219 6069
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 14366 6060 14372 6112
rect 14424 6100 14430 6112
rect 14844 6100 14872 6128
rect 14936 6109 14964 6140
rect 15933 6137 15945 6140
rect 15979 6137 15991 6171
rect 15933 6131 15991 6137
rect 17954 6128 17960 6180
rect 18012 6168 18018 6180
rect 18524 6168 18552 6208
rect 19444 6208 21496 6236
rect 19153 6171 19211 6177
rect 18012 6140 18164 6168
rect 18524 6140 19104 6168
rect 18012 6128 18018 6140
rect 14424 6072 14872 6100
rect 14921 6103 14979 6109
rect 14424 6060 14430 6072
rect 14921 6069 14933 6103
rect 14967 6069 14979 6103
rect 14921 6063 14979 6069
rect 15289 6103 15347 6109
rect 15289 6069 15301 6103
rect 15335 6100 15347 6103
rect 15378 6100 15384 6112
rect 15335 6072 15384 6100
rect 15335 6069 15347 6072
rect 15289 6063 15347 6069
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 16393 6103 16451 6109
rect 16393 6069 16405 6103
rect 16439 6100 16451 6103
rect 16758 6100 16764 6112
rect 16439 6072 16764 6100
rect 16439 6069 16451 6072
rect 16393 6063 16451 6069
rect 16758 6060 16764 6072
rect 16816 6060 16822 6112
rect 16942 6100 16948 6112
rect 16903 6072 16948 6100
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 17034 6060 17040 6112
rect 17092 6100 17098 6112
rect 17313 6103 17371 6109
rect 17313 6100 17325 6103
rect 17092 6072 17325 6100
rect 17092 6060 17098 6072
rect 17313 6069 17325 6072
rect 17359 6069 17371 6103
rect 17313 6063 17371 6069
rect 17402 6060 17408 6112
rect 17460 6100 17466 6112
rect 17460 6072 17505 6100
rect 17460 6060 17466 6072
rect 17678 6060 17684 6112
rect 17736 6100 17742 6112
rect 18136 6109 18164 6140
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 17736 6072 18061 6100
rect 17736 6060 17742 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18136 6103 18199 6109
rect 18136 6072 18153 6103
rect 18049 6063 18107 6069
rect 18141 6069 18153 6072
rect 18187 6069 18199 6103
rect 18782 6100 18788 6112
rect 18743 6072 18788 6100
rect 18141 6063 18199 6069
rect 18782 6060 18788 6072
rect 18840 6060 18846 6112
rect 18966 6100 18972 6112
rect 18927 6072 18972 6100
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 19076 6100 19104 6140
rect 19153 6137 19165 6171
rect 19199 6168 19211 6171
rect 19444 6168 19472 6208
rect 19199 6140 19472 6168
rect 19512 6171 19570 6177
rect 19199 6137 19211 6140
rect 19153 6131 19211 6137
rect 19512 6137 19524 6171
rect 19558 6137 19570 6171
rect 19512 6131 19570 6137
rect 19536 6100 19564 6131
rect 20162 6128 20168 6180
rect 20220 6168 20226 6180
rect 20901 6171 20959 6177
rect 20901 6168 20913 6171
rect 20220 6140 20913 6168
rect 20220 6128 20226 6140
rect 20901 6137 20913 6140
rect 20947 6137 20959 6171
rect 21082 6168 21088 6180
rect 21043 6140 21088 6168
rect 20901 6131 20959 6137
rect 21082 6128 21088 6140
rect 21140 6128 21146 6180
rect 21468 6177 21496 6208
rect 21453 6171 21511 6177
rect 21453 6137 21465 6171
rect 21499 6168 21511 6171
rect 21542 6168 21548 6180
rect 21499 6140 21548 6168
rect 21499 6137 21511 6140
rect 21453 6131 21511 6137
rect 21542 6128 21548 6140
rect 21600 6128 21606 6180
rect 19076 6072 19564 6100
rect 19978 6060 19984 6112
rect 20036 6100 20042 6112
rect 20714 6100 20720 6112
rect 20036 6072 20720 6100
rect 20036 6060 20042 6072
rect 20714 6060 20720 6072
rect 20772 6100 20778 6112
rect 21174 6100 21180 6112
rect 20772 6072 21180 6100
rect 20772 6060 20778 6072
rect 21174 6060 21180 6072
rect 21232 6060 21238 6112
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 2866 5896 2872 5908
rect 1627 5868 2872 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3142 5896 3148 5908
rect 3103 5868 3148 5896
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3752 5868 3893 5896
rect 3752 5856 3758 5868
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 3881 5859 3939 5865
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 5442 5896 5448 5908
rect 4028 5868 5448 5896
rect 4028 5856 4034 5868
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5592 5868 5637 5896
rect 5592 5856 5598 5868
rect 5810 5856 5816 5908
rect 5868 5896 5874 5908
rect 6365 5899 6423 5905
rect 6365 5896 6377 5899
rect 5868 5868 6377 5896
rect 5868 5856 5874 5868
rect 6365 5865 6377 5868
rect 6411 5865 6423 5899
rect 6730 5896 6736 5908
rect 6691 5868 6736 5896
rect 6365 5859 6423 5865
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 6825 5899 6883 5905
rect 6825 5865 6837 5899
rect 6871 5896 6883 5899
rect 6871 5868 9352 5896
rect 6871 5865 6883 5868
rect 6825 5859 6883 5865
rect 1946 5788 1952 5840
rect 2004 5837 2010 5840
rect 2004 5831 2068 5837
rect 2004 5797 2022 5831
rect 2056 5797 2068 5831
rect 7469 5831 7527 5837
rect 7469 5828 7481 5831
rect 2004 5791 2068 5797
rect 2746 5800 7481 5828
rect 2004 5788 2010 5791
rect 1302 5720 1308 5772
rect 1360 5760 1366 5772
rect 1397 5763 1455 5769
rect 1397 5760 1409 5763
rect 1360 5732 1409 5760
rect 1360 5720 1366 5732
rect 1397 5729 1409 5732
rect 1443 5760 1455 5763
rect 2746 5760 2774 5800
rect 7469 5797 7481 5800
rect 7515 5797 7527 5831
rect 7469 5791 7527 5797
rect 7926 5788 7932 5840
rect 7984 5828 7990 5840
rect 8113 5831 8171 5837
rect 8113 5828 8125 5831
rect 7984 5800 8125 5828
rect 7984 5788 7990 5800
rect 8113 5797 8125 5800
rect 8159 5828 8171 5831
rect 8573 5831 8631 5837
rect 8159 5800 8340 5828
rect 8159 5797 8171 5800
rect 8113 5791 8171 5797
rect 1443 5732 2774 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 3234 5720 3240 5772
rect 3292 5760 3298 5772
rect 3329 5763 3387 5769
rect 3329 5760 3341 5763
rect 3292 5732 3341 5760
rect 3292 5720 3298 5732
rect 3329 5729 3341 5732
rect 3375 5760 3387 5763
rect 3970 5760 3976 5772
rect 3375 5732 3976 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 4157 5763 4215 5769
rect 4157 5729 4169 5763
rect 4203 5760 4215 5763
rect 4246 5760 4252 5772
rect 4203 5732 4252 5760
rect 4203 5729 4215 5732
rect 4157 5723 4215 5729
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 1780 5556 1808 5655
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3605 5695 3663 5701
rect 3605 5692 3617 5695
rect 3200 5664 3617 5692
rect 3200 5652 3206 5664
rect 3605 5661 3617 5664
rect 3651 5661 3663 5695
rect 3605 5655 3663 5661
rect 4172 5624 4200 5723
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 4424 5763 4482 5769
rect 4424 5729 4436 5763
rect 4470 5760 4482 5763
rect 4798 5760 4804 5772
rect 4470 5732 4804 5760
rect 4470 5729 4482 5732
rect 4424 5723 4482 5729
rect 4798 5720 4804 5732
rect 4856 5760 4862 5772
rect 4856 5732 5488 5760
rect 4856 5720 4862 5732
rect 5460 5692 5488 5732
rect 5718 5720 5724 5772
rect 5776 5760 5782 5772
rect 5813 5763 5871 5769
rect 5813 5760 5825 5763
rect 5776 5732 5825 5760
rect 5776 5720 5782 5732
rect 5813 5729 5825 5732
rect 5859 5729 5871 5763
rect 5813 5723 5871 5729
rect 6089 5763 6147 5769
rect 6089 5729 6101 5763
rect 6135 5760 6147 5763
rect 6178 5760 6184 5772
rect 6135 5732 6184 5760
rect 6135 5729 6147 5732
rect 6089 5723 6147 5729
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 7340 5732 7389 5760
rect 7340 5720 7346 5732
rect 7377 5729 7389 5732
rect 7423 5760 7435 5763
rect 8018 5760 8024 5772
rect 7423 5732 8024 5760
rect 7423 5729 7435 5732
rect 7377 5723 7435 5729
rect 8018 5720 8024 5732
rect 8076 5720 8082 5772
rect 8312 5760 8340 5800
rect 8573 5797 8585 5831
rect 8619 5828 8631 5831
rect 8938 5828 8944 5840
rect 8619 5800 8944 5828
rect 8619 5797 8631 5800
rect 8573 5791 8631 5797
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 9324 5828 9352 5868
rect 9784 5868 10456 5896
rect 9784 5828 9812 5868
rect 10318 5828 10324 5840
rect 9324 5800 9812 5828
rect 9968 5800 10324 5828
rect 9968 5760 9996 5800
rect 10318 5788 10324 5800
rect 10376 5788 10382 5840
rect 10428 5828 10456 5868
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 11701 5899 11759 5905
rect 11701 5896 11713 5899
rect 11020 5868 11713 5896
rect 11020 5856 11026 5868
rect 11701 5865 11713 5868
rect 11747 5865 11759 5899
rect 11701 5859 11759 5865
rect 12161 5899 12219 5905
rect 12161 5865 12173 5899
rect 12207 5896 12219 5899
rect 12342 5896 12348 5908
rect 12207 5868 12348 5896
rect 12207 5865 12219 5868
rect 12161 5859 12219 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12492 5868 14228 5896
rect 12492 5856 12498 5868
rect 11238 5828 11244 5840
rect 10428 5800 11244 5828
rect 11238 5788 11244 5800
rect 11296 5788 11302 5840
rect 11790 5788 11796 5840
rect 11848 5828 11854 5840
rect 12774 5831 12832 5837
rect 12774 5828 12786 5831
rect 11848 5800 12786 5828
rect 11848 5788 11854 5800
rect 12774 5797 12786 5800
rect 12820 5797 12832 5831
rect 12774 5791 12832 5797
rect 12894 5788 12900 5840
rect 12952 5788 12958 5840
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 14093 5831 14151 5837
rect 14093 5828 14105 5831
rect 13872 5800 14105 5828
rect 13872 5788 13878 5800
rect 14093 5797 14105 5800
rect 14139 5797 14151 5831
rect 14093 5791 14151 5797
rect 8312 5732 9996 5760
rect 10502 5720 10508 5772
rect 10560 5769 10566 5772
rect 10560 5760 10572 5769
rect 10560 5732 11468 5760
rect 10560 5723 10572 5732
rect 10560 5720 10566 5723
rect 6822 5692 6828 5704
rect 5460 5664 6828 5692
rect 6822 5652 6828 5664
rect 6880 5692 6886 5704
rect 6917 5695 6975 5701
rect 6917 5692 6929 5695
rect 6880 5664 6929 5692
rect 6880 5652 6886 5664
rect 6917 5661 6929 5664
rect 6963 5661 6975 5695
rect 6917 5655 6975 5661
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 8570 5692 8576 5704
rect 8435 5664 8576 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 7193 5627 7251 5633
rect 7193 5624 7205 5627
rect 2700 5596 4200 5624
rect 5092 5596 7205 5624
rect 2700 5568 2728 5596
rect 2682 5556 2688 5568
rect 1780 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 3513 5559 3571 5565
rect 3513 5525 3525 5559
rect 3559 5556 3571 5559
rect 3694 5556 3700 5568
rect 3559 5528 3700 5556
rect 3559 5525 3571 5528
rect 3513 5519 3571 5525
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 3786 5516 3792 5568
rect 3844 5556 3850 5568
rect 5092 5556 5120 5596
rect 7193 5593 7205 5596
rect 7239 5593 7251 5627
rect 8220 5624 8248 5655
rect 7193 5587 7251 5593
rect 7576 5596 8248 5624
rect 3844 5528 5120 5556
rect 3844 5516 3850 5528
rect 5166 5516 5172 5568
rect 5224 5556 5230 5568
rect 5629 5559 5687 5565
rect 5629 5556 5641 5559
rect 5224 5528 5641 5556
rect 5224 5516 5230 5528
rect 5629 5525 5641 5528
rect 5675 5525 5687 5559
rect 5629 5519 5687 5525
rect 5810 5516 5816 5568
rect 5868 5556 5874 5568
rect 5905 5559 5963 5565
rect 5905 5556 5917 5559
rect 5868 5528 5917 5556
rect 5868 5516 5874 5528
rect 5905 5525 5917 5528
rect 5951 5525 5963 5559
rect 6178 5556 6184 5568
rect 6139 5528 6184 5556
rect 5905 5519 5963 5525
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 7576 5556 7604 5596
rect 6972 5528 7604 5556
rect 6972 5516 6978 5528
rect 7650 5516 7656 5568
rect 7708 5556 7714 5568
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 7708 5528 7757 5556
rect 7708 5516 7714 5528
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 7745 5519 7803 5525
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 8404 5556 8432 5655
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 10778 5692 10784 5704
rect 10739 5664 10784 5692
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 11440 5701 11468 5732
rect 11606 5720 11612 5772
rect 11664 5760 11670 5772
rect 11882 5760 11888 5772
rect 11664 5732 11888 5760
rect 11664 5720 11670 5732
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 12069 5763 12127 5769
rect 12069 5729 12081 5763
rect 12115 5760 12127 5763
rect 12342 5760 12348 5772
rect 12115 5732 12348 5760
rect 12115 5729 12127 5732
rect 12069 5723 12127 5729
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 12529 5763 12587 5769
rect 12529 5729 12541 5763
rect 12575 5760 12587 5763
rect 12912 5760 12940 5788
rect 13262 5760 13268 5772
rect 12575 5732 13268 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 13262 5720 13268 5732
rect 13320 5760 13326 5772
rect 14200 5760 14228 5868
rect 15470 5856 15476 5908
rect 15528 5896 15534 5908
rect 16209 5899 16267 5905
rect 16209 5896 16221 5899
rect 15528 5868 16221 5896
rect 15528 5856 15534 5868
rect 16209 5865 16221 5868
rect 16255 5865 16267 5899
rect 16209 5859 16267 5865
rect 16577 5899 16635 5905
rect 16577 5865 16589 5899
rect 16623 5896 16635 5899
rect 17034 5896 17040 5908
rect 16623 5868 17040 5896
rect 16623 5865 16635 5868
rect 16577 5859 16635 5865
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 17402 5896 17408 5908
rect 17363 5868 17408 5896
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 18049 5899 18107 5905
rect 18049 5865 18061 5899
rect 18095 5896 18107 5899
rect 18138 5896 18144 5908
rect 18095 5868 18144 5896
rect 18095 5865 18107 5868
rect 18049 5859 18107 5865
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 19978 5896 19984 5908
rect 18984 5868 19984 5896
rect 14274 5788 14280 5840
rect 14332 5828 14338 5840
rect 14614 5831 14672 5837
rect 14614 5828 14626 5831
rect 14332 5800 14626 5828
rect 14332 5788 14338 5800
rect 14614 5797 14626 5800
rect 14660 5828 14672 5831
rect 14660 5800 15976 5828
rect 14660 5797 14672 5800
rect 14614 5791 14672 5797
rect 15948 5760 15976 5800
rect 16666 5760 16672 5772
rect 13320 5732 13584 5760
rect 14200 5732 15875 5760
rect 13320 5720 13326 5732
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5661 11391 5695
rect 11333 5655 11391 5661
rect 11425 5695 11483 5701
rect 11425 5661 11437 5695
rect 11471 5692 11483 5695
rect 12253 5695 12311 5701
rect 12253 5692 12265 5695
rect 11471 5664 12265 5692
rect 11471 5661 11483 5664
rect 11425 5655 11483 5661
rect 12253 5661 12265 5664
rect 12299 5661 12311 5695
rect 13556 5692 13584 5732
rect 13998 5692 14004 5704
rect 13556 5664 14004 5692
rect 12253 5655 12311 5661
rect 8662 5584 8668 5636
rect 8720 5624 8726 5636
rect 8849 5627 8907 5633
rect 8849 5624 8861 5627
rect 8720 5596 8861 5624
rect 8720 5584 8726 5596
rect 8849 5593 8861 5596
rect 8895 5593 8907 5627
rect 8849 5587 8907 5593
rect 9401 5627 9459 5633
rect 9401 5593 9413 5627
rect 9447 5624 9459 5627
rect 9766 5624 9772 5636
rect 9447 5596 9772 5624
rect 9447 5593 9459 5596
rect 9401 5587 9459 5593
rect 9766 5584 9772 5596
rect 9824 5584 9830 5636
rect 10873 5627 10931 5633
rect 10873 5593 10885 5627
rect 10919 5624 10931 5627
rect 11238 5624 11244 5636
rect 10919 5596 11244 5624
rect 10919 5593 10931 5596
rect 10873 5587 10931 5593
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 8260 5528 8432 5556
rect 8260 5516 8266 5528
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 9125 5559 9183 5565
rect 9125 5556 9137 5559
rect 8536 5528 9137 5556
rect 8536 5516 8542 5528
rect 9125 5525 9137 5528
rect 9171 5525 9183 5559
rect 9125 5519 9183 5525
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 11348 5556 11376 5655
rect 13998 5652 14004 5664
rect 14056 5692 14062 5704
rect 14369 5695 14427 5701
rect 14369 5692 14381 5695
rect 14056 5664 14381 5692
rect 14056 5652 14062 5664
rect 14369 5661 14381 5664
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 11790 5584 11796 5636
rect 11848 5624 11854 5636
rect 12066 5624 12072 5636
rect 11848 5596 12072 5624
rect 11848 5584 11854 5596
rect 12066 5584 12072 5596
rect 12124 5584 12130 5636
rect 12526 5624 12532 5636
rect 12176 5596 12532 5624
rect 12176 5556 12204 5596
rect 12526 5584 12532 5596
rect 12584 5584 12590 5636
rect 14090 5624 14096 5636
rect 13740 5596 14096 5624
rect 9548 5528 12204 5556
rect 9548 5516 9554 5528
rect 12250 5516 12256 5568
rect 12308 5556 12314 5568
rect 12802 5556 12808 5568
rect 12308 5528 12808 5556
rect 12308 5516 12314 5528
rect 12802 5516 12808 5528
rect 12860 5556 12866 5568
rect 13740 5556 13768 5596
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 15746 5624 15752 5636
rect 15707 5596 15752 5624
rect 15746 5584 15752 5596
rect 15804 5584 15810 5636
rect 15847 5624 15875 5732
rect 15948 5732 16672 5760
rect 15948 5701 15976 5732
rect 16666 5720 16672 5732
rect 16724 5760 16730 5772
rect 16724 5732 16804 5760
rect 16724 5720 16730 5732
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5692 16175 5695
rect 16206 5692 16212 5704
rect 16163 5664 16212 5692
rect 16163 5661 16175 5664
rect 16117 5655 16175 5661
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 16776 5701 16804 5732
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 16945 5763 17003 5769
rect 16945 5760 16957 5763
rect 16908 5732 16957 5760
rect 16908 5720 16914 5732
rect 16945 5729 16957 5732
rect 16991 5729 17003 5763
rect 16945 5723 17003 5729
rect 17037 5763 17095 5769
rect 17037 5729 17049 5763
rect 17083 5760 17095 5763
rect 17218 5760 17224 5772
rect 17083 5732 17224 5760
rect 17083 5729 17095 5732
rect 17037 5723 17095 5729
rect 17218 5720 17224 5732
rect 17276 5760 17282 5772
rect 18984 5760 19012 5868
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 20070 5856 20076 5908
rect 20128 5896 20134 5908
rect 20165 5899 20223 5905
rect 20165 5896 20177 5899
rect 20128 5868 20177 5896
rect 20128 5856 20134 5868
rect 20165 5865 20177 5868
rect 20211 5865 20223 5899
rect 20622 5896 20628 5908
rect 20583 5868 20628 5896
rect 20165 5859 20223 5865
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 19058 5788 19064 5840
rect 19116 5828 19122 5840
rect 20901 5831 20959 5837
rect 20901 5828 20913 5831
rect 19116 5800 20913 5828
rect 19116 5788 19122 5800
rect 20901 5797 20913 5800
rect 20947 5797 20959 5831
rect 20901 5791 20959 5797
rect 21085 5831 21143 5837
rect 21085 5797 21097 5831
rect 21131 5828 21143 5831
rect 22005 5831 22063 5837
rect 22005 5828 22017 5831
rect 21131 5800 22017 5828
rect 21131 5797 21143 5800
rect 21085 5791 21143 5797
rect 22005 5797 22017 5800
rect 22051 5797 22063 5831
rect 22005 5791 22063 5797
rect 19150 5760 19156 5772
rect 19208 5769 19214 5772
rect 17276 5732 19012 5760
rect 19120 5732 19156 5760
rect 17276 5720 17282 5732
rect 19150 5720 19156 5732
rect 19208 5723 19220 5769
rect 20441 5763 20499 5769
rect 19628 5732 20300 5760
rect 19208 5720 19214 5723
rect 16761 5695 16819 5701
rect 16761 5661 16773 5695
rect 16807 5661 16819 5695
rect 19426 5692 19432 5704
rect 19387 5664 19432 5692
rect 16761 5655 16819 5661
rect 19426 5652 19432 5664
rect 19484 5652 19490 5704
rect 17681 5627 17739 5633
rect 17681 5624 17693 5627
rect 15847 5596 17693 5624
rect 17681 5593 17693 5596
rect 17727 5624 17739 5627
rect 17770 5624 17776 5636
rect 17727 5596 17776 5624
rect 17727 5593 17739 5596
rect 17681 5587 17739 5593
rect 17770 5584 17776 5596
rect 17828 5584 17834 5636
rect 17957 5627 18015 5633
rect 17957 5593 17969 5627
rect 18003 5624 18015 5627
rect 18138 5624 18144 5636
rect 18003 5596 18144 5624
rect 18003 5593 18015 5596
rect 17957 5587 18015 5593
rect 18138 5584 18144 5596
rect 18196 5584 18202 5636
rect 13906 5556 13912 5568
rect 12860 5528 13768 5556
rect 13867 5528 13912 5556
rect 12860 5516 12866 5528
rect 13906 5516 13912 5528
rect 13964 5516 13970 5568
rect 14108 5556 14136 5584
rect 19628 5556 19656 5732
rect 19889 5695 19947 5701
rect 19889 5661 19901 5695
rect 19935 5692 19947 5695
rect 19978 5692 19984 5704
rect 19935 5664 19984 5692
rect 19935 5661 19947 5664
rect 19889 5655 19947 5661
rect 19978 5652 19984 5664
rect 20036 5652 20042 5704
rect 19705 5627 19763 5633
rect 19705 5593 19717 5627
rect 19751 5624 19763 5627
rect 20162 5624 20168 5636
rect 19751 5596 20168 5624
rect 19751 5593 19763 5596
rect 19705 5587 19763 5593
rect 20162 5584 20168 5596
rect 20220 5584 20226 5636
rect 20070 5556 20076 5568
rect 14108 5528 19656 5556
rect 20031 5528 20076 5556
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 20272 5556 20300 5732
rect 20441 5729 20453 5763
rect 20487 5729 20499 5763
rect 21450 5760 21456 5772
rect 21411 5732 21456 5760
rect 20441 5723 20499 5729
rect 20464 5636 20492 5723
rect 21450 5720 21456 5732
rect 21508 5720 21514 5772
rect 21269 5695 21327 5701
rect 21269 5692 21281 5695
rect 20548 5664 21281 5692
rect 20438 5584 20444 5636
rect 20496 5584 20502 5636
rect 20548 5556 20576 5664
rect 21269 5661 21281 5664
rect 21315 5661 21327 5695
rect 21269 5655 21327 5661
rect 21284 5596 21588 5624
rect 20272 5528 20576 5556
rect 20809 5559 20867 5565
rect 20809 5525 20821 5559
rect 20855 5556 20867 5559
rect 21284 5556 21312 5596
rect 21560 5568 21588 5596
rect 20855 5528 21312 5556
rect 20855 5525 20867 5528
rect 20809 5519 20867 5525
rect 21542 5516 21548 5568
rect 21600 5516 21606 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 1762 5312 1768 5364
rect 1820 5352 1826 5364
rect 1857 5355 1915 5361
rect 1857 5352 1869 5355
rect 1820 5324 1869 5352
rect 1820 5312 1826 5324
rect 1857 5321 1869 5324
rect 1903 5321 1915 5355
rect 3786 5352 3792 5364
rect 1857 5315 1915 5321
rect 2700 5324 3792 5352
rect 1581 5287 1639 5293
rect 1581 5253 1593 5287
rect 1627 5284 1639 5287
rect 2700 5284 2728 5324
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 4062 5352 4068 5364
rect 4023 5324 4068 5352
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 6733 5355 6791 5361
rect 6733 5352 6745 5355
rect 4632 5324 6745 5352
rect 1627 5256 2728 5284
rect 1627 5253 1639 5256
rect 1581 5247 1639 5253
rect 1946 5176 1952 5228
rect 2004 5216 2010 5228
rect 2409 5219 2467 5225
rect 2409 5216 2421 5219
rect 2004 5188 2421 5216
rect 2004 5176 2010 5188
rect 2409 5185 2421 5188
rect 2455 5185 2467 5219
rect 2682 5216 2688 5228
rect 2643 5188 2688 5216
rect 2409 5179 2467 5185
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 3970 5216 3976 5228
rect 3712 5188 3976 5216
rect 1302 5108 1308 5160
rect 1360 5148 1366 5160
rect 1397 5151 1455 5157
rect 1397 5148 1409 5151
rect 1360 5120 1409 5148
rect 1360 5108 1366 5120
rect 1397 5117 1409 5120
rect 1443 5148 1455 5151
rect 3510 5148 3516 5160
rect 1443 5120 3516 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 3510 5108 3516 5120
rect 3568 5108 3574 5160
rect 2866 5040 2872 5092
rect 2924 5089 2930 5092
rect 2924 5083 2988 5089
rect 2924 5049 2942 5083
rect 2976 5080 2988 5083
rect 3712 5080 3740 5188
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4080 5148 4108 5312
rect 4632 5225 4660 5324
rect 6733 5321 6745 5324
rect 6779 5321 6791 5355
rect 6733 5315 6791 5321
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 8849 5355 8907 5361
rect 8849 5352 8861 5355
rect 6972 5324 8861 5352
rect 6972 5312 6978 5324
rect 8849 5321 8861 5324
rect 8895 5321 8907 5355
rect 10410 5352 10416 5364
rect 8849 5315 8907 5321
rect 9600 5324 10416 5352
rect 9033 5287 9091 5293
rect 9033 5284 9045 5287
rect 6472 5256 9045 5284
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5185 4675 5219
rect 4798 5216 4804 5228
rect 4759 5188 4804 5216
rect 4617 5179 4675 5185
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 4982 5176 4988 5228
rect 5040 5216 5046 5228
rect 5040 5188 5212 5216
rect 5040 5176 5046 5188
rect 2976 5052 3740 5080
rect 3804 5120 4108 5148
rect 2976 5049 2988 5052
rect 2924 5043 2988 5049
rect 2924 5040 2930 5043
rect 2222 5012 2228 5024
rect 2183 4984 2228 5012
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2372 4984 2417 5012
rect 2372 4972 2378 4984
rect 2498 4972 2504 5024
rect 2556 5012 2562 5024
rect 3804 5012 3832 5120
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 4525 5151 4583 5157
rect 4525 5148 4537 5151
rect 4304 5120 4537 5148
rect 4304 5108 4310 5120
rect 4525 5117 4537 5120
rect 4571 5148 4583 5151
rect 5074 5148 5080 5160
rect 4571 5120 5080 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5184 5157 5212 5188
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5316 5188 6009 5216
rect 5316 5176 5322 5188
rect 5997 5185 6009 5188
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 5169 5151 5227 5157
rect 5169 5117 5181 5151
rect 5215 5117 5227 5151
rect 5810 5148 5816 5160
rect 5771 5120 5816 5148
rect 5169 5111 5227 5117
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 6472 5157 6500 5256
rect 9033 5253 9045 5256
rect 9079 5253 9091 5287
rect 9033 5247 9091 5253
rect 7006 5216 7012 5228
rect 6967 5188 7012 5216
rect 7006 5176 7012 5188
rect 7064 5216 7070 5228
rect 7558 5216 7564 5228
rect 7064 5188 7564 5216
rect 7064 5176 7070 5188
rect 7558 5176 7564 5188
rect 7616 5176 7622 5228
rect 7852 5188 8156 5216
rect 6457 5151 6515 5157
rect 6457 5148 6469 5151
rect 5960 5120 6469 5148
rect 5960 5108 5966 5120
rect 6457 5117 6469 5120
rect 6503 5117 6515 5151
rect 6457 5111 6515 5117
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5148 6791 5151
rect 7852 5148 7880 5188
rect 8018 5148 8024 5160
rect 6779 5120 7880 5148
rect 7979 5120 8024 5148
rect 6779 5117 6791 5120
rect 6733 5111 6791 5117
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 8128 5148 8156 5188
rect 8202 5176 8208 5228
rect 8260 5216 8266 5228
rect 9600 5216 9628 5324
rect 10410 5312 10416 5324
rect 10468 5352 10474 5364
rect 10468 5324 14044 5352
rect 10468 5312 10474 5324
rect 13170 5284 13176 5296
rect 12176 5256 13176 5284
rect 8260 5188 8305 5216
rect 8496 5188 9628 5216
rect 10781 5219 10839 5225
rect 8260 5176 8266 5188
rect 8496 5148 8524 5188
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 10965 5219 11023 5225
rect 10965 5185 10977 5219
rect 11011 5216 11023 5219
rect 11146 5216 11152 5228
rect 11011 5188 11152 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 8128 5120 8524 5148
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5148 8631 5151
rect 8662 5148 8668 5160
rect 8619 5120 8668 5148
rect 8619 5117 8631 5120
rect 8573 5111 8631 5117
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 8938 5108 8944 5160
rect 8996 5148 9002 5160
rect 9214 5148 9220 5160
rect 8996 5120 9220 5148
rect 8996 5108 9002 5120
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 10330 5151 10388 5157
rect 10330 5148 10342 5151
rect 9824 5120 10342 5148
rect 9824 5108 9830 5120
rect 10330 5117 10342 5120
rect 10376 5117 10388 5151
rect 10330 5111 10388 5117
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5148 10655 5151
rect 10686 5148 10692 5160
rect 10643 5120 10692 5148
rect 10643 5117 10655 5120
rect 10597 5111 10655 5117
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 3878 5040 3884 5092
rect 3936 5080 3942 5092
rect 6178 5080 6184 5092
rect 3936 5052 6184 5080
rect 3936 5040 3942 5052
rect 6178 5040 6184 5052
rect 6236 5040 6242 5092
rect 7466 5080 7472 5092
rect 6564 5052 7472 5080
rect 2556 4984 3832 5012
rect 2556 4972 2562 4984
rect 3970 4972 3976 5024
rect 4028 5012 4034 5024
rect 4157 5015 4215 5021
rect 4157 5012 4169 5015
rect 4028 4984 4169 5012
rect 4028 4972 4034 4984
rect 4157 4981 4169 4984
rect 4203 4981 4215 5015
rect 4157 4975 4215 4981
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4764 4984 4997 5012
rect 4764 4972 4770 4984
rect 4985 4981 4997 4984
rect 5031 4981 5043 5015
rect 4985 4975 5043 4981
rect 5074 4972 5080 5024
rect 5132 5012 5138 5024
rect 5261 5015 5319 5021
rect 5261 5012 5273 5015
rect 5132 4984 5273 5012
rect 5132 4972 5138 4984
rect 5261 4981 5273 4984
rect 5307 4981 5319 5015
rect 5442 5012 5448 5024
rect 5403 4984 5448 5012
rect 5261 4975 5319 4981
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 5905 5015 5963 5021
rect 5905 4981 5917 5015
rect 5951 5012 5963 5015
rect 6564 5012 6592 5052
rect 7466 5040 7472 5052
rect 7524 5040 7530 5092
rect 9122 5080 9128 5092
rect 7576 5052 9128 5080
rect 5951 4984 6592 5012
rect 6641 5015 6699 5021
rect 5951 4981 5963 4984
rect 5905 4975 5963 4981
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 6730 5012 6736 5024
rect 6687 4984 6736 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 7101 5015 7159 5021
rect 7101 5012 7113 5015
rect 6880 4984 7113 5012
rect 6880 4972 6886 4984
rect 7101 4981 7113 4984
rect 7147 4981 7159 5015
rect 7101 4975 7159 4981
rect 7190 4972 7196 5024
rect 7248 5012 7254 5024
rect 7576 5021 7604 5052
rect 9122 5040 9128 5052
rect 9180 5040 9186 5092
rect 10796 5080 10824 5179
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 12176 5225 12204 5256
rect 13170 5244 13176 5256
rect 13228 5244 13234 5296
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5185 12219 5219
rect 12161 5179 12219 5185
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 12308 5188 12357 5216
rect 12308 5176 12314 5188
rect 12345 5185 12357 5188
rect 12391 5216 12403 5219
rect 12713 5219 12771 5225
rect 12713 5216 12725 5219
rect 12391 5188 12725 5216
rect 12391 5185 12403 5188
rect 12345 5179 12403 5185
rect 12713 5185 12725 5188
rect 12759 5185 12771 5219
rect 12713 5179 12771 5185
rect 11054 5148 11060 5160
rect 11015 5120 11060 5148
rect 11054 5108 11060 5120
rect 11112 5108 11118 5160
rect 11882 5108 11888 5160
rect 11940 5148 11946 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11940 5120 12081 5148
rect 11940 5108 11946 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12728 5148 12756 5179
rect 12802 5176 12808 5228
rect 12860 5216 12866 5228
rect 12860 5188 12905 5216
rect 12860 5176 12866 5188
rect 13078 5176 13084 5228
rect 13136 5216 13142 5228
rect 13538 5216 13544 5228
rect 13136 5188 13544 5216
rect 13136 5176 13142 5188
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 13906 5216 13912 5228
rect 13867 5188 13912 5216
rect 13906 5176 13912 5188
rect 13964 5176 13970 5228
rect 12897 5151 12955 5157
rect 12728 5120 12817 5148
rect 12069 5111 12127 5117
rect 12526 5080 12532 5092
rect 9646 5052 10824 5080
rect 11440 5052 12532 5080
rect 7561 5015 7619 5021
rect 7248 4984 7293 5012
rect 7248 4972 7254 4984
rect 7561 4981 7573 5015
rect 7607 4981 7619 5015
rect 7561 4975 7619 4981
rect 7653 5015 7711 5021
rect 7653 4981 7665 5015
rect 7699 5012 7711 5015
rect 7742 5012 7748 5024
rect 7699 4984 7748 5012
rect 7699 4981 7711 4984
rect 7653 4975 7711 4981
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 8113 5015 8171 5021
rect 8113 4981 8125 5015
rect 8159 5012 8171 5015
rect 8294 5012 8300 5024
rect 8159 4984 8300 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 8665 5015 8723 5021
rect 8665 5012 8677 5015
rect 8628 4984 8677 5012
rect 8628 4972 8634 4984
rect 8665 4981 8677 4984
rect 8711 4981 8723 5015
rect 9214 5012 9220 5024
rect 9175 4984 9220 5012
rect 8665 4975 8723 4981
rect 9214 4972 9220 4984
rect 9272 5012 9278 5024
rect 9646 5012 9674 5052
rect 11440 5021 11468 5052
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 12789 5080 12817 5120
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 13814 5148 13820 5160
rect 12943 5120 13820 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14016 5148 14044 5324
rect 14734 5312 14740 5364
rect 14792 5352 14798 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14792 5324 14933 5352
rect 14792 5312 14798 5324
rect 14921 5321 14933 5324
rect 14967 5321 14979 5355
rect 15654 5352 15660 5364
rect 14921 5315 14979 5321
rect 15028 5324 15660 5352
rect 14274 5216 14280 5228
rect 14235 5188 14280 5216
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 15028 5225 15056 5324
rect 15654 5312 15660 5324
rect 15712 5352 15718 5364
rect 16390 5352 16396 5364
rect 15712 5324 15976 5352
rect 16351 5324 16396 5352
rect 15712 5312 15718 5324
rect 15948 5284 15976 5324
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 17678 5352 17684 5364
rect 17639 5324 17684 5352
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 17957 5355 18015 5361
rect 17957 5321 17969 5355
rect 18003 5352 18015 5355
rect 19242 5352 19248 5364
rect 18003 5324 19248 5352
rect 18003 5321 18015 5324
rect 17957 5315 18015 5321
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19429 5355 19487 5361
rect 19429 5352 19441 5355
rect 19392 5324 19441 5352
rect 19392 5312 19398 5324
rect 19429 5321 19441 5324
rect 19475 5321 19487 5355
rect 19429 5315 19487 5321
rect 15948 5256 18092 5284
rect 18064 5228 18092 5256
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5185 15071 5219
rect 15013 5179 15071 5185
rect 16390 5176 16396 5228
rect 16448 5216 16454 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16448 5188 17049 5216
rect 16448 5176 16454 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 18046 5216 18052 5228
rect 18007 5188 18052 5216
rect 17037 5179 17095 5185
rect 18046 5176 18052 5188
rect 18104 5176 18110 5228
rect 19444 5216 19472 5315
rect 19610 5312 19616 5364
rect 19668 5352 19674 5364
rect 20162 5352 20168 5364
rect 19668 5324 20168 5352
rect 19668 5312 19674 5324
rect 20162 5312 20168 5324
rect 20220 5312 20226 5364
rect 20257 5355 20315 5361
rect 20257 5321 20269 5355
rect 20303 5352 20315 5355
rect 20438 5352 20444 5364
rect 20303 5324 20444 5352
rect 20303 5321 20315 5324
rect 20257 5315 20315 5321
rect 20438 5312 20444 5324
rect 20496 5312 20502 5364
rect 20717 5355 20775 5361
rect 20717 5352 20729 5355
rect 20548 5324 20729 5352
rect 19518 5244 19524 5296
rect 19576 5284 19582 5296
rect 20548 5284 20576 5324
rect 20717 5321 20729 5324
rect 20763 5321 20775 5355
rect 20717 5315 20775 5321
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 21910 5352 21916 5364
rect 20864 5324 21916 5352
rect 20864 5312 20870 5324
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 19576 5256 20576 5284
rect 20625 5287 20683 5293
rect 19576 5244 19582 5256
rect 20625 5253 20637 5287
rect 20671 5284 20683 5287
rect 22278 5284 22284 5296
rect 20671 5256 22284 5284
rect 20671 5253 20683 5256
rect 20625 5247 20683 5253
rect 22278 5244 22284 5256
rect 22336 5244 22342 5296
rect 19613 5219 19671 5225
rect 19613 5216 19625 5219
rect 19444 5188 19625 5216
rect 19613 5185 19625 5188
rect 19659 5185 19671 5219
rect 21266 5216 21272 5228
rect 19613 5179 19671 5185
rect 19720 5188 20944 5216
rect 21227 5188 21272 5216
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 14016 5120 14565 5148
rect 14553 5117 14565 5120
rect 14599 5117 14611 5151
rect 14553 5111 14611 5117
rect 15280 5151 15338 5157
rect 15280 5117 15292 5151
rect 15326 5148 15338 5151
rect 15746 5148 15752 5160
rect 15326 5120 15752 5148
rect 15326 5117 15338 5120
rect 15280 5111 15338 5117
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 16942 5108 16948 5160
rect 17000 5148 17006 5160
rect 17313 5151 17371 5157
rect 17313 5148 17325 5151
rect 17000 5120 17325 5148
rect 17000 5108 17006 5120
rect 17313 5117 17325 5120
rect 17359 5117 17371 5151
rect 17313 5111 17371 5117
rect 18782 5108 18788 5160
rect 18840 5148 18846 5160
rect 19720 5148 19748 5188
rect 18840 5120 19748 5148
rect 20441 5151 20499 5157
rect 18840 5108 18846 5120
rect 20441 5117 20453 5151
rect 20487 5148 20499 5151
rect 20806 5148 20812 5160
rect 20487 5120 20812 5148
rect 20487 5117 20499 5120
rect 20441 5111 20499 5117
rect 20806 5108 20812 5120
rect 20864 5108 20870 5160
rect 20916 5157 20944 5188
rect 21266 5176 21272 5188
rect 21324 5176 21330 5228
rect 20901 5151 20959 5157
rect 20901 5117 20913 5151
rect 20947 5148 20959 5151
rect 21082 5148 21088 5160
rect 20947 5120 21088 5148
rect 20947 5117 20959 5120
rect 20901 5111 20959 5117
rect 21082 5108 21088 5120
rect 21140 5108 21146 5160
rect 21177 5151 21235 5157
rect 21177 5117 21189 5151
rect 21223 5148 21235 5151
rect 21726 5148 21732 5160
rect 21223 5120 21732 5148
rect 21223 5117 21235 5120
rect 21177 5111 21235 5117
rect 21726 5108 21732 5120
rect 21784 5108 21790 5160
rect 13906 5080 13912 5092
rect 12789 5052 13912 5080
rect 13906 5040 13912 5052
rect 13964 5040 13970 5092
rect 14734 5040 14740 5092
rect 14792 5080 14798 5092
rect 16669 5083 16727 5089
rect 16669 5080 16681 5083
rect 14792 5052 16681 5080
rect 14792 5040 14798 5052
rect 16669 5049 16681 5052
rect 16715 5049 16727 5083
rect 16669 5043 16727 5049
rect 16758 5040 16764 5092
rect 16816 5080 16822 5092
rect 17221 5083 17279 5089
rect 17221 5080 17233 5083
rect 16816 5052 17233 5080
rect 16816 5040 16822 5052
rect 17221 5049 17233 5052
rect 17267 5049 17279 5083
rect 17221 5043 17279 5049
rect 18230 5040 18236 5092
rect 18288 5089 18294 5092
rect 18288 5083 18352 5089
rect 18288 5049 18306 5083
rect 18340 5049 18352 5083
rect 18288 5043 18352 5049
rect 18288 5040 18294 5043
rect 18414 5040 18420 5092
rect 18472 5080 18478 5092
rect 19889 5083 19947 5089
rect 19889 5080 19901 5083
rect 18472 5052 19901 5080
rect 18472 5040 18478 5052
rect 19889 5049 19901 5052
rect 19935 5049 19947 5083
rect 19889 5043 19947 5049
rect 20070 5040 20076 5092
rect 20128 5080 20134 5092
rect 21450 5080 21456 5092
rect 20128 5052 21456 5080
rect 20128 5040 20134 5052
rect 21450 5040 21456 5052
rect 21508 5040 21514 5092
rect 9272 4984 9674 5012
rect 11425 5015 11483 5021
rect 9272 4972 9278 4984
rect 11425 4981 11437 5015
rect 11471 4981 11483 5015
rect 11425 4975 11483 4981
rect 11606 4972 11612 5024
rect 11664 5012 11670 5024
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11664 4984 11713 5012
rect 11664 4972 11670 4984
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 11701 4975 11759 4981
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 12342 5012 12348 5024
rect 11940 4984 12348 5012
rect 11940 4972 11946 4984
rect 12342 4972 12348 4984
rect 12400 4972 12406 5024
rect 13262 5012 13268 5024
rect 13223 4984 13268 5012
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 13354 4972 13360 5024
rect 13412 5012 13418 5024
rect 13412 4984 13457 5012
rect 13412 4972 13418 4984
rect 13538 4972 13544 5024
rect 13596 5012 13602 5024
rect 13725 5015 13783 5021
rect 13725 5012 13737 5015
rect 13596 4984 13737 5012
rect 13596 4972 13602 4984
rect 13725 4981 13737 4984
rect 13771 4981 13783 5015
rect 13725 4975 13783 4981
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 14090 5012 14096 5024
rect 13872 4984 14096 5012
rect 13872 4972 13878 4984
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14366 4972 14372 5024
rect 14424 5012 14430 5024
rect 14461 5015 14519 5021
rect 14461 5012 14473 5015
rect 14424 4984 14473 5012
rect 14424 4972 14430 4984
rect 14461 4981 14473 4984
rect 14507 5012 14519 5015
rect 16577 5015 16635 5021
rect 16577 5012 16589 5015
rect 14507 4984 16589 5012
rect 14507 4981 14519 4984
rect 14461 4975 14519 4981
rect 16577 4981 16589 4984
rect 16623 5012 16635 5015
rect 17034 5012 17040 5024
rect 16623 4984 17040 5012
rect 16623 4981 16635 4984
rect 16577 4975 16635 4981
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 17310 4972 17316 5024
rect 17368 5012 17374 5024
rect 18138 5012 18144 5024
rect 17368 4984 18144 5012
rect 17368 4972 17374 4984
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 19797 5015 19855 5021
rect 19797 5012 19809 5015
rect 18840 4984 19809 5012
rect 18840 4972 18846 4984
rect 19797 4981 19809 4984
rect 19843 4981 19855 5015
rect 19797 4975 19855 4981
rect 20162 4972 20168 5024
rect 20220 5012 20226 5024
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20220 4984 21005 5012
rect 20220 4972 20226 4984
rect 20993 4981 21005 4984
rect 21039 4981 21051 5015
rect 20993 4975 21051 4981
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 1397 4811 1455 4817
rect 1397 4777 1409 4811
rect 1443 4808 1455 4811
rect 1946 4808 1952 4820
rect 1443 4780 1952 4808
rect 1443 4777 1455 4780
rect 1397 4771 1455 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2314 4768 2320 4820
rect 2372 4808 2378 4820
rect 2961 4811 3019 4817
rect 2961 4808 2973 4811
rect 2372 4780 2973 4808
rect 2372 4768 2378 4780
rect 2961 4777 2973 4780
rect 3007 4777 3019 4811
rect 2961 4771 3019 4777
rect 3329 4811 3387 4817
rect 3329 4777 3341 4811
rect 3375 4808 3387 4811
rect 3881 4811 3939 4817
rect 3881 4808 3893 4811
rect 3375 4780 3893 4808
rect 3375 4777 3387 4780
rect 3329 4771 3387 4777
rect 3881 4777 3893 4780
rect 3927 4777 3939 4811
rect 3881 4771 3939 4777
rect 4341 4811 4399 4817
rect 4341 4777 4353 4811
rect 4387 4808 4399 4811
rect 4709 4811 4767 4817
rect 4709 4808 4721 4811
rect 4387 4780 4721 4808
rect 4387 4777 4399 4780
rect 4341 4771 4399 4777
rect 4709 4777 4721 4780
rect 4755 4777 4767 4811
rect 4709 4771 4767 4777
rect 5169 4811 5227 4817
rect 5169 4777 5181 4811
rect 5215 4808 5227 4811
rect 6270 4808 6276 4820
rect 5215 4780 6276 4808
rect 5215 4777 5227 4780
rect 5169 4771 5227 4777
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 7282 4808 7288 4820
rect 7243 4780 7288 4808
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 7742 4808 7748 4820
rect 7703 4780 7748 4808
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 9674 4808 9680 4820
rect 8619 4780 9680 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 9916 4780 10241 4808
rect 9916 4768 9922 4780
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 10229 4771 10287 4777
rect 10689 4811 10747 4817
rect 10689 4777 10701 4811
rect 10735 4808 10747 4811
rect 11149 4811 11207 4817
rect 11149 4808 11161 4811
rect 10735 4780 11161 4808
rect 10735 4777 10747 4780
rect 10689 4771 10747 4777
rect 11149 4777 11161 4780
rect 11195 4777 11207 4811
rect 11149 4771 11207 4777
rect 12253 4811 12311 4817
rect 12253 4777 12265 4811
rect 12299 4808 12311 4811
rect 13078 4808 13084 4820
rect 12299 4780 13084 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 13170 4768 13176 4820
rect 13228 4808 13234 4820
rect 14921 4811 14979 4817
rect 14921 4808 14933 4811
rect 13228 4780 14933 4808
rect 13228 4768 13234 4780
rect 14921 4777 14933 4780
rect 14967 4777 14979 4811
rect 14921 4771 14979 4777
rect 16945 4811 17003 4817
rect 16945 4777 16957 4811
rect 16991 4808 17003 4811
rect 17218 4808 17224 4820
rect 16991 4780 17224 4808
rect 16991 4777 17003 4780
rect 16945 4771 17003 4777
rect 17218 4768 17224 4780
rect 17276 4808 17282 4820
rect 17862 4808 17868 4820
rect 17276 4780 17868 4808
rect 17276 4768 17282 4780
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 17957 4811 18015 4817
rect 17957 4777 17969 4811
rect 18003 4808 18015 4811
rect 18414 4808 18420 4820
rect 18003 4780 18420 4808
rect 18003 4777 18015 4780
rect 17957 4771 18015 4777
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 18782 4808 18788 4820
rect 18743 4780 18788 4808
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 18874 4768 18880 4820
rect 18932 4808 18938 4820
rect 19058 4808 19064 4820
rect 18932 4780 19064 4808
rect 18932 4768 18938 4780
rect 19058 4768 19064 4780
rect 19116 4768 19122 4820
rect 19613 4811 19671 4817
rect 19613 4777 19625 4811
rect 19659 4777 19671 4811
rect 19613 4771 19671 4777
rect 3050 4700 3056 4752
rect 3108 4740 3114 4752
rect 4249 4743 4307 4749
rect 3108 4712 4200 4740
rect 3108 4700 3114 4712
rect 2521 4675 2579 4681
rect 2521 4641 2533 4675
rect 2567 4672 2579 4675
rect 2682 4672 2688 4684
rect 2567 4644 2688 4672
rect 2567 4641 2579 4644
rect 2521 4635 2579 4641
rect 2682 4632 2688 4644
rect 2740 4672 2746 4684
rect 4172 4672 4200 4712
rect 4249 4709 4261 4743
rect 4295 4740 4307 4743
rect 5626 4740 5632 4752
rect 4295 4712 5632 4740
rect 4295 4709 4307 4712
rect 4249 4703 4307 4709
rect 5626 4700 5632 4712
rect 5684 4700 5690 4752
rect 6764 4743 6822 4749
rect 6764 4709 6776 4743
rect 6810 4740 6822 4743
rect 6810 4712 7604 4740
rect 6810 4709 6822 4712
rect 6764 4703 6822 4709
rect 4706 4672 4712 4684
rect 2740 4644 3556 4672
rect 4172 4644 4712 4672
rect 2740 4632 2746 4644
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4573 2835 4607
rect 3418 4604 3424 4616
rect 3379 4576 3424 4604
rect 2777 4567 2835 4573
rect 2590 4428 2596 4480
rect 2648 4468 2654 4480
rect 2792 4468 2820 4567
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 3528 4613 3556 4644
rect 4706 4632 4712 4644
rect 4764 4632 4770 4684
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 5810 4672 5816 4684
rect 5123 4644 5816 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 7098 4672 7104 4684
rect 7011 4644 7104 4672
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7576 4672 7604 4712
rect 7650 4700 7656 4752
rect 7708 4740 7714 4752
rect 7837 4743 7895 4749
rect 7837 4740 7849 4743
rect 7708 4712 7849 4740
rect 7708 4700 7714 4712
rect 7837 4709 7849 4712
rect 7883 4709 7895 4743
rect 9214 4740 9220 4752
rect 7837 4703 7895 4709
rect 8956 4712 9220 4740
rect 8956 4672 8984 4712
rect 9214 4700 9220 4712
rect 9272 4700 9278 4752
rect 10502 4740 10508 4752
rect 9646 4712 10508 4740
rect 9122 4672 9128 4684
rect 7576 4644 8984 4672
rect 9083 4644 9128 4672
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 9646 4672 9674 4712
rect 10502 4700 10508 4712
rect 10560 4700 10566 4752
rect 10597 4743 10655 4749
rect 10597 4709 10609 4743
rect 10643 4740 10655 4743
rect 11606 4740 11612 4752
rect 10643 4712 11612 4740
rect 10643 4709 10655 4712
rect 10597 4703 10655 4709
rect 11606 4700 11612 4712
rect 11664 4700 11670 4752
rect 11977 4743 12035 4749
rect 11977 4709 11989 4743
rect 12023 4740 12035 4743
rect 14369 4743 14427 4749
rect 14369 4740 14381 4743
rect 12023 4712 12296 4740
rect 12023 4709 12035 4712
rect 11977 4703 12035 4709
rect 12268 4684 12296 4712
rect 12544 4712 14381 4740
rect 9600 4644 9674 4672
rect 9861 4675 9919 4681
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 4338 4564 4344 4616
rect 4396 4604 4402 4616
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4396 4576 4445 4604
rect 4396 4564 4402 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 7009 4607 7067 4613
rect 5316 4576 5672 4604
rect 5316 4564 5322 4576
rect 3050 4496 3056 4548
rect 3108 4536 3114 4548
rect 4982 4536 4988 4548
rect 3108 4508 4988 4536
rect 3108 4496 3114 4508
rect 4982 4496 4988 4508
rect 5040 4496 5046 4548
rect 5644 4545 5672 4576
rect 7009 4573 7021 4607
rect 7055 4573 7067 4607
rect 7116 4604 7144 4632
rect 7282 4604 7288 4616
rect 7116 4576 7288 4604
rect 7009 4567 7067 4573
rect 5629 4539 5687 4545
rect 5629 4505 5641 4539
rect 5675 4505 5687 4539
rect 5629 4499 5687 4505
rect 3786 4468 3792 4480
rect 2648 4440 3792 4468
rect 2648 4428 2654 4440
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 4246 4428 4252 4480
rect 4304 4468 4310 4480
rect 5718 4468 5724 4480
rect 4304 4440 5724 4468
rect 4304 4428 4310 4440
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 6730 4428 6736 4480
rect 6788 4468 6794 4480
rect 7024 4468 7052 4567
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 7374 4564 7380 4616
rect 7432 4564 7438 4616
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4604 8079 4607
rect 8202 4604 8208 4616
rect 8067 4576 8208 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8481 4607 8539 4613
rect 8352 4576 8397 4604
rect 8352 4564 8358 4576
rect 8481 4573 8493 4607
rect 8527 4604 8539 4607
rect 9490 4604 9496 4616
rect 8527 4576 9496 4604
rect 8527 4573 8539 4576
rect 8481 4567 8539 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 9600 4613 9628 4644
rect 9861 4641 9873 4675
rect 9907 4641 9919 4675
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 9861 4635 9919 4641
rect 10980 4644 11529 4672
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4573 9643 4607
rect 9766 4604 9772 4616
rect 9727 4576 9772 4604
rect 9585 4567 9643 4573
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 7392 4536 7420 4564
rect 9876 4536 9904 4635
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 7392 4508 9904 4536
rect 10520 4536 10548 4567
rect 10778 4564 10784 4616
rect 10836 4604 10842 4616
rect 10980 4604 11008 4644
rect 11517 4641 11529 4644
rect 11563 4641 11575 4675
rect 11882 4672 11888 4684
rect 11517 4635 11575 4641
rect 11624 4644 11888 4672
rect 11054 4604 11060 4616
rect 10836 4576 11060 4604
rect 10836 4564 10842 4576
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 11238 4564 11244 4616
rect 11296 4604 11302 4616
rect 11624 4613 11652 4644
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 12066 4672 12072 4684
rect 12027 4644 12072 4672
rect 12066 4632 12072 4644
rect 12124 4632 12130 4684
rect 12250 4632 12256 4684
rect 12308 4632 12314 4684
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 12544 4681 12572 4712
rect 14369 4709 14381 4712
rect 14415 4709 14427 4743
rect 15832 4743 15890 4749
rect 14369 4703 14427 4709
rect 15396 4712 15792 4740
rect 12529 4675 12587 4681
rect 12529 4672 12541 4675
rect 12492 4644 12541 4672
rect 12492 4632 12498 4644
rect 12529 4641 12541 4644
rect 12575 4641 12587 4675
rect 12529 4635 12587 4641
rect 13814 4632 13820 4684
rect 13872 4681 13878 4684
rect 13872 4672 13884 4681
rect 13872 4644 13917 4672
rect 13872 4635 13884 4644
rect 13872 4632 13878 4635
rect 13998 4632 14004 4684
rect 14056 4672 14062 4684
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 14056 4644 14105 4672
rect 14056 4632 14062 4644
rect 14093 4641 14105 4644
rect 14139 4641 14151 4675
rect 14093 4635 14151 4641
rect 14550 4632 14556 4684
rect 14608 4672 14614 4684
rect 15197 4675 15255 4681
rect 15197 4672 15209 4675
rect 14608 4644 15209 4672
rect 14608 4632 14614 4644
rect 15197 4641 15209 4644
rect 15243 4641 15255 4675
rect 15197 4635 15255 4641
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 11296 4576 11621 4604
rect 11296 4564 11302 4576
rect 11609 4573 11621 4576
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 12158 4604 12164 4616
rect 11839 4576 12164 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 14366 4564 14372 4616
rect 14424 4604 14430 4616
rect 14645 4607 14703 4613
rect 14645 4604 14657 4607
rect 14424 4576 14657 4604
rect 14424 4564 14430 4576
rect 14645 4573 14657 4576
rect 14691 4604 14703 4607
rect 15396 4604 15424 4712
rect 15565 4675 15623 4681
rect 15565 4641 15577 4675
rect 15611 4672 15623 4675
rect 15654 4672 15660 4684
rect 15611 4644 15660 4672
rect 15611 4641 15623 4644
rect 15565 4635 15623 4641
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 15764 4672 15792 4712
rect 15832 4709 15844 4743
rect 15878 4740 15890 4743
rect 16390 4740 16396 4752
rect 15878 4712 16396 4740
rect 15878 4709 15890 4712
rect 15832 4703 15890 4709
rect 16390 4700 16396 4712
rect 16448 4700 16454 4752
rect 17589 4743 17647 4749
rect 17589 4709 17601 4743
rect 17635 4740 17647 4743
rect 19628 4740 19656 4771
rect 19978 4768 19984 4820
rect 20036 4808 20042 4820
rect 20073 4811 20131 4817
rect 20073 4808 20085 4811
rect 20036 4780 20085 4808
rect 20036 4768 20042 4780
rect 20073 4777 20085 4780
rect 20119 4777 20131 4811
rect 20073 4771 20131 4777
rect 20254 4768 20260 4820
rect 20312 4808 20318 4820
rect 20441 4811 20499 4817
rect 20441 4808 20453 4811
rect 20312 4780 20453 4808
rect 20312 4768 20318 4780
rect 20441 4777 20453 4780
rect 20487 4777 20499 4811
rect 20714 4808 20720 4820
rect 20675 4780 20720 4808
rect 20441 4771 20499 4777
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 21361 4811 21419 4817
rect 21361 4777 21373 4811
rect 21407 4808 21419 4811
rect 21818 4808 21824 4820
rect 21407 4780 21824 4808
rect 21407 4777 21419 4780
rect 21361 4771 21419 4777
rect 21818 4768 21824 4780
rect 21876 4768 21882 4820
rect 17635 4712 19656 4740
rect 19812 4712 21220 4740
rect 17635 4709 17647 4712
rect 17589 4703 17647 4709
rect 17310 4672 17316 4684
rect 15764 4644 17316 4672
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 17678 4672 17684 4684
rect 17420 4644 17684 4672
rect 17420 4613 17448 4644
rect 17678 4632 17684 4644
rect 17736 4672 17742 4684
rect 18417 4675 18475 4681
rect 17736 4644 18276 4672
rect 17736 4632 17742 4644
rect 18248 4616 18276 4644
rect 18417 4641 18429 4675
rect 18463 4672 18475 4675
rect 18782 4672 18788 4684
rect 18463 4644 18788 4672
rect 18463 4641 18475 4644
rect 18417 4635 18475 4641
rect 18782 4632 18788 4644
rect 18840 4632 18846 4684
rect 19150 4672 19156 4684
rect 19111 4644 19156 4672
rect 19150 4632 19156 4644
rect 19208 4632 19214 4684
rect 19242 4632 19248 4684
rect 19300 4672 19306 4684
rect 19812 4672 19840 4712
rect 19978 4672 19984 4684
rect 19300 4644 19840 4672
rect 19939 4644 19984 4672
rect 19300 4632 19306 4644
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 20625 4675 20683 4681
rect 20625 4641 20637 4675
rect 20671 4641 20683 4675
rect 20898 4672 20904 4684
rect 20859 4644 20904 4672
rect 20625 4635 20683 4641
rect 14691 4576 15424 4604
rect 17405 4607 17463 4613
rect 14691 4573 14703 4576
rect 14645 4567 14703 4573
rect 17405 4573 17417 4607
rect 17451 4573 17463 4607
rect 17405 4567 17463 4573
rect 17497 4607 17555 4613
rect 17497 4573 17509 4607
rect 17543 4604 17555 4607
rect 18046 4604 18052 4616
rect 17543 4576 18052 4604
rect 17543 4573 17555 4576
rect 17497 4567 17555 4573
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 18230 4604 18236 4616
rect 18191 4576 18236 4604
rect 18230 4564 18236 4576
rect 18288 4564 18294 4616
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4604 18383 4607
rect 19610 4604 19616 4616
rect 18371 4576 19616 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 19610 4564 19616 4576
rect 19668 4564 19674 4616
rect 20165 4607 20223 4613
rect 20165 4573 20177 4607
rect 20211 4573 20223 4607
rect 20165 4567 20223 4573
rect 12618 4536 12624 4548
rect 10520 4508 12624 4536
rect 12618 4496 12624 4508
rect 12676 4536 12682 4548
rect 12713 4539 12771 4545
rect 12713 4536 12725 4539
rect 12676 4508 12725 4536
rect 12676 4496 12682 4508
rect 12713 4505 12725 4508
rect 12759 4505 12771 4539
rect 18874 4536 18880 4548
rect 12713 4499 12771 4505
rect 17052 4508 18880 4536
rect 7374 4468 7380 4480
rect 6788 4440 7052 4468
rect 7335 4440 7380 4468
rect 6788 4428 6794 4440
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 8754 4428 8760 4480
rect 8812 4468 8818 4480
rect 8941 4471 8999 4477
rect 8941 4468 8953 4471
rect 8812 4440 8953 4468
rect 8812 4428 8818 4440
rect 8941 4437 8953 4440
rect 8987 4437 8999 4471
rect 9306 4468 9312 4480
rect 9267 4440 9312 4468
rect 8941 4431 8999 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 11057 4471 11115 4477
rect 11057 4437 11069 4471
rect 11103 4468 11115 4471
rect 11977 4471 12035 4477
rect 11977 4468 11989 4471
rect 11103 4440 11989 4468
rect 11103 4437 11115 4440
rect 11057 4431 11115 4437
rect 11977 4437 11989 4440
rect 12023 4437 12035 4471
rect 12342 4468 12348 4480
rect 12303 4440 12348 4468
rect 11977 4431 12035 4437
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 14737 4471 14795 4477
rect 14737 4468 14749 4471
rect 14240 4440 14749 4468
rect 14240 4428 14246 4440
rect 14737 4437 14749 4440
rect 14783 4468 14795 4471
rect 15286 4468 15292 4480
rect 14783 4440 15292 4468
rect 14783 4437 14795 4440
rect 14737 4431 14795 4437
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 15381 4471 15439 4477
rect 15381 4437 15393 4471
rect 15427 4468 15439 4471
rect 17052 4468 17080 4508
rect 18874 4496 18880 4508
rect 18932 4496 18938 4548
rect 18984 4508 19288 4536
rect 15427 4440 17080 4468
rect 17129 4471 17187 4477
rect 15427 4437 15439 4440
rect 15381 4431 15439 4437
rect 17129 4437 17141 4471
rect 17175 4468 17187 4471
rect 18984 4468 19012 4508
rect 17175 4440 19012 4468
rect 19061 4471 19119 4477
rect 17175 4437 17187 4440
rect 17129 4431 17187 4437
rect 19061 4437 19073 4471
rect 19107 4468 19119 4471
rect 19150 4468 19156 4480
rect 19107 4440 19156 4468
rect 19107 4437 19119 4440
rect 19061 4431 19119 4437
rect 19150 4428 19156 4440
rect 19208 4428 19214 4480
rect 19260 4468 19288 4508
rect 19794 4496 19800 4548
rect 19852 4536 19858 4548
rect 20180 4536 20208 4567
rect 19852 4508 20208 4536
rect 19852 4496 19858 4508
rect 19334 4468 19340 4480
rect 19260 4440 19340 4468
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 19429 4471 19487 4477
rect 19429 4437 19441 4471
rect 19475 4468 19487 4471
rect 20070 4468 20076 4480
rect 19475 4440 20076 4468
rect 19475 4437 19487 4440
rect 19429 4431 19487 4437
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 20162 4428 20168 4480
rect 20220 4468 20226 4480
rect 20640 4468 20668 4635
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 21192 4681 21220 4712
rect 21177 4675 21235 4681
rect 21177 4641 21189 4675
rect 21223 4641 21235 4675
rect 21450 4672 21456 4684
rect 21411 4644 21456 4672
rect 21177 4635 21235 4641
rect 21192 4604 21220 4635
rect 21450 4632 21456 4644
rect 21508 4632 21514 4684
rect 21818 4604 21824 4616
rect 21192 4576 21824 4604
rect 21818 4564 21824 4576
rect 21876 4564 21882 4616
rect 20990 4468 20996 4480
rect 20220 4440 20668 4468
rect 20951 4440 20996 4468
rect 20220 4428 20226 4440
rect 20990 4428 20996 4440
rect 21048 4428 21054 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 2682 4264 2688 4276
rect 2643 4236 2688 4264
rect 2682 4224 2688 4236
rect 2740 4224 2746 4276
rect 6273 4267 6331 4273
rect 6273 4233 6285 4267
rect 6319 4264 6331 4267
rect 7190 4264 7196 4276
rect 6319 4236 7196 4264
rect 6319 4233 6331 4236
rect 6273 4227 6331 4233
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 7558 4224 7564 4276
rect 7616 4264 7622 4276
rect 8205 4267 8263 4273
rect 8205 4264 8217 4267
rect 7616 4236 8217 4264
rect 7616 4224 7622 4236
rect 8205 4233 8217 4236
rect 8251 4233 8263 4267
rect 8205 4227 8263 4233
rect 8846 4224 8852 4276
rect 8904 4264 8910 4276
rect 8904 4236 8984 4264
rect 8904 4224 8910 4236
rect 2866 4196 2872 4208
rect 1964 4168 2872 4196
rect 1964 4137 1992 4168
rect 2866 4156 2872 4168
rect 2924 4156 2930 4208
rect 4706 4196 4712 4208
rect 4080 4168 4712 4196
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 2958 4128 2964 4140
rect 1949 4091 2007 4097
rect 2056 4100 2964 4128
rect 1302 4020 1308 4072
rect 1360 4060 1366 4072
rect 1397 4063 1455 4069
rect 1397 4060 1409 4063
rect 1360 4032 1409 4060
rect 1360 4020 1366 4032
rect 1397 4029 1409 4032
rect 1443 4060 1455 4063
rect 2056 4060 2084 4100
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 4080 4137 4108 4168
rect 4706 4156 4712 4168
rect 4764 4196 4770 4208
rect 6730 4196 6736 4208
rect 4764 4168 6736 4196
rect 4764 4156 4770 4168
rect 6730 4156 6736 4168
rect 6788 4196 6794 4208
rect 8297 4199 8355 4205
rect 6788 4168 6868 4196
rect 6788 4156 6794 4168
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4097 4123 4131
rect 5074 4128 5080 4140
rect 4065 4091 4123 4097
rect 4356 4100 5080 4128
rect 1443 4032 2084 4060
rect 2133 4063 2191 4069
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 2133 4029 2145 4063
rect 2179 4060 2191 4063
rect 3970 4060 3976 4072
rect 2179 4032 3976 4060
rect 2179 4029 2191 4032
rect 2133 4023 2191 4029
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 4356 4069 4384 4100
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5258 4128 5264 4140
rect 5219 4100 5264 4128
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 5994 4128 6000 4140
rect 5767 4100 6000 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 6840 4137 6868 4168
rect 8297 4165 8309 4199
rect 8343 4165 8355 4199
rect 8297 4159 8355 4165
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 4430 4020 4436 4072
rect 4488 4020 4494 4072
rect 4614 4060 4620 4072
rect 4575 4032 4620 4060
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 6641 4063 6699 4069
rect 6641 4060 6653 4063
rect 5736 4032 6653 4060
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 3326 3992 3332 4004
rect 2271 3964 3332 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 3326 3952 3332 3964
rect 3384 3952 3390 4004
rect 3602 3952 3608 4004
rect 3660 3992 3666 4004
rect 3820 3995 3878 4001
rect 3820 3992 3832 3995
rect 3660 3964 3832 3992
rect 3660 3952 3666 3964
rect 3820 3961 3832 3964
rect 3866 3992 3878 3995
rect 4448 3992 4476 4020
rect 5736 4004 5764 4032
rect 6641 4029 6653 4032
rect 6687 4029 6699 4063
rect 7374 4060 7380 4072
rect 6641 4023 6699 4029
rect 6748 4032 7380 4060
rect 3866 3964 4384 3992
rect 4448 3964 4752 3992
rect 3866 3961 3878 3964
rect 3820 3955 3878 3961
rect 4356 3936 4384 3964
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 1854 3924 1860 3936
rect 1811 3896 1860 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 2593 3927 2651 3933
rect 2593 3893 2605 3927
rect 2639 3924 2651 3927
rect 3970 3924 3976 3936
rect 2639 3896 3976 3924
rect 2639 3893 2651 3896
rect 2593 3887 2651 3893
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 4154 3924 4160 3936
rect 4115 3896 4160 3924
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4338 3884 4344 3936
rect 4396 3884 4402 3936
rect 4430 3884 4436 3936
rect 4488 3924 4494 3936
rect 4724 3933 4752 3964
rect 5718 3952 5724 4004
rect 5776 3952 5782 4004
rect 5905 3995 5963 4001
rect 5905 3961 5917 3995
rect 5951 3992 5963 3995
rect 6748 3992 6776 4032
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 7466 4020 7472 4072
rect 7524 4060 7530 4072
rect 8312 4060 8340 4159
rect 8754 4128 8760 4140
rect 8715 4100 8760 4128
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4097 8907 4131
rect 8956 4128 8984 4236
rect 9306 4224 9312 4276
rect 9364 4264 9370 4276
rect 14366 4264 14372 4276
rect 9364 4236 14372 4264
rect 9364 4224 9370 4236
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 15286 4224 15292 4276
rect 15344 4264 15350 4276
rect 15746 4264 15752 4276
rect 15344 4236 15752 4264
rect 15344 4224 15350 4236
rect 15746 4224 15752 4236
rect 15804 4224 15810 4276
rect 17678 4264 17684 4276
rect 17639 4236 17684 4264
rect 17678 4224 17684 4236
rect 17736 4224 17742 4276
rect 18046 4224 18052 4276
rect 18104 4264 18110 4276
rect 19153 4267 19211 4273
rect 19153 4264 19165 4267
rect 18104 4236 19165 4264
rect 18104 4224 18110 4236
rect 19153 4233 19165 4236
rect 19199 4233 19211 4267
rect 19153 4227 19211 4233
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 20898 4264 20904 4276
rect 19392 4236 20904 4264
rect 19392 4224 19398 4236
rect 20898 4224 20904 4236
rect 20956 4264 20962 4276
rect 21450 4264 21456 4276
rect 20956 4236 21456 4264
rect 20956 4224 20962 4236
rect 21450 4224 21456 4236
rect 21508 4224 21514 4276
rect 9490 4196 9496 4208
rect 9451 4168 9496 4196
rect 9490 4156 9496 4168
rect 9548 4156 9554 4208
rect 9858 4156 9864 4208
rect 9916 4196 9922 4208
rect 9916 4168 12296 4196
rect 9916 4156 9922 4168
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 8956 4100 9137 4128
rect 8849 4091 8907 4097
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 7524 4032 8340 4060
rect 7524 4020 7530 4032
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8444 4032 8677 4060
rect 8444 4020 8450 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 8665 4023 8723 4029
rect 7070 3995 7128 4001
rect 7070 3992 7082 3995
rect 5951 3964 6776 3992
rect 6840 3964 7082 3992
rect 5951 3961 5963 3964
rect 5905 3955 5963 3961
rect 4709 3927 4767 3933
rect 4488 3896 4533 3924
rect 4488 3884 4494 3896
rect 4709 3893 4721 3927
rect 4755 3893 4767 3927
rect 4709 3887 4767 3893
rect 4982 3884 4988 3936
rect 5040 3924 5046 3936
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 5040 3896 5089 3924
rect 5040 3884 5046 3896
rect 5077 3893 5089 3896
rect 5123 3893 5135 3927
rect 5077 3887 5135 3893
rect 5169 3927 5227 3933
rect 5169 3893 5181 3927
rect 5215 3924 5227 3927
rect 5350 3924 5356 3936
rect 5215 3896 5356 3924
rect 5215 3893 5227 3896
rect 5169 3887 5227 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 5810 3924 5816 3936
rect 5771 3896 5816 3924
rect 5810 3884 5816 3896
rect 5868 3884 5874 3936
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 6638 3924 6644 3936
rect 6503 3896 6644 3924
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 6840 3924 6868 3964
rect 7070 3961 7082 3964
rect 7116 3961 7128 3995
rect 7070 3955 7128 3961
rect 8202 3952 8208 4004
rect 8260 3992 8266 4004
rect 8864 3992 8892 4091
rect 9674 4088 9680 4140
rect 9732 4128 9738 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9732 4100 10057 4128
rect 9732 4088 9738 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10870 4088 10876 4140
rect 10928 4128 10934 4140
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 10928 4100 11069 4128
rect 10928 4088 10934 4100
rect 11057 4097 11069 4100
rect 11103 4097 11115 4131
rect 12158 4128 12164 4140
rect 12119 4100 12164 4128
rect 11057 4091 11115 4097
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12268 4137 12296 4168
rect 12526 4156 12532 4208
rect 12584 4196 12590 4208
rect 16942 4196 16948 4208
rect 12584 4168 16948 4196
rect 12584 4156 12590 4168
rect 16942 4156 16948 4168
rect 17000 4156 17006 4208
rect 20441 4199 20499 4205
rect 20441 4165 20453 4199
rect 20487 4196 20499 4199
rect 20530 4196 20536 4208
rect 20487 4168 20536 4196
rect 20487 4165 20499 4168
rect 20441 4159 20499 4165
rect 20530 4156 20536 4168
rect 20588 4156 20594 4208
rect 20806 4196 20812 4208
rect 20767 4168 20812 4196
rect 20806 4156 20812 4168
rect 20864 4156 20870 4208
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4097 12311 4131
rect 12253 4091 12311 4097
rect 12618 4088 12624 4140
rect 12676 4128 12682 4140
rect 13357 4131 13415 4137
rect 13357 4128 13369 4131
rect 12676 4100 13369 4128
rect 12676 4088 12682 4100
rect 13357 4097 13369 4100
rect 13403 4097 13415 4131
rect 13357 4091 13415 4097
rect 13446 4088 13452 4140
rect 13504 4128 13510 4140
rect 14093 4131 14151 4137
rect 14093 4128 14105 4131
rect 13504 4100 14105 4128
rect 13504 4088 13510 4100
rect 14093 4097 14105 4100
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 15105 4131 15163 4137
rect 15105 4097 15117 4131
rect 15151 4128 15163 4131
rect 15286 4128 15292 4140
rect 15151 4100 15292 4128
rect 15151 4097 15163 4100
rect 15105 4091 15163 4097
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 17586 4128 17592 4140
rect 15856 4100 17592 4128
rect 8938 4020 8944 4072
rect 8996 4060 9002 4072
rect 10505 4063 10563 4069
rect 10505 4060 10517 4063
rect 8996 4032 10517 4060
rect 8996 4020 9002 4032
rect 10505 4029 10517 4032
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 8260 3964 8892 3992
rect 9309 3995 9367 4001
rect 8260 3952 8266 3964
rect 9309 3961 9321 3995
rect 9355 3992 9367 3995
rect 9398 3992 9404 4004
rect 9355 3964 9404 3992
rect 9355 3961 9367 3964
rect 9309 3955 9367 3961
rect 9398 3952 9404 3964
rect 9456 3952 9462 4004
rect 9953 3995 10011 4001
rect 9953 3961 9965 3995
rect 9999 3992 10011 3995
rect 10226 3992 10232 4004
rect 9999 3964 10232 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 10226 3952 10232 3964
rect 10284 3952 10290 4004
rect 10520 3992 10548 4023
rect 10594 4020 10600 4072
rect 10652 4060 10658 4072
rect 10781 4063 10839 4069
rect 10781 4060 10793 4063
rect 10652 4032 10793 4060
rect 10652 4020 10658 4032
rect 10781 4029 10793 4032
rect 10827 4060 10839 4063
rect 11425 4063 11483 4069
rect 11425 4060 11437 4063
rect 10827 4032 11437 4060
rect 10827 4029 10839 4032
rect 10781 4023 10839 4029
rect 11425 4029 11437 4032
rect 11471 4029 11483 4063
rect 11698 4060 11704 4072
rect 11659 4032 11704 4060
rect 11425 4023 11483 4029
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 13078 4060 13084 4072
rect 12084 4032 13084 4060
rect 10873 3995 10931 4001
rect 10873 3992 10885 3995
rect 10520 3964 10885 3992
rect 10873 3961 10885 3964
rect 10919 3961 10931 3995
rect 10873 3955 10931 3961
rect 10962 3952 10968 4004
rect 11020 3992 11026 4004
rect 11241 3995 11299 4001
rect 11241 3992 11253 3995
rect 11020 3964 11253 3992
rect 11020 3952 11026 3964
rect 11241 3961 11253 3964
rect 11287 3961 11299 3995
rect 11241 3955 11299 3961
rect 6788 3896 6868 3924
rect 6788 3884 6794 3896
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9824 3896 9873 3924
rect 9824 3884 9830 3896
rect 9861 3893 9873 3896
rect 9907 3893 9919 3927
rect 9861 3887 9919 3893
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10100 3896 10333 3924
rect 10100 3884 10106 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10321 3887 10379 3893
rect 10410 3884 10416 3936
rect 10468 3924 10474 3936
rect 10597 3927 10655 3933
rect 10597 3924 10609 3927
rect 10468 3896 10609 3924
rect 10468 3884 10474 3896
rect 10597 3893 10609 3896
rect 10643 3893 10655 3927
rect 10597 3887 10655 3893
rect 11885 3927 11943 3933
rect 11885 3893 11897 3927
rect 11931 3924 11943 3927
rect 12084 3924 12112 4032
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13173 4063 13231 4069
rect 13173 4029 13185 4063
rect 13219 4060 13231 4063
rect 13262 4060 13268 4072
rect 13219 4032 13268 4060
rect 13219 4029 13231 4032
rect 13173 4023 13231 4029
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4029 13691 4063
rect 13633 4023 13691 4029
rect 14369 4063 14427 4069
rect 14369 4029 14381 4063
rect 14415 4060 14427 4063
rect 14458 4060 14464 4072
rect 14415 4032 14464 4060
rect 14415 4029 14427 4032
rect 14369 4023 14427 4029
rect 12526 3952 12532 4004
rect 12584 3992 12590 4004
rect 13648 3992 13676 4023
rect 14458 4020 14464 4032
rect 14516 4020 14522 4072
rect 14642 4060 14648 4072
rect 14603 4032 14648 4060
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 15856 4060 15884 4100
rect 17586 4088 17592 4100
rect 17644 4088 17650 4140
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4128 19119 4131
rect 19150 4128 19156 4140
rect 19107 4100 19156 4128
rect 19107 4097 19119 4100
rect 19061 4091 19119 4097
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 19794 4128 19800 4140
rect 19260 4100 19800 4128
rect 14844 4032 15884 4060
rect 12584 3964 13676 3992
rect 12584 3952 12590 3964
rect 13722 3952 13728 4004
rect 13780 3992 13786 4004
rect 13909 3995 13967 4001
rect 13909 3992 13921 3995
rect 13780 3964 13921 3992
rect 13780 3952 13786 3964
rect 13909 3961 13921 3964
rect 13955 3961 13967 3995
rect 13909 3955 13967 3961
rect 14384 3964 14688 3992
rect 11931 3896 12112 3924
rect 11931 3893 11943 3896
rect 11885 3887 11943 3893
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 12216 3896 12357 3924
rect 12216 3884 12222 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12710 3924 12716 3936
rect 12671 3896 12716 3924
rect 12345 3887 12403 3893
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 12802 3884 12808 3936
rect 12860 3924 12866 3936
rect 13265 3927 13323 3933
rect 12860 3896 12905 3924
rect 12860 3884 12866 3896
rect 13265 3893 13277 3927
rect 13311 3924 13323 3927
rect 13354 3924 13360 3936
rect 13311 3896 13360 3924
rect 13311 3893 13323 3896
rect 13265 3887 13323 3893
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 14384 3924 14412 3964
rect 14660 3936 14688 3964
rect 14550 3924 14556 3936
rect 13863 3896 14412 3924
rect 14511 3896 14556 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 14642 3884 14648 3936
rect 14700 3884 14706 3936
rect 14844 3933 14872 4032
rect 15930 4020 15936 4072
rect 15988 4060 15994 4072
rect 16301 4063 16359 4069
rect 15988 4032 16033 4060
rect 15988 4020 15994 4032
rect 16301 4029 16313 4063
rect 16347 4060 16359 4063
rect 16390 4060 16396 4072
rect 16347 4032 16396 4060
rect 16347 4029 16359 4032
rect 16301 4023 16359 4029
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 16574 4060 16580 4072
rect 16535 4032 16580 4060
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 16942 4060 16948 4072
rect 16903 4032 16948 4060
rect 16942 4020 16948 4032
rect 17000 4020 17006 4072
rect 17405 4063 17463 4069
rect 17405 4029 17417 4063
rect 17451 4060 17463 4063
rect 17954 4060 17960 4072
rect 17451 4032 17960 4060
rect 17451 4029 17463 4032
rect 17405 4023 17463 4029
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 18794 4063 18852 4069
rect 18794 4029 18806 4063
rect 18840 4060 18852 4063
rect 19260 4060 19288 4100
rect 19794 4088 19800 4100
rect 19852 4088 19858 4140
rect 19978 4128 19984 4140
rect 19939 4100 19984 4128
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20070 4088 20076 4140
rect 20128 4128 20134 4140
rect 20128 4100 21312 4128
rect 20128 4088 20134 4100
rect 21284 4072 21312 4100
rect 18840 4032 19288 4060
rect 18840 4029 18852 4032
rect 18794 4023 18852 4029
rect 18892 4004 18920 4032
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 20257 4063 20315 4069
rect 19392 4032 20208 4060
rect 19392 4020 19398 4032
rect 15289 3995 15347 4001
rect 15289 3961 15301 3995
rect 15335 3992 15347 3995
rect 15378 3992 15384 4004
rect 15335 3964 15384 3992
rect 15335 3961 15347 3964
rect 15289 3955 15347 3961
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 15672 3964 18837 3992
rect 14829 3927 14887 3933
rect 14829 3893 14841 3927
rect 14875 3893 14887 3927
rect 15194 3924 15200 3936
rect 15155 3896 15200 3924
rect 14829 3887 14887 3893
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 15672 3933 15700 3964
rect 15657 3927 15715 3933
rect 15657 3893 15669 3927
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 16117 3927 16175 3933
rect 16117 3893 16129 3927
rect 16163 3924 16175 3927
rect 16298 3924 16304 3936
rect 16163 3896 16304 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 16482 3924 16488 3936
rect 16443 3896 16488 3924
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 16758 3924 16764 3936
rect 16719 3896 16764 3924
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 17126 3924 17132 3936
rect 17087 3896 17132 3924
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 17589 3927 17647 3933
rect 17589 3893 17601 3927
rect 17635 3924 17647 3927
rect 18690 3924 18696 3936
rect 17635 3896 18696 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 18690 3884 18696 3896
rect 18748 3884 18754 3936
rect 18809 3924 18837 3964
rect 18874 3952 18880 4004
rect 18932 3952 18938 4004
rect 19613 3995 19671 4001
rect 19613 3992 19625 3995
rect 19306 3964 19625 3992
rect 19306 3924 19334 3964
rect 19613 3961 19625 3964
rect 19659 3961 19671 3995
rect 20180 3992 20208 4032
rect 20257 4029 20269 4063
rect 20303 4060 20315 4063
rect 20438 4060 20444 4072
rect 20303 4032 20444 4060
rect 20303 4029 20315 4032
rect 20257 4023 20315 4029
rect 20438 4020 20444 4032
rect 20496 4020 20502 4072
rect 20714 4060 20720 4072
rect 20675 4032 20720 4060
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 20993 4063 21051 4069
rect 20993 4029 21005 4063
rect 21039 4029 21051 4063
rect 21266 4060 21272 4072
rect 21227 4032 21272 4060
rect 20993 4023 21051 4029
rect 21008 3992 21036 4023
rect 21266 4020 21272 4032
rect 21324 4020 21330 4072
rect 21542 4060 21548 4072
rect 21503 4032 21548 4060
rect 21542 4020 21548 4032
rect 21600 4020 21606 4072
rect 22005 3995 22063 4001
rect 22005 3992 22017 3995
rect 20180 3964 22017 3992
rect 19613 3955 19671 3961
rect 22005 3961 22017 3964
rect 22051 3961 22063 3995
rect 22005 3955 22063 3961
rect 19518 3924 19524 3936
rect 18809 3896 19334 3924
rect 19479 3896 19524 3924
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 19702 3884 19708 3936
rect 19760 3924 19766 3936
rect 20533 3927 20591 3933
rect 20533 3924 20545 3927
rect 19760 3896 20545 3924
rect 19760 3884 19766 3896
rect 20533 3893 20545 3896
rect 20579 3893 20591 3927
rect 20533 3887 20591 3893
rect 20898 3884 20904 3936
rect 20956 3924 20962 3936
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 20956 3896 21097 3924
rect 20956 3884 20962 3896
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 21085 3887 21143 3893
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3924 21419 3927
rect 22094 3924 22100 3936
rect 21407 3896 22100 3924
rect 21407 3893 21419 3896
rect 21361 3887 21419 3893
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 2038 3720 2044 3732
rect 1627 3692 2044 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 2222 3720 2228 3732
rect 2179 3692 2228 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 2961 3723 3019 3729
rect 2961 3689 2973 3723
rect 3007 3720 3019 3723
rect 3418 3720 3424 3732
rect 3007 3692 3424 3720
rect 3007 3689 3019 3692
rect 2961 3683 3019 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 4249 3723 4307 3729
rect 4249 3689 4261 3723
rect 4295 3720 4307 3723
rect 4338 3720 4344 3732
rect 4295 3692 4344 3720
rect 4295 3689 4307 3692
rect 4249 3683 4307 3689
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 5442 3720 5448 3732
rect 4448 3692 5448 3720
rect 2774 3652 2780 3664
rect 1688 3624 2780 3652
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 1688 3593 1716 3624
rect 2774 3612 2780 3624
rect 2832 3612 2838 3664
rect 3329 3655 3387 3661
rect 3329 3621 3341 3655
rect 3375 3652 3387 3655
rect 4448 3652 4476 3692
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 6273 3723 6331 3729
rect 6273 3689 6285 3723
rect 6319 3720 6331 3723
rect 8205 3723 8263 3729
rect 8205 3720 8217 3723
rect 6319 3692 8217 3720
rect 6319 3689 6331 3692
rect 6273 3683 6331 3689
rect 8205 3689 8217 3692
rect 8251 3689 8263 3723
rect 8205 3683 8263 3689
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 8754 3720 8760 3732
rect 8352 3692 8760 3720
rect 8352 3680 8358 3692
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 9309 3723 9367 3729
rect 9309 3720 9321 3723
rect 9088 3692 9321 3720
rect 9088 3680 9094 3692
rect 9309 3689 9321 3692
rect 9355 3689 9367 3723
rect 9309 3683 9367 3689
rect 9766 3680 9772 3732
rect 9824 3720 9830 3732
rect 10318 3720 10324 3732
rect 9824 3692 10324 3720
rect 9824 3680 9830 3692
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 11974 3680 11980 3732
rect 12032 3720 12038 3732
rect 12526 3720 12532 3732
rect 12032 3692 12532 3720
rect 12032 3680 12038 3692
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 12710 3720 12716 3732
rect 12671 3692 12716 3720
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 14182 3720 14188 3732
rect 12820 3692 14188 3720
rect 3375 3624 4476 3652
rect 3375 3621 3387 3624
rect 3329 3615 3387 3621
rect 4706 3612 4712 3664
rect 4764 3652 4770 3664
rect 4764 3624 5212 3652
rect 4764 3612 4770 3624
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3553 1731 3587
rect 1673 3547 1731 3553
rect 2501 3587 2559 3593
rect 2501 3553 2513 3587
rect 2547 3584 2559 3587
rect 2866 3584 2872 3596
rect 2547 3556 2872 3584
rect 2547 3553 2559 3556
rect 2501 3547 2559 3553
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 3421 3587 3479 3593
rect 3421 3553 3433 3587
rect 3467 3584 3479 3587
rect 4522 3584 4528 3596
rect 3467 3556 4528 3584
rect 3467 3553 3479 3556
rect 3421 3547 3479 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 4890 3584 4896 3596
rect 4632 3556 4896 3584
rect 2590 3516 2596 3528
rect 2551 3488 2596 3516
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 2682 3476 2688 3528
rect 2740 3516 2746 3528
rect 3602 3516 3608 3528
rect 2740 3488 2785 3516
rect 3563 3488 3608 3516
rect 2740 3476 2746 3488
rect 3602 3476 3608 3488
rect 3660 3476 3666 3528
rect 3878 3516 3884 3528
rect 3839 3488 3884 3516
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 3970 3476 3976 3528
rect 4028 3516 4034 3528
rect 4632 3516 4660 3556
rect 4890 3544 4896 3556
rect 4948 3544 4954 3596
rect 5184 3584 5212 3624
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 5362 3655 5420 3661
rect 5362 3652 5374 3655
rect 5316 3624 5374 3652
rect 5316 3612 5322 3624
rect 5362 3621 5374 3624
rect 5408 3621 5420 3655
rect 5362 3615 5420 3621
rect 5718 3612 5724 3664
rect 5776 3652 5782 3664
rect 6086 3652 6092 3664
rect 5776 3624 6092 3652
rect 5776 3612 5782 3624
rect 6086 3612 6092 3624
rect 6144 3612 6150 3664
rect 6181 3655 6239 3661
rect 6181 3621 6193 3655
rect 6227 3652 6239 3655
rect 7466 3652 7472 3664
rect 6227 3624 7472 3652
rect 6227 3621 6239 3624
rect 6181 3615 6239 3621
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 9214 3652 9220 3664
rect 8404 3624 8708 3652
rect 9175 3624 9220 3652
rect 5629 3587 5687 3593
rect 5629 3584 5641 3587
rect 5184 3556 5641 3584
rect 5629 3553 5641 3556
rect 5675 3553 5687 3587
rect 5629 3547 5687 3553
rect 7098 3544 7104 3596
rect 7156 3584 7162 3596
rect 7846 3587 7904 3593
rect 7846 3584 7858 3587
rect 7156 3556 7858 3584
rect 7156 3544 7162 3556
rect 7846 3553 7858 3556
rect 7892 3584 7904 3587
rect 8202 3584 8208 3596
rect 7892 3556 8208 3584
rect 7892 3553 7904 3556
rect 7846 3547 7904 3553
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 5994 3516 6000 3528
rect 4028 3488 4660 3516
rect 5955 3488 6000 3516
rect 4028 3476 4034 3488
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 6914 3516 6920 3528
rect 6144 3488 6920 3516
rect 6144 3476 6150 3488
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 8110 3516 8116 3528
rect 8023 3488 8116 3516
rect 8110 3476 8116 3488
rect 8168 3516 8174 3528
rect 8404 3516 8432 3624
rect 8570 3584 8576 3596
rect 8531 3556 8576 3584
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 8680 3584 8708 3624
rect 9214 3612 9220 3624
rect 9272 3612 9278 3664
rect 10042 3612 10048 3664
rect 10100 3652 10106 3664
rect 10778 3652 10784 3664
rect 10100 3624 10784 3652
rect 10100 3612 10106 3624
rect 10778 3612 10784 3624
rect 10836 3612 10842 3664
rect 12434 3612 12440 3664
rect 12492 3652 12498 3664
rect 12820 3661 12848 3692
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 14921 3723 14979 3729
rect 14921 3720 14933 3723
rect 14792 3692 14933 3720
rect 14792 3680 14798 3692
rect 14921 3689 14933 3692
rect 14967 3689 14979 3723
rect 14921 3683 14979 3689
rect 15381 3723 15439 3729
rect 15381 3689 15393 3723
rect 15427 3720 15439 3723
rect 18693 3723 18751 3729
rect 15427 3692 18644 3720
rect 15427 3689 15439 3692
rect 15381 3683 15439 3689
rect 12805 3655 12863 3661
rect 12805 3652 12817 3655
rect 12492 3624 12817 3652
rect 12492 3612 12498 3624
rect 12805 3621 12817 3624
rect 12851 3621 12863 3655
rect 12805 3615 12863 3621
rect 12894 3612 12900 3664
rect 12952 3612 12958 3664
rect 13633 3655 13691 3661
rect 13633 3621 13645 3655
rect 13679 3652 13691 3655
rect 13679 3624 13860 3652
rect 13679 3621 13691 3624
rect 13633 3615 13691 3621
rect 10617 3587 10675 3593
rect 8680 3556 9812 3584
rect 8168 3488 8432 3516
rect 8168 3476 8174 3488
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8665 3519 8723 3525
rect 8665 3516 8677 3519
rect 8536 3488 8677 3516
rect 8536 3476 8542 3488
rect 8665 3485 8677 3488
rect 8711 3485 8723 3519
rect 8665 3479 8723 3485
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 1857 3451 1915 3457
rect 1857 3417 1869 3451
rect 1903 3448 1915 3451
rect 2498 3448 2504 3460
rect 1903 3420 2504 3448
rect 1903 3417 1915 3420
rect 1857 3411 1915 3417
rect 2498 3408 2504 3420
rect 2556 3408 2562 3460
rect 2746 3420 4384 3448
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 1949 3383 2007 3389
rect 1949 3380 1961 3383
rect 1728 3352 1961 3380
rect 1728 3340 1734 3352
rect 1949 3349 1961 3352
rect 1995 3349 2007 3383
rect 1949 3343 2007 3349
rect 2222 3340 2228 3392
rect 2280 3380 2286 3392
rect 2746 3380 2774 3420
rect 2280 3352 2774 3380
rect 2280 3340 2286 3352
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 3418 3380 3424 3392
rect 3292 3352 3424 3380
rect 3292 3340 3298 3352
rect 3418 3340 3424 3352
rect 3476 3340 3482 3392
rect 4356 3380 4384 3420
rect 5721 3383 5779 3389
rect 5721 3380 5733 3383
rect 4356 3352 5733 3380
rect 5721 3349 5733 3352
rect 5767 3349 5779 3383
rect 6012 3380 6040 3476
rect 6641 3451 6699 3457
rect 6641 3417 6653 3451
rect 6687 3448 6699 3451
rect 6822 3448 6828 3460
rect 6687 3420 6828 3448
rect 6687 3417 6699 3420
rect 6641 3411 6699 3417
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 8202 3408 8208 3460
rect 8260 3448 8266 3460
rect 8772 3448 8800 3479
rect 8260 3420 8800 3448
rect 8260 3408 8266 3420
rect 6730 3380 6736 3392
rect 6012 3352 6736 3380
rect 5721 3343 5779 3349
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 7742 3340 7748 3392
rect 7800 3380 7806 3392
rect 9214 3380 9220 3392
rect 7800 3352 9220 3380
rect 7800 3340 7806 3352
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 9493 3383 9551 3389
rect 9493 3349 9505 3383
rect 9539 3380 9551 3383
rect 9674 3380 9680 3392
rect 9539 3352 9680 3380
rect 9539 3349 9551 3352
rect 9493 3343 9551 3349
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 9784 3380 9812 3556
rect 10617 3553 10629 3587
rect 10663 3584 10675 3587
rect 10663 3556 11008 3584
rect 10663 3553 10675 3556
rect 10617 3547 10675 3553
rect 10873 3519 10931 3525
rect 10873 3485 10885 3519
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 10686 3380 10692 3392
rect 9784 3352 10692 3380
rect 10686 3340 10692 3352
rect 10744 3380 10750 3392
rect 10888 3380 10916 3479
rect 10980 3389 11008 3556
rect 11698 3544 11704 3596
rect 11756 3584 11762 3596
rect 12078 3587 12136 3593
rect 12078 3584 12090 3587
rect 11756 3556 12090 3584
rect 11756 3544 11762 3556
rect 12078 3553 12090 3556
rect 12124 3553 12136 3587
rect 12078 3547 12136 3553
rect 12345 3587 12403 3593
rect 12345 3553 12357 3587
rect 12391 3584 12403 3587
rect 12912 3584 12940 3612
rect 13354 3584 13360 3596
rect 12391 3556 13360 3584
rect 12391 3553 12403 3556
rect 12345 3547 12403 3553
rect 13354 3544 13360 3556
rect 13412 3544 13418 3596
rect 13538 3544 13544 3596
rect 13596 3584 13602 3596
rect 13725 3587 13783 3593
rect 13725 3584 13737 3587
rect 13596 3556 13737 3584
rect 13596 3544 13602 3556
rect 13725 3553 13737 3556
rect 13771 3553 13783 3587
rect 13832 3584 13860 3624
rect 14090 3612 14096 3664
rect 14148 3652 14154 3664
rect 14148 3624 14504 3652
rect 14148 3612 14154 3624
rect 14369 3587 14427 3593
rect 14369 3584 14381 3587
rect 13832 3556 14381 3584
rect 13725 3547 13783 3553
rect 14369 3553 14381 3556
rect 14415 3553 14427 3587
rect 14476 3584 14504 3624
rect 14550 3612 14556 3664
rect 14608 3652 14614 3664
rect 14608 3624 15792 3652
rect 14608 3612 14614 3624
rect 15013 3587 15071 3593
rect 15013 3584 15025 3587
rect 14476 3556 15025 3584
rect 14369 3547 14427 3553
rect 15013 3553 15025 3556
rect 15059 3584 15071 3587
rect 15102 3584 15108 3596
rect 15059 3556 15108 3584
rect 15059 3553 15071 3556
rect 15013 3547 15071 3553
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 15764 3593 15792 3624
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 18616 3652 18644 3692
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 18782 3720 18788 3732
rect 18739 3692 18788 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 18782 3680 18788 3692
rect 18840 3680 18846 3732
rect 20073 3723 20131 3729
rect 20073 3720 20085 3723
rect 18892 3692 20085 3720
rect 18892 3652 18920 3692
rect 20073 3689 20085 3692
rect 20119 3689 20131 3723
rect 20073 3683 20131 3689
rect 20530 3652 20536 3664
rect 17184 3624 17908 3652
rect 18616 3624 18920 3652
rect 19352 3624 20536 3652
rect 17184 3612 17190 3624
rect 15473 3587 15531 3593
rect 15473 3553 15485 3587
rect 15519 3553 15531 3587
rect 15473 3547 15531 3553
rect 15749 3587 15807 3593
rect 15749 3553 15761 3587
rect 15795 3553 15807 3587
rect 15749 3547 15807 3553
rect 12618 3516 12624 3528
rect 12579 3488 12624 3516
rect 12618 3476 12624 3488
rect 12676 3516 12682 3528
rect 12894 3516 12900 3528
rect 12676 3488 12900 3516
rect 12676 3476 12682 3488
rect 12894 3476 12900 3488
rect 12952 3516 12958 3528
rect 13817 3519 13875 3525
rect 13817 3516 13829 3519
rect 12952 3488 13829 3516
rect 12952 3476 12958 3488
rect 13817 3485 13829 3488
rect 13863 3485 13875 3519
rect 13817 3479 13875 3485
rect 14829 3519 14887 3525
rect 14829 3485 14841 3519
rect 14875 3485 14887 3519
rect 15488 3516 15516 3547
rect 17218 3544 17224 3596
rect 17276 3593 17282 3596
rect 17276 3584 17288 3593
rect 17586 3584 17592 3596
rect 17276 3556 17321 3584
rect 17547 3556 17592 3584
rect 17276 3547 17288 3556
rect 17276 3544 17282 3547
rect 17586 3544 17592 3556
rect 17644 3544 17650 3596
rect 17880 3593 17908 3624
rect 17865 3587 17923 3593
rect 17865 3553 17877 3587
rect 17911 3553 17923 3587
rect 18230 3584 18236 3596
rect 17865 3547 17923 3553
rect 17972 3556 18236 3584
rect 16206 3516 16212 3528
rect 15488 3488 16212 3516
rect 14829 3479 14887 3485
rect 12986 3408 12992 3460
rect 13044 3448 13050 3460
rect 14093 3451 14151 3457
rect 14093 3448 14105 3451
rect 13044 3420 14105 3448
rect 13044 3408 13050 3420
rect 14093 3417 14105 3420
rect 14139 3417 14151 3451
rect 14844 3448 14872 3479
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 17497 3519 17555 3525
rect 17497 3485 17509 3519
rect 17543 3516 17555 3519
rect 17972 3516 18000 3556
rect 18230 3544 18236 3556
rect 18288 3544 18294 3596
rect 18506 3544 18512 3596
rect 18564 3584 18570 3596
rect 19153 3587 19211 3593
rect 19153 3584 19165 3587
rect 18564 3556 19165 3584
rect 18564 3544 18570 3556
rect 19153 3553 19165 3556
rect 19199 3553 19211 3587
rect 19153 3547 19211 3553
rect 17543 3488 18000 3516
rect 17543 3485 17555 3488
rect 17497 3479 17555 3485
rect 17604 3460 17632 3488
rect 18138 3476 18144 3528
rect 18196 3516 18202 3528
rect 18417 3519 18475 3525
rect 18417 3516 18429 3519
rect 18196 3488 18429 3516
rect 18196 3476 18202 3488
rect 18417 3485 18429 3488
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 18601 3519 18659 3525
rect 18601 3485 18613 3519
rect 18647 3516 18659 3519
rect 19352 3516 19380 3624
rect 20530 3612 20536 3624
rect 20588 3612 20594 3664
rect 21358 3652 21364 3664
rect 21319 3624 21364 3652
rect 21358 3612 21364 3624
rect 21416 3612 21422 3664
rect 19978 3584 19984 3596
rect 19939 3556 19984 3584
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 20441 3587 20499 3593
rect 20441 3553 20453 3587
rect 20487 3584 20499 3587
rect 20622 3584 20628 3596
rect 20487 3556 20628 3584
rect 20487 3553 20499 3556
rect 20441 3547 20499 3553
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 20993 3587 21051 3593
rect 20993 3553 21005 3587
rect 21039 3584 21051 3587
rect 21634 3584 21640 3596
rect 21039 3556 21640 3584
rect 21039 3553 21051 3556
rect 20993 3547 21051 3553
rect 21634 3544 21640 3556
rect 21692 3544 21698 3596
rect 18647 3488 19380 3516
rect 18647 3485 18659 3488
rect 18601 3479 18659 3485
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 19576 3488 19748 3516
rect 19576 3476 19582 3488
rect 15286 3448 15292 3460
rect 14844 3420 15292 3448
rect 14093 3411 14151 3417
rect 15286 3408 15292 3420
rect 15344 3448 15350 3460
rect 16117 3451 16175 3457
rect 16117 3448 16129 3451
rect 15344 3420 16129 3448
rect 15344 3408 15350 3420
rect 16117 3417 16129 3420
rect 16163 3448 16175 3451
rect 16390 3448 16396 3460
rect 16163 3420 16396 3448
rect 16163 3417 16175 3420
rect 16117 3411 16175 3417
rect 16390 3408 16396 3420
rect 16448 3408 16454 3460
rect 17586 3408 17592 3460
rect 17644 3408 17650 3460
rect 18049 3451 18107 3457
rect 18049 3417 18061 3451
rect 18095 3448 18107 3451
rect 19610 3448 19616 3460
rect 18095 3420 19472 3448
rect 19571 3420 19616 3448
rect 18095 3417 18107 3420
rect 18049 3411 18107 3417
rect 10744 3352 10916 3380
rect 10965 3383 11023 3389
rect 10744 3340 10750 3352
rect 10965 3349 10977 3383
rect 11011 3380 11023 3383
rect 11054 3380 11060 3392
rect 11011 3352 11060 3380
rect 11011 3349 11023 3352
rect 10965 3343 11023 3349
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 13170 3380 13176 3392
rect 13131 3352 13176 3380
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 13265 3383 13323 3389
rect 13265 3349 13277 3383
rect 13311 3380 13323 3383
rect 13538 3380 13544 3392
rect 13311 3352 13544 3380
rect 13311 3349 13323 3352
rect 13265 3343 13323 3349
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 15657 3383 15715 3389
rect 15657 3349 15669 3383
rect 15703 3380 15715 3383
rect 15838 3380 15844 3392
rect 15703 3352 15844 3380
rect 15703 3349 15715 3352
rect 15657 3343 15715 3349
rect 15838 3340 15844 3352
rect 15896 3340 15902 3392
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 15988 3352 16033 3380
rect 15988 3340 15994 3352
rect 16298 3340 16304 3392
rect 16356 3380 16362 3392
rect 17310 3380 17316 3392
rect 16356 3352 17316 3380
rect 16356 3340 16362 3352
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 17678 3340 17684 3392
rect 17736 3380 17742 3392
rect 17773 3383 17831 3389
rect 17773 3380 17785 3383
rect 17736 3352 17785 3380
rect 17736 3340 17742 3352
rect 17773 3349 17785 3352
rect 17819 3349 17831 3383
rect 17773 3343 17831 3349
rect 18233 3383 18291 3389
rect 18233 3349 18245 3383
rect 18279 3380 18291 3383
rect 18782 3380 18788 3392
rect 18279 3352 18788 3380
rect 18279 3349 18291 3352
rect 18233 3343 18291 3349
rect 18782 3340 18788 3352
rect 18840 3340 18846 3392
rect 19058 3380 19064 3392
rect 19019 3352 19064 3380
rect 19058 3340 19064 3352
rect 19116 3340 19122 3392
rect 19334 3380 19340 3392
rect 19295 3352 19340 3380
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 19444 3380 19472 3420
rect 19610 3408 19616 3420
rect 19668 3408 19674 3460
rect 19720 3448 19748 3488
rect 19794 3476 19800 3528
rect 19852 3516 19858 3528
rect 20165 3519 20223 3525
rect 20165 3516 20177 3519
rect 19852 3488 20177 3516
rect 19852 3476 19858 3488
rect 20165 3485 20177 3488
rect 20211 3485 20223 3519
rect 20165 3479 20223 3485
rect 20809 3519 20867 3525
rect 20809 3485 20821 3519
rect 20855 3516 20867 3519
rect 21082 3516 21088 3528
rect 20855 3488 21088 3516
rect 20855 3485 20867 3488
rect 20809 3479 20867 3485
rect 21082 3476 21088 3488
rect 21140 3476 21146 3528
rect 20254 3448 20260 3460
rect 19720 3420 20260 3448
rect 20254 3408 20260 3420
rect 20312 3408 20318 3460
rect 20990 3448 20996 3460
rect 20456 3420 20996 3448
rect 20456 3380 20484 3420
rect 20990 3408 20996 3420
rect 21048 3408 21054 3460
rect 21545 3451 21603 3457
rect 21545 3417 21557 3451
rect 21591 3448 21603 3451
rect 21910 3448 21916 3460
rect 21591 3420 21916 3448
rect 21591 3417 21603 3420
rect 21545 3411 21603 3417
rect 21910 3408 21916 3420
rect 21968 3408 21974 3460
rect 20622 3380 20628 3392
rect 19444 3352 20484 3380
rect 20583 3352 20628 3380
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 21085 3383 21143 3389
rect 21085 3349 21097 3383
rect 21131 3380 21143 3383
rect 22738 3380 22744 3392
rect 21131 3352 22744 3380
rect 21131 3349 21143 3352
rect 21085 3343 21143 3349
rect 22738 3340 22744 3352
rect 22796 3340 22802 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 2590 3136 2596 3188
rect 2648 3176 2654 3188
rect 3053 3179 3111 3185
rect 3053 3176 3065 3179
rect 2648 3148 3065 3176
rect 2648 3136 2654 3148
rect 3053 3145 3065 3148
rect 3099 3145 3111 3179
rect 3053 3139 3111 3145
rect 3694 3136 3700 3188
rect 3752 3176 3758 3188
rect 5074 3176 5080 3188
rect 3752 3148 5080 3176
rect 3752 3136 3758 3148
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5261 3179 5319 3185
rect 5261 3145 5273 3179
rect 5307 3176 5319 3179
rect 5718 3176 5724 3188
rect 5307 3148 5724 3176
rect 5307 3145 5319 3148
rect 5261 3139 5319 3145
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 6273 3179 6331 3185
rect 6273 3176 6285 3179
rect 5868 3148 6285 3176
rect 5868 3136 5874 3148
rect 6273 3145 6285 3148
rect 6319 3145 6331 3179
rect 6273 3139 6331 3145
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 8294 3176 8300 3188
rect 6696 3148 8300 3176
rect 6696 3136 6702 3148
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 8478 3176 8484 3188
rect 8439 3148 8484 3176
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 9766 3176 9772 3188
rect 9600 3148 9772 3176
rect 1581 3111 1639 3117
rect 1581 3077 1593 3111
rect 1627 3108 1639 3111
rect 3510 3108 3516 3120
rect 1627 3080 3372 3108
rect 1627 3077 1639 3080
rect 1581 3071 1639 3077
rect 2130 3040 2136 3052
rect 1412 3012 2136 3040
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 1412 2981 1440 3012
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 1360 2944 1409 2972
rect 1360 2932 1366 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1854 2972 1860 2984
rect 1815 2944 1860 2972
rect 1397 2935 1455 2941
rect 1854 2932 1860 2944
rect 1912 2932 1918 2984
rect 2222 2972 2228 2984
rect 2183 2944 2228 2972
rect 2222 2932 2228 2944
rect 2280 2932 2286 2984
rect 2682 2972 2688 2984
rect 2595 2944 2688 2972
rect 2682 2932 2688 2944
rect 2740 2972 2746 2984
rect 3142 2972 3148 2984
rect 2740 2944 3148 2972
rect 2740 2932 2746 2944
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 198 2864 204 2916
rect 256 2904 262 2916
rect 1486 2904 1492 2916
rect 256 2876 1492 2904
rect 256 2864 262 2876
rect 1486 2864 1492 2876
rect 1544 2904 1550 2916
rect 1673 2907 1731 2913
rect 1673 2904 1685 2907
rect 1544 2876 1685 2904
rect 1544 2864 1550 2876
rect 1673 2873 1685 2876
rect 1719 2873 1731 2907
rect 3234 2904 3240 2916
rect 1673 2867 1731 2873
rect 2884 2876 3240 2904
rect 2406 2836 2412 2848
rect 2367 2808 2412 2836
rect 2406 2796 2412 2808
rect 2464 2796 2470 2848
rect 2498 2796 2504 2848
rect 2556 2836 2562 2848
rect 2884 2845 2912 2876
rect 3234 2864 3240 2876
rect 3292 2864 3298 2916
rect 3344 2904 3372 3080
rect 3436 3080 3516 3108
rect 3436 2972 3464 3080
rect 3510 3068 3516 3080
rect 3568 3068 3574 3120
rect 5442 3068 5448 3120
rect 5500 3108 5506 3120
rect 6086 3108 6092 3120
rect 5500 3080 6092 3108
rect 5500 3068 5506 3080
rect 6086 3068 6092 3080
rect 6144 3068 6150 3120
rect 6362 3068 6368 3120
rect 6420 3108 6426 3120
rect 6457 3111 6515 3117
rect 6457 3108 6469 3111
rect 6420 3080 6469 3108
rect 6420 3068 6426 3080
rect 6457 3077 6469 3080
rect 6503 3077 6515 3111
rect 6457 3071 6515 3077
rect 6825 3111 6883 3117
rect 6825 3077 6837 3111
rect 6871 3108 6883 3111
rect 7098 3108 7104 3120
rect 6871 3080 7104 3108
rect 6871 3077 6883 3080
rect 6825 3071 6883 3077
rect 3602 3040 3608 3052
rect 3563 3012 3608 3040
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3844 3012 3893 3040
rect 3844 3000 3850 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3040 5779 3043
rect 6840 3040 6868 3071
rect 7098 3068 7104 3080
rect 7156 3068 7162 3120
rect 8202 3068 8208 3120
rect 8260 3108 8266 3120
rect 9398 3108 9404 3120
rect 8260 3080 9404 3108
rect 8260 3068 8266 3080
rect 9398 3068 9404 3080
rect 9456 3068 9462 3120
rect 8754 3040 8760 3052
rect 5767 3012 6868 3040
rect 8128 3012 8760 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 4154 2981 4160 2984
rect 3513 2975 3571 2981
rect 3513 2972 3525 2975
rect 3436 2944 3525 2972
rect 3513 2941 3525 2944
rect 3559 2941 3571 2975
rect 4148 2972 4160 2981
rect 4115 2944 4160 2972
rect 3513 2935 3571 2941
rect 4148 2935 4160 2944
rect 4154 2932 4160 2935
rect 4212 2932 4218 2984
rect 4706 2932 4712 2984
rect 4764 2972 4770 2984
rect 5166 2972 5172 2984
rect 4764 2944 5172 2972
rect 4764 2932 4770 2944
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 5905 2975 5963 2981
rect 5905 2941 5917 2975
rect 5951 2972 5963 2975
rect 7650 2972 7656 2984
rect 5951 2944 7656 2972
rect 5951 2941 5963 2944
rect 5905 2935 5963 2941
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 7949 2975 8007 2981
rect 7949 2941 7961 2975
rect 7995 2972 8007 2975
rect 8128 2972 8156 3012
rect 8754 3000 8760 3012
rect 8812 3040 8818 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8812 3012 9045 3040
rect 8812 3000 8818 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 7995 2944 8156 2972
rect 8205 2975 8263 2981
rect 7995 2941 8007 2944
rect 7949 2935 8007 2941
rect 8205 2941 8217 2975
rect 8251 2941 8263 2975
rect 8846 2972 8852 2984
rect 8759 2944 8852 2972
rect 8205 2935 8263 2941
rect 3344 2876 4200 2904
rect 4172 2848 4200 2876
rect 4890 2864 4896 2916
rect 4948 2904 4954 2916
rect 6638 2904 6644 2916
rect 4948 2876 5948 2904
rect 6599 2876 6644 2904
rect 4948 2864 4954 2876
rect 2869 2839 2927 2845
rect 2556 2808 2601 2836
rect 2556 2796 2562 2808
rect 2869 2805 2881 2839
rect 2915 2805 2927 2839
rect 3418 2836 3424 2848
rect 3379 2808 3424 2836
rect 2869 2799 2927 2805
rect 3418 2796 3424 2808
rect 3476 2796 3482 2848
rect 4154 2796 4160 2848
rect 4212 2796 4218 2848
rect 5810 2836 5816 2848
rect 5771 2808 5816 2836
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 5920 2836 5948 2876
rect 6638 2864 6644 2876
rect 6696 2864 6702 2916
rect 6748 2876 6960 2904
rect 6748 2836 6776 2876
rect 5920 2808 6776 2836
rect 6932 2836 6960 2876
rect 8110 2864 8116 2916
rect 8168 2904 8174 2916
rect 8220 2904 8248 2935
rect 8846 2932 8852 2944
rect 8904 2972 8910 2984
rect 9600 2972 9628 3148
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10965 3179 11023 3185
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 11146 3176 11152 3188
rect 11011 3148 11152 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 11698 3176 11704 3188
rect 11659 3148 11704 3176
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 15194 3176 15200 3188
rect 11808 3148 15200 3176
rect 10778 3068 10784 3120
rect 10836 3108 10842 3120
rect 11808 3108 11836 3148
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 17586 3176 17592 3188
rect 16960 3148 17592 3176
rect 10836 3080 11836 3108
rect 10836 3068 10842 3080
rect 13078 3068 13084 3120
rect 13136 3108 13142 3120
rect 15565 3111 15623 3117
rect 13136 3080 14228 3108
rect 13136 3068 13142 3080
rect 13170 3000 13176 3052
rect 13228 3040 13234 3052
rect 13633 3043 13691 3049
rect 13633 3040 13645 3043
rect 13228 3012 13645 3040
rect 13228 3000 13234 3012
rect 13633 3009 13645 3012
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 8904 2944 9628 2972
rect 8904 2932 8910 2944
rect 9674 2932 9680 2984
rect 9732 2972 9738 2984
rect 10514 2975 10572 2981
rect 10514 2972 10526 2975
rect 9732 2944 10526 2972
rect 9732 2932 9738 2944
rect 10514 2941 10526 2944
rect 10560 2941 10572 2975
rect 10514 2935 10572 2941
rect 10686 2932 10692 2984
rect 10744 2972 10750 2984
rect 10781 2975 10839 2981
rect 10781 2972 10793 2975
rect 10744 2944 10793 2972
rect 10744 2932 10750 2944
rect 10781 2941 10793 2944
rect 10827 2941 10839 2975
rect 10781 2935 10839 2941
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 11020 2944 11253 2972
rect 11020 2932 11026 2944
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 12986 2972 12992 2984
rect 11241 2935 11299 2941
rect 12406 2944 12992 2972
rect 8168 2876 8248 2904
rect 8941 2907 8999 2913
rect 8168 2864 8174 2876
rect 8941 2873 8953 2907
rect 8987 2904 8999 2907
rect 10134 2904 10140 2916
rect 8987 2876 10140 2904
rect 8987 2873 8999 2876
rect 8941 2867 8999 2873
rect 10134 2864 10140 2876
rect 10192 2864 10198 2916
rect 10226 2864 10232 2916
rect 10284 2904 10290 2916
rect 10980 2904 11008 2932
rect 10284 2876 11008 2904
rect 11057 2907 11115 2913
rect 10284 2864 10290 2876
rect 11057 2873 11069 2907
rect 11103 2873 11115 2907
rect 11057 2867 11115 2873
rect 8297 2839 8355 2845
rect 8297 2836 8309 2839
rect 6932 2808 8309 2836
rect 8297 2805 8309 2808
rect 8343 2805 8355 2839
rect 8297 2799 8355 2805
rect 8754 2796 8760 2848
rect 8812 2836 8818 2848
rect 9401 2839 9459 2845
rect 9401 2836 9413 2839
rect 8812 2808 9413 2836
rect 8812 2796 8818 2808
rect 9401 2805 9413 2808
rect 9447 2805 9459 2839
rect 9401 2799 9459 2805
rect 9766 2796 9772 2848
rect 9824 2836 9830 2848
rect 10870 2836 10876 2848
rect 9824 2808 10876 2836
rect 9824 2796 9830 2808
rect 10870 2796 10876 2808
rect 10928 2836 10934 2848
rect 11072 2836 11100 2867
rect 11146 2864 11152 2916
rect 11204 2904 11210 2916
rect 12406 2904 12434 2944
rect 12728 2916 12756 2944
rect 12986 2932 12992 2944
rect 13044 2932 13050 2984
rect 13081 2975 13139 2981
rect 13081 2941 13093 2975
rect 13127 2972 13139 2975
rect 13354 2972 13360 2984
rect 13127 2944 13360 2972
rect 13127 2941 13139 2944
rect 13081 2935 13139 2941
rect 13354 2932 13360 2944
rect 13412 2932 13418 2984
rect 13538 2972 13544 2984
rect 13499 2944 13544 2972
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 11204 2876 12434 2904
rect 11204 2864 11210 2876
rect 12710 2864 12716 2916
rect 12768 2864 12774 2916
rect 12894 2913 12900 2916
rect 12836 2907 12900 2913
rect 12836 2873 12848 2907
rect 12882 2873 12900 2907
rect 12836 2867 12900 2873
rect 12894 2864 12900 2867
rect 12952 2864 12958 2916
rect 13740 2904 13768 3003
rect 14200 2981 14228 3080
rect 15565 3077 15577 3111
rect 15611 3108 15623 3111
rect 16574 3108 16580 3120
rect 15611 3080 16580 3108
rect 15611 3077 15623 3080
rect 15565 3071 15623 3077
rect 16574 3068 16580 3080
rect 16632 3068 16638 3120
rect 16960 3049 16988 3148
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 18325 3179 18383 3185
rect 18325 3145 18337 3179
rect 18371 3176 18383 3179
rect 18874 3176 18880 3188
rect 18371 3148 18880 3176
rect 18371 3145 18383 3148
rect 18325 3139 18383 3145
rect 18874 3136 18880 3148
rect 18932 3136 18938 3188
rect 19153 3179 19211 3185
rect 19153 3145 19165 3179
rect 19199 3176 19211 3179
rect 19978 3176 19984 3188
rect 19199 3148 19984 3176
rect 19199 3145 19211 3148
rect 19153 3139 19211 3145
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 19242 3108 19248 3120
rect 18064 3080 19248 3108
rect 18064 3052 18092 3080
rect 19242 3068 19248 3080
rect 19300 3068 19306 3120
rect 19429 3111 19487 3117
rect 19429 3077 19441 3111
rect 19475 3108 19487 3111
rect 19610 3108 19616 3120
rect 19475 3080 19616 3108
rect 19475 3077 19487 3080
rect 19429 3071 19487 3077
rect 19610 3068 19616 3080
rect 19668 3068 19674 3120
rect 19705 3111 19763 3117
rect 19705 3077 19717 3111
rect 19751 3108 19763 3111
rect 20806 3108 20812 3120
rect 19751 3080 20812 3108
rect 19751 3077 19763 3080
rect 19705 3071 19763 3077
rect 20806 3068 20812 3080
rect 20864 3068 20870 3120
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3009 17003 3043
rect 16945 3003 17003 3009
rect 18046 3000 18052 3052
rect 18104 3000 18110 3052
rect 18230 3000 18236 3052
rect 18288 3040 18294 3052
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 18288 3012 18521 3040
rect 18288 3000 18294 3012
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 18509 3003 18567 3009
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 19392 3012 20024 3040
rect 19392 3000 19398 3012
rect 14185 2975 14243 2981
rect 14185 2941 14197 2975
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 14277 2975 14335 2981
rect 14277 2941 14289 2975
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 14292 2904 14320 2935
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 14553 2975 14611 2981
rect 14553 2972 14565 2975
rect 14424 2944 14565 2972
rect 14424 2932 14430 2944
rect 14553 2941 14565 2944
rect 14599 2941 14611 2975
rect 14553 2935 14611 2941
rect 14642 2932 14648 2984
rect 14700 2972 14706 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14700 2944 14841 2972
rect 14700 2932 14706 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 15102 2972 15108 2984
rect 15063 2944 15108 2972
rect 14829 2935 14887 2941
rect 15102 2932 15108 2944
rect 15160 2932 15166 2984
rect 15378 2972 15384 2984
rect 15339 2944 15384 2972
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 15838 2972 15844 2984
rect 15799 2944 15844 2972
rect 15838 2932 15844 2944
rect 15896 2932 15902 2984
rect 15930 2932 15936 2984
rect 15988 2972 15994 2984
rect 16209 2975 16267 2981
rect 16209 2972 16221 2975
rect 15988 2944 16221 2972
rect 15988 2932 15994 2944
rect 16209 2941 16221 2944
rect 16255 2941 16267 2975
rect 16209 2935 16267 2941
rect 16482 2932 16488 2984
rect 16540 2972 16546 2984
rect 16669 2975 16727 2981
rect 16669 2972 16681 2975
rect 16540 2944 16681 2972
rect 16540 2932 16546 2944
rect 16669 2941 16681 2944
rect 16715 2941 16727 2975
rect 16669 2935 16727 2941
rect 18414 2932 18420 2984
rect 18472 2972 18478 2984
rect 19245 2975 19303 2981
rect 19245 2972 19257 2975
rect 18472 2944 19257 2972
rect 18472 2932 18478 2944
rect 19245 2941 19257 2944
rect 19291 2941 19303 2975
rect 19518 2972 19524 2984
rect 19479 2944 19524 2972
rect 19245 2935 19303 2941
rect 19518 2932 19524 2944
rect 19576 2932 19582 2984
rect 19996 2981 20024 3012
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 20680 3012 20852 3040
rect 20680 3000 20686 3012
rect 20824 2981 20852 3012
rect 19981 2975 20039 2981
rect 19981 2941 19993 2975
rect 20027 2941 20039 2975
rect 20809 2975 20867 2981
rect 19981 2935 20039 2941
rect 20088 2944 20760 2972
rect 15654 2904 15660 2916
rect 13004 2876 13768 2904
rect 13832 2876 14320 2904
rect 15615 2876 15660 2904
rect 10928 2808 11100 2836
rect 10928 2796 10934 2808
rect 11330 2796 11336 2848
rect 11388 2836 11394 2848
rect 11425 2839 11483 2845
rect 11425 2836 11437 2839
rect 11388 2808 11437 2836
rect 11388 2796 11394 2808
rect 11425 2805 11437 2808
rect 11471 2805 11483 2839
rect 11425 2799 11483 2805
rect 11698 2796 11704 2848
rect 11756 2836 11762 2848
rect 12342 2836 12348 2848
rect 11756 2808 12348 2836
rect 11756 2796 11762 2808
rect 12342 2796 12348 2808
rect 12400 2836 12406 2848
rect 13004 2836 13032 2876
rect 13170 2836 13176 2848
rect 12400 2808 13032 2836
rect 13131 2808 13176 2836
rect 12400 2796 12406 2808
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 13832 2836 13860 2876
rect 15654 2864 15660 2876
rect 15712 2864 15718 2916
rect 16022 2904 16028 2916
rect 15983 2876 16028 2904
rect 16022 2864 16028 2876
rect 16080 2864 16086 2916
rect 16390 2864 16396 2916
rect 16448 2904 16454 2916
rect 17190 2907 17248 2913
rect 17190 2904 17202 2907
rect 16448 2876 17202 2904
rect 16448 2864 16454 2876
rect 17190 2873 17202 2876
rect 17236 2904 17248 2907
rect 17236 2876 18092 2904
rect 17236 2873 17248 2876
rect 17190 2867 17248 2873
rect 13998 2836 14004 2848
rect 13320 2808 13860 2836
rect 13959 2808 14004 2836
rect 13320 2796 13326 2808
rect 13998 2796 14004 2808
rect 14056 2796 14062 2848
rect 14458 2836 14464 2848
rect 14419 2808 14464 2836
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 14734 2836 14740 2848
rect 14695 2808 14740 2836
rect 14734 2796 14740 2808
rect 14792 2796 14798 2848
rect 15013 2839 15071 2845
rect 15013 2805 15025 2839
rect 15059 2836 15071 2839
rect 15194 2836 15200 2848
rect 15059 2808 15200 2836
rect 15059 2805 15071 2808
rect 15013 2799 15071 2805
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 15289 2839 15347 2845
rect 15289 2805 15301 2839
rect 15335 2836 15347 2839
rect 15470 2836 15476 2848
rect 15335 2808 15476 2836
rect 15335 2805 15347 2808
rect 15289 2799 15347 2805
rect 15470 2796 15476 2808
rect 15528 2796 15534 2848
rect 16482 2796 16488 2848
rect 16540 2836 16546 2848
rect 16577 2839 16635 2845
rect 16577 2836 16589 2839
rect 16540 2808 16589 2836
rect 16540 2796 16546 2808
rect 16577 2805 16589 2808
rect 16623 2805 16635 2839
rect 16577 2799 16635 2805
rect 17678 2796 17684 2848
rect 17736 2836 17742 2848
rect 17954 2836 17960 2848
rect 17736 2808 17960 2836
rect 17736 2796 17742 2808
rect 17954 2796 17960 2808
rect 18012 2796 18018 2848
rect 18064 2836 18092 2876
rect 18138 2864 18144 2916
rect 18196 2904 18202 2916
rect 19334 2904 19340 2916
rect 18196 2876 19340 2904
rect 18196 2864 18202 2876
rect 19334 2864 19340 2876
rect 19392 2864 19398 2916
rect 19794 2904 19800 2916
rect 19755 2876 19800 2904
rect 19794 2864 19800 2876
rect 19852 2864 19858 2916
rect 19886 2864 19892 2916
rect 19944 2904 19950 2916
rect 20088 2904 20116 2944
rect 20254 2904 20260 2916
rect 19944 2876 20116 2904
rect 20215 2876 20260 2904
rect 19944 2864 19950 2876
rect 20254 2864 20260 2876
rect 20312 2864 20318 2916
rect 20441 2907 20499 2913
rect 20441 2873 20453 2907
rect 20487 2873 20499 2907
rect 20622 2904 20628 2916
rect 20583 2876 20628 2904
rect 20441 2867 20499 2873
rect 18230 2836 18236 2848
rect 18064 2808 18236 2836
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 18506 2796 18512 2848
rect 18564 2836 18570 2848
rect 18693 2839 18751 2845
rect 18693 2836 18705 2839
rect 18564 2808 18705 2836
rect 18564 2796 18570 2808
rect 18693 2805 18705 2808
rect 18739 2805 18751 2839
rect 18693 2799 18751 2805
rect 18785 2839 18843 2845
rect 18785 2805 18797 2839
rect 18831 2836 18843 2839
rect 19702 2836 19708 2848
rect 18831 2808 19708 2836
rect 18831 2805 18843 2808
rect 18785 2799 18843 2805
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 20456 2836 20484 2867
rect 20622 2864 20628 2876
rect 20680 2864 20686 2916
rect 20732 2904 20760 2944
rect 20809 2941 20821 2975
rect 20855 2941 20867 2975
rect 20809 2935 20867 2941
rect 21177 2975 21235 2981
rect 21177 2941 21189 2975
rect 21223 2972 21235 2975
rect 22186 2972 22192 2984
rect 21223 2944 22192 2972
rect 21223 2941 21235 2944
rect 21177 2935 21235 2941
rect 22186 2932 22192 2944
rect 22244 2932 22250 2984
rect 21361 2907 21419 2913
rect 21361 2904 21373 2907
rect 20732 2876 21373 2904
rect 21361 2873 21373 2876
rect 21407 2873 21419 2907
rect 21361 2867 21419 2873
rect 20993 2839 21051 2845
rect 20993 2836 21005 2839
rect 20456 2808 21005 2836
rect 20993 2805 21005 2808
rect 21039 2805 21051 2839
rect 21450 2836 21456 2848
rect 21411 2808 21456 2836
rect 20993 2799 21051 2805
rect 21450 2796 21456 2808
rect 21508 2796 21514 2848
rect 22002 2836 22008 2848
rect 21963 2808 22008 2836
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 1394 2592 1400 2644
rect 1452 2592 1458 2644
rect 2866 2632 2872 2644
rect 2827 2604 2872 2632
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 3510 2592 3516 2644
rect 3568 2632 3574 2644
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 3568 2604 4077 2632
rect 3568 2592 3574 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 4065 2595 4123 2601
rect 4433 2635 4491 2641
rect 4433 2601 4445 2635
rect 4479 2632 4491 2635
rect 4798 2632 4804 2644
rect 4479 2604 4804 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 5626 2632 5632 2644
rect 5587 2604 5632 2632
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6270 2632 6276 2644
rect 5736 2604 6276 2632
rect 1412 2564 1440 2592
rect 3237 2567 3295 2573
rect 1412 2536 2728 2564
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1486 2496 1492 2508
rect 1443 2468 1492 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1486 2456 1492 2468
rect 1544 2456 1550 2508
rect 1670 2496 1676 2508
rect 1583 2468 1676 2496
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 2240 2505 2268 2536
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2465 2007 2499
rect 1949 2459 2007 2465
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2465 2283 2499
rect 2590 2496 2596 2508
rect 2551 2468 2596 2496
rect 2225 2459 2283 2465
rect 566 2388 572 2440
rect 624 2428 630 2440
rect 1688 2428 1716 2456
rect 624 2400 1716 2428
rect 1964 2428 1992 2459
rect 2590 2456 2596 2468
rect 2648 2456 2654 2508
rect 2700 2496 2728 2536
rect 3237 2533 3249 2567
rect 3283 2564 3295 2567
rect 3878 2564 3884 2576
rect 3283 2536 3884 2564
rect 3283 2533 3295 2536
rect 3237 2527 3295 2533
rect 3878 2524 3884 2536
rect 3936 2524 3942 2576
rect 4154 2524 4160 2576
rect 4212 2564 4218 2576
rect 4525 2567 4583 2573
rect 4525 2564 4537 2567
rect 4212 2536 4537 2564
rect 4212 2524 4218 2536
rect 4525 2533 4537 2536
rect 4571 2564 4583 2567
rect 4706 2564 4712 2576
rect 4571 2536 4712 2564
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 5169 2567 5227 2573
rect 5169 2533 5181 2567
rect 5215 2564 5227 2567
rect 5736 2564 5764 2604
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 6730 2632 6736 2644
rect 6691 2604 6736 2632
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 7006 2632 7012 2644
rect 6967 2604 7012 2632
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 7285 2635 7343 2641
rect 7285 2601 7297 2635
rect 7331 2601 7343 2635
rect 7285 2595 7343 2601
rect 5215 2536 5764 2564
rect 5215 2533 5227 2536
rect 5169 2527 5227 2533
rect 5810 2524 5816 2576
rect 5868 2564 5874 2576
rect 7300 2564 7328 2595
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 7653 2635 7711 2641
rect 7653 2632 7665 2635
rect 7524 2604 7665 2632
rect 7524 2592 7530 2604
rect 7653 2601 7665 2604
rect 7699 2601 7711 2635
rect 7653 2595 7711 2601
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 8662 2632 8668 2644
rect 8619 2604 8668 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9088 2604 9904 2632
rect 9088 2592 9094 2604
rect 5868 2536 7328 2564
rect 5868 2524 5874 2536
rect 7558 2524 7564 2576
rect 7616 2564 7622 2576
rect 7745 2567 7803 2573
rect 7745 2564 7757 2567
rect 7616 2536 7757 2564
rect 7616 2524 7622 2536
rect 7745 2533 7757 2536
rect 7791 2533 7803 2567
rect 9582 2564 9588 2576
rect 9543 2536 9588 2564
rect 7745 2527 7803 2533
rect 9582 2524 9588 2536
rect 9640 2524 9646 2576
rect 9876 2564 9904 2604
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 10100 2604 10241 2632
rect 10100 2592 10106 2604
rect 10229 2601 10241 2604
rect 10275 2601 10287 2635
rect 10502 2632 10508 2644
rect 10463 2604 10508 2632
rect 10229 2595 10287 2601
rect 10502 2592 10508 2604
rect 10560 2592 10566 2644
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11885 2635 11943 2641
rect 11885 2632 11897 2635
rect 11287 2604 11897 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 11885 2601 11897 2604
rect 11931 2601 11943 2635
rect 11885 2595 11943 2601
rect 12158 2592 12164 2644
rect 12216 2632 12222 2644
rect 12253 2635 12311 2641
rect 12253 2632 12265 2635
rect 12216 2604 12265 2632
rect 12216 2592 12222 2604
rect 12253 2601 12265 2604
rect 12299 2601 12311 2635
rect 12253 2595 12311 2601
rect 12345 2635 12403 2641
rect 12345 2601 12357 2635
rect 12391 2632 12403 2635
rect 12434 2632 12440 2644
rect 12391 2604 12440 2632
rect 12391 2601 12403 2604
rect 12345 2595 12403 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 12802 2632 12808 2644
rect 12763 2604 12808 2632
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 13078 2592 13084 2644
rect 13136 2632 13142 2644
rect 14369 2635 14427 2641
rect 13136 2604 14320 2632
rect 13136 2592 13142 2604
rect 10137 2567 10195 2573
rect 10137 2564 10149 2567
rect 9876 2536 10149 2564
rect 10137 2533 10149 2536
rect 10183 2533 10195 2567
rect 10137 2527 10195 2533
rect 11333 2567 11391 2573
rect 11333 2533 11345 2567
rect 11379 2564 11391 2567
rect 13170 2564 13176 2576
rect 11379 2536 13176 2564
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 13722 2564 13728 2576
rect 13280 2536 13728 2564
rect 13280 2508 13308 2536
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 13998 2564 14004 2576
rect 13959 2536 14004 2564
rect 13998 2524 14004 2536
rect 14056 2524 14062 2576
rect 3973 2499 4031 2505
rect 3973 2496 3985 2499
rect 2700 2468 3985 2496
rect 3973 2465 3985 2468
rect 4019 2465 4031 2499
rect 4890 2496 4896 2508
rect 4851 2468 4896 2496
rect 3973 2459 4031 2465
rect 4890 2456 4896 2468
rect 4948 2456 4954 2508
rect 5353 2499 5411 2505
rect 5353 2465 5365 2499
rect 5399 2496 5411 2499
rect 5442 2496 5448 2508
rect 5399 2468 5448 2496
rect 5399 2465 5411 2468
rect 5353 2459 5411 2465
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5994 2496 6000 2508
rect 5955 2468 6000 2496
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6546 2456 6552 2508
rect 6604 2496 6610 2508
rect 6641 2499 6699 2505
rect 6641 2496 6653 2499
rect 6604 2468 6653 2496
rect 6604 2456 6610 2468
rect 6641 2465 6653 2468
rect 6687 2465 6699 2499
rect 7190 2496 7196 2508
rect 7151 2468 7196 2496
rect 6641 2459 6699 2465
rect 7190 2456 7196 2468
rect 7248 2456 7254 2508
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 7576 2468 8493 2496
rect 2498 2428 2504 2440
rect 1964 2400 2504 2428
rect 624 2388 630 2400
rect 1026 2320 1032 2372
rect 1084 2360 1090 2372
rect 1964 2360 1992 2400
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 3602 2428 3608 2440
rect 3559 2400 3608 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 3602 2388 3608 2400
rect 3660 2388 3666 2440
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2397 4767 2431
rect 6086 2428 6092 2440
rect 6047 2400 6092 2428
rect 4709 2391 4767 2397
rect 1084 2332 1992 2360
rect 2777 2363 2835 2369
rect 1084 2320 1090 2332
rect 2777 2329 2789 2363
rect 2823 2360 2835 2363
rect 3786 2360 3792 2372
rect 2823 2332 3792 2360
rect 2823 2329 2835 2332
rect 2777 2323 2835 2329
rect 3786 2320 3792 2332
rect 3844 2320 3850 2372
rect 4724 2360 4752 2391
rect 6086 2388 6092 2400
rect 6144 2388 6150 2440
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 5258 2360 5264 2372
rect 4724 2332 5264 2360
rect 5258 2320 5264 2332
rect 5316 2360 5322 2372
rect 6196 2360 6224 2391
rect 5316 2332 6224 2360
rect 5316 2320 5322 2332
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 1857 2295 1915 2301
rect 1857 2261 1869 2295
rect 1903 2292 1915 2295
rect 2038 2292 2044 2304
rect 1903 2264 2044 2292
rect 1903 2261 1915 2264
rect 1857 2255 1915 2261
rect 2038 2252 2044 2264
rect 2096 2252 2102 2304
rect 2130 2252 2136 2304
rect 2188 2292 2194 2304
rect 2409 2295 2467 2301
rect 2188 2264 2233 2292
rect 2188 2252 2194 2264
rect 2409 2261 2421 2295
rect 2455 2292 2467 2295
rect 4798 2292 4804 2304
rect 2455 2264 4804 2292
rect 2455 2261 2467 2264
rect 2409 2255 2467 2261
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 5077 2295 5135 2301
rect 5077 2261 5089 2295
rect 5123 2292 5135 2295
rect 7576 2292 7604 2468
rect 8481 2465 8493 2468
rect 8527 2496 8539 2499
rect 8662 2496 8668 2508
rect 8527 2468 8668 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 8662 2456 8668 2468
rect 8720 2456 8726 2508
rect 10597 2499 10655 2505
rect 8772 2468 9812 2496
rect 8772 2440 8800 2468
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8754 2428 8760 2440
rect 7975 2400 8760 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9674 2428 9680 2440
rect 9635 2400 9680 2428
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 9784 2437 9812 2468
rect 10597 2465 10609 2499
rect 10643 2465 10655 2499
rect 10597 2459 10655 2465
rect 9769 2431 9827 2437
rect 9769 2397 9781 2431
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 7650 2320 7656 2372
rect 7708 2360 7714 2372
rect 8113 2363 8171 2369
rect 8113 2360 8125 2363
rect 7708 2332 8125 2360
rect 7708 2320 7714 2332
rect 8113 2329 8125 2332
rect 8159 2329 8171 2363
rect 8113 2323 8171 2329
rect 8570 2320 8576 2372
rect 8628 2360 8634 2372
rect 9217 2363 9275 2369
rect 9217 2360 9229 2363
rect 8628 2332 9229 2360
rect 8628 2320 8634 2332
rect 9217 2329 9229 2332
rect 9263 2329 9275 2363
rect 9217 2323 9275 2329
rect 9398 2320 9404 2372
rect 9456 2360 9462 2372
rect 10612 2360 10640 2459
rect 12710 2456 12716 2508
rect 12768 2496 12774 2508
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12768 2468 12909 2496
rect 12768 2456 12774 2468
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 12986 2456 12992 2508
rect 13044 2496 13050 2508
rect 13081 2499 13139 2505
rect 13081 2496 13093 2499
rect 13044 2468 13093 2496
rect 13044 2456 13050 2468
rect 13081 2465 13093 2468
rect 13127 2465 13139 2499
rect 13262 2496 13268 2508
rect 13223 2468 13268 2496
rect 13081 2459 13139 2465
rect 13262 2456 13268 2468
rect 13320 2456 13326 2508
rect 13446 2496 13452 2508
rect 13359 2468 13452 2496
rect 11054 2428 11060 2440
rect 11015 2400 11060 2428
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 12437 2431 12495 2437
rect 12437 2428 12449 2431
rect 12400 2400 12449 2428
rect 12400 2388 12406 2400
rect 12437 2397 12449 2400
rect 12483 2397 12495 2431
rect 13372 2428 13400 2468
rect 13446 2456 13452 2468
rect 13504 2496 13510 2508
rect 13633 2499 13691 2505
rect 13633 2496 13645 2499
rect 13504 2468 13645 2496
rect 13504 2456 13510 2468
rect 13633 2465 13645 2468
rect 13679 2465 13691 2499
rect 14182 2496 14188 2508
rect 14143 2468 14188 2496
rect 13633 2459 13691 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14292 2496 14320 2604
rect 14369 2601 14381 2635
rect 14415 2632 14427 2635
rect 14415 2604 15516 2632
rect 14415 2601 14427 2604
rect 14369 2595 14427 2601
rect 14458 2524 14464 2576
rect 14516 2564 14522 2576
rect 14737 2567 14795 2573
rect 14737 2564 14749 2567
rect 14516 2536 14749 2564
rect 14516 2524 14522 2536
rect 14737 2533 14749 2536
rect 14783 2533 14795 2567
rect 14737 2527 14795 2533
rect 14826 2524 14832 2576
rect 14884 2564 14890 2576
rect 15488 2573 15516 2604
rect 17034 2592 17040 2644
rect 17092 2632 17098 2644
rect 17589 2635 17647 2641
rect 17589 2632 17601 2635
rect 17092 2604 17601 2632
rect 17092 2592 17098 2604
rect 17589 2601 17601 2604
rect 17635 2601 17647 2635
rect 17589 2595 17647 2601
rect 17954 2592 17960 2644
rect 18012 2632 18018 2644
rect 18049 2635 18107 2641
rect 18049 2632 18061 2635
rect 18012 2604 18061 2632
rect 18012 2592 18018 2604
rect 18049 2601 18061 2604
rect 18095 2601 18107 2635
rect 18049 2595 18107 2601
rect 18509 2635 18567 2641
rect 18509 2601 18521 2635
rect 18555 2601 18567 2635
rect 18509 2595 18567 2601
rect 15105 2567 15163 2573
rect 15105 2564 15117 2567
rect 14884 2536 15117 2564
rect 14884 2524 14890 2536
rect 15105 2533 15117 2536
rect 15151 2533 15163 2567
rect 15105 2527 15163 2533
rect 15473 2567 15531 2573
rect 15473 2533 15485 2567
rect 15519 2533 15531 2567
rect 15473 2527 15531 2533
rect 15562 2524 15568 2576
rect 15620 2564 15626 2576
rect 16209 2567 16267 2573
rect 16209 2564 16221 2567
rect 15620 2536 16221 2564
rect 15620 2524 15626 2536
rect 16209 2533 16221 2536
rect 16255 2533 16267 2567
rect 16209 2527 16267 2533
rect 16574 2524 16580 2576
rect 16632 2564 16638 2576
rect 16632 2536 16677 2564
rect 16632 2524 16638 2536
rect 16758 2524 16764 2576
rect 16816 2564 16822 2576
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 16816 2536 16865 2564
rect 16816 2524 16822 2536
rect 16853 2533 16865 2536
rect 16899 2533 16911 2567
rect 17402 2564 17408 2576
rect 17363 2536 17408 2564
rect 16853 2527 16911 2533
rect 17402 2524 17408 2536
rect 17460 2524 17466 2576
rect 17770 2524 17776 2576
rect 17828 2564 17834 2576
rect 18141 2567 18199 2573
rect 18141 2564 18153 2567
rect 17828 2536 18153 2564
rect 17828 2524 17834 2536
rect 18141 2533 18153 2536
rect 18187 2533 18199 2567
rect 18524 2564 18552 2595
rect 18598 2592 18604 2644
rect 18656 2632 18662 2644
rect 19058 2632 19064 2644
rect 18656 2604 18701 2632
rect 19019 2604 19064 2632
rect 18656 2592 18662 2604
rect 19058 2592 19064 2604
rect 19116 2592 19122 2644
rect 19334 2592 19340 2644
rect 19392 2632 19398 2644
rect 19981 2635 20039 2641
rect 19981 2632 19993 2635
rect 19392 2604 19993 2632
rect 19392 2592 19398 2604
rect 19981 2601 19993 2604
rect 20027 2601 20039 2635
rect 19981 2595 20039 2601
rect 20346 2592 20352 2644
rect 20404 2632 20410 2644
rect 21361 2635 21419 2641
rect 21361 2632 21373 2635
rect 20404 2604 21373 2632
rect 20404 2592 20410 2604
rect 21361 2601 21373 2604
rect 21407 2601 21419 2635
rect 21361 2595 21419 2601
rect 18969 2567 19027 2573
rect 18969 2564 18981 2567
rect 18524 2536 18981 2564
rect 18141 2527 18199 2533
rect 18969 2533 18981 2536
rect 19015 2533 19027 2567
rect 18969 2527 19027 2533
rect 19426 2524 19432 2576
rect 19484 2564 19490 2576
rect 20441 2567 20499 2573
rect 20441 2564 20453 2567
rect 19484 2536 20453 2564
rect 19484 2524 19490 2536
rect 20441 2533 20453 2536
rect 20487 2533 20499 2567
rect 20806 2564 20812 2576
rect 20767 2536 20812 2564
rect 20441 2527 20499 2533
rect 20806 2524 20812 2536
rect 20864 2524 20870 2576
rect 20990 2524 20996 2576
rect 21048 2564 21054 2576
rect 21177 2567 21235 2573
rect 21177 2564 21189 2567
rect 21048 2536 21189 2564
rect 21048 2524 21054 2536
rect 21177 2533 21189 2536
rect 21223 2533 21235 2567
rect 21177 2527 21235 2533
rect 14553 2499 14611 2505
rect 14553 2496 14565 2499
rect 14292 2468 14565 2496
rect 14553 2465 14565 2468
rect 14599 2465 14611 2499
rect 14553 2459 14611 2465
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 15252 2468 15853 2496
rect 15252 2456 15258 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 18230 2496 18236 2508
rect 15841 2459 15899 2465
rect 17972 2468 18236 2496
rect 12437 2391 12495 2397
rect 12636 2400 13400 2428
rect 10781 2363 10839 2369
rect 10781 2360 10793 2363
rect 9456 2332 10793 2360
rect 9456 2320 9462 2332
rect 10781 2329 10793 2332
rect 10827 2329 10839 2363
rect 10781 2323 10839 2329
rect 11701 2363 11759 2369
rect 11701 2329 11713 2363
rect 11747 2360 11759 2363
rect 12066 2360 12072 2372
rect 11747 2332 12072 2360
rect 11747 2329 11759 2332
rect 11701 2323 11759 2329
rect 12066 2320 12072 2332
rect 12124 2320 12130 2372
rect 5123 2264 7604 2292
rect 5123 2261 5135 2264
rect 5077 2255 5135 2261
rect 8478 2252 8484 2304
rect 8536 2292 8542 2304
rect 8941 2295 8999 2301
rect 8941 2292 8953 2295
rect 8536 2264 8953 2292
rect 8536 2252 8542 2264
rect 8941 2261 8953 2264
rect 8987 2292 8999 2295
rect 9030 2292 9036 2304
rect 8987 2264 9036 2292
rect 8987 2261 8999 2264
rect 8941 2255 8999 2261
rect 9030 2252 9036 2264
rect 9088 2252 9094 2304
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 12636 2292 12664 2400
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 13596 2400 14933 2428
rect 13596 2388 13602 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 15286 2388 15292 2440
rect 15344 2428 15350 2440
rect 16393 2431 16451 2437
rect 16393 2428 16405 2431
rect 15344 2400 16405 2428
rect 15344 2388 15350 2400
rect 16393 2397 16405 2400
rect 16439 2397 16451 2431
rect 16393 2391 16451 2397
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2428 17095 2431
rect 17310 2428 17316 2440
rect 17083 2400 17316 2428
rect 17083 2397 17095 2400
rect 17037 2391 17095 2397
rect 17310 2388 17316 2400
rect 17368 2388 17374 2440
rect 17972 2437 18000 2468
rect 18230 2456 18236 2468
rect 18288 2456 18294 2508
rect 19613 2499 19671 2505
rect 19613 2496 19625 2499
rect 18708 2468 19625 2496
rect 17957 2431 18015 2437
rect 17957 2397 17969 2431
rect 18003 2397 18015 2431
rect 17957 2391 18015 2397
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18708 2428 18736 2468
rect 19613 2465 19625 2468
rect 19659 2465 19671 2499
rect 19613 2459 19671 2465
rect 19702 2456 19708 2508
rect 19760 2496 19766 2508
rect 20073 2499 20131 2505
rect 20073 2496 20085 2499
rect 19760 2468 20085 2496
rect 19760 2456 19766 2468
rect 20073 2465 20085 2468
rect 20119 2465 20131 2499
rect 20073 2459 20131 2465
rect 21545 2499 21603 2505
rect 21545 2465 21557 2499
rect 21591 2465 21603 2499
rect 21545 2459 21603 2465
rect 18104 2400 18736 2428
rect 18104 2388 18110 2400
rect 18874 2388 18880 2440
rect 18932 2428 18938 2440
rect 19153 2431 19211 2437
rect 19153 2428 19165 2431
rect 18932 2400 19165 2428
rect 18932 2388 18938 2400
rect 19153 2397 19165 2400
rect 19199 2397 19211 2431
rect 19153 2391 19211 2397
rect 19242 2388 19248 2440
rect 19300 2428 19306 2440
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 19300 2400 20637 2428
rect 19300 2388 19306 2400
rect 20625 2397 20637 2400
rect 20671 2397 20683 2431
rect 20625 2391 20683 2397
rect 21082 2388 21088 2440
rect 21140 2428 21146 2440
rect 21560 2428 21588 2459
rect 21140 2400 21588 2428
rect 21140 2388 21146 2400
rect 12710 2320 12716 2372
rect 12768 2360 12774 2372
rect 13817 2363 13875 2369
rect 13817 2360 13829 2363
rect 12768 2332 13829 2360
rect 12768 2320 12774 2332
rect 13817 2329 13829 2332
rect 13863 2329 13875 2363
rect 13817 2323 13875 2329
rect 14826 2320 14832 2372
rect 14884 2360 14890 2372
rect 16025 2363 16083 2369
rect 16025 2360 16037 2363
rect 14884 2332 16037 2360
rect 14884 2320 14890 2332
rect 16025 2329 16037 2332
rect 16071 2329 16083 2363
rect 16025 2323 16083 2329
rect 16850 2320 16856 2372
rect 16908 2360 16914 2372
rect 17221 2363 17279 2369
rect 17221 2360 17233 2363
rect 16908 2332 17233 2360
rect 16908 2320 16914 2332
rect 17221 2329 17233 2332
rect 17267 2329 17279 2363
rect 17221 2323 17279 2329
rect 17678 2320 17684 2372
rect 17736 2360 17742 2372
rect 19429 2363 19487 2369
rect 19429 2360 19441 2363
rect 17736 2332 19441 2360
rect 17736 2320 17742 2332
rect 19429 2329 19441 2332
rect 19475 2329 19487 2363
rect 20257 2363 20315 2369
rect 20257 2360 20269 2363
rect 19429 2323 19487 2329
rect 19536 2332 20269 2360
rect 11940 2264 12664 2292
rect 13541 2295 13599 2301
rect 11940 2252 11946 2264
rect 13541 2261 13553 2295
rect 13587 2292 13599 2295
rect 14366 2292 14372 2304
rect 13587 2264 14372 2292
rect 13587 2261 13599 2264
rect 13541 2255 13599 2261
rect 14366 2252 14372 2264
rect 14424 2252 14430 2304
rect 15378 2292 15384 2304
rect 15339 2264 15384 2292
rect 15378 2252 15384 2264
rect 15436 2252 15442 2304
rect 15746 2292 15752 2304
rect 15707 2264 15752 2292
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 18598 2252 18604 2304
rect 18656 2292 18662 2304
rect 19536 2292 19564 2332
rect 20257 2329 20269 2332
rect 20303 2329 20315 2363
rect 20257 2323 20315 2329
rect 18656 2264 19564 2292
rect 18656 2252 18662 2264
rect 19610 2252 19616 2304
rect 19668 2292 19674 2304
rect 21085 2295 21143 2301
rect 21085 2292 21097 2295
rect 19668 2264 21097 2292
rect 19668 2252 19674 2264
rect 21085 2261 21097 2264
rect 21131 2261 21143 2295
rect 21085 2255 21143 2261
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 1578 2048 1584 2100
rect 1636 2088 1642 2100
rect 1636 2060 5948 2088
rect 1636 2048 1642 2060
rect 5920 1952 5948 2060
rect 5994 2048 6000 2100
rect 6052 2088 6058 2100
rect 11790 2088 11796 2100
rect 6052 2060 11796 2088
rect 6052 2048 6058 2060
rect 11790 2048 11796 2060
rect 11848 2048 11854 2100
rect 6086 1980 6092 2032
rect 6144 2020 6150 2032
rect 6454 2020 6460 2032
rect 6144 1992 6460 2020
rect 6144 1980 6150 1992
rect 6454 1980 6460 1992
rect 6512 2020 6518 2032
rect 10502 2020 10508 2032
rect 6512 1992 10508 2020
rect 6512 1980 6518 1992
rect 10502 1980 10508 1992
rect 10560 1980 10566 2032
rect 11422 1980 11428 2032
rect 11480 2020 11486 2032
rect 13262 2020 13268 2032
rect 11480 1992 13268 2020
rect 11480 1980 11486 1992
rect 13262 1980 13268 1992
rect 13320 1980 13326 2032
rect 5920 1924 6776 1952
rect 2038 1844 2044 1896
rect 2096 1884 2102 1896
rect 6641 1887 6699 1893
rect 6641 1884 6653 1887
rect 2096 1856 6653 1884
rect 2096 1844 2102 1856
rect 6641 1853 6653 1856
rect 6687 1853 6699 1887
rect 6641 1847 6699 1853
rect 3050 1776 3056 1828
rect 3108 1816 3114 1828
rect 4890 1816 4896 1828
rect 3108 1788 4896 1816
rect 3108 1776 3114 1788
rect 4890 1776 4896 1788
rect 4948 1776 4954 1828
rect 5994 1776 6000 1828
rect 6052 1816 6058 1828
rect 6546 1816 6552 1828
rect 6052 1788 6552 1816
rect 6052 1776 6058 1788
rect 6546 1776 6552 1788
rect 6604 1776 6610 1828
rect 6748 1816 6776 1924
rect 8662 1912 8668 1964
rect 8720 1952 8726 1964
rect 9858 1952 9864 1964
rect 8720 1924 9864 1952
rect 8720 1912 8726 1924
rect 9858 1912 9864 1924
rect 9916 1912 9922 1964
rect 6825 1887 6883 1893
rect 6825 1853 6837 1887
rect 6871 1884 6883 1887
rect 8846 1884 8852 1896
rect 6871 1856 8852 1884
rect 6871 1853 6883 1856
rect 6825 1847 6883 1853
rect 8846 1844 8852 1856
rect 8904 1844 8910 1896
rect 10134 1816 10140 1828
rect 6748 1788 10140 1816
rect 10134 1776 10140 1788
rect 10192 1776 10198 1828
rect 2130 1708 2136 1760
rect 2188 1748 2194 1760
rect 2188 1720 2774 1748
rect 2188 1708 2194 1720
rect 2746 1680 2774 1720
rect 6454 1708 6460 1760
rect 6512 1748 6518 1760
rect 7190 1748 7196 1760
rect 6512 1720 7196 1748
rect 6512 1708 6518 1720
rect 7190 1708 7196 1720
rect 7248 1708 7254 1760
rect 9674 1680 9680 1692
rect 2746 1652 9680 1680
rect 9674 1640 9680 1652
rect 9732 1640 9738 1692
rect 9582 1572 9588 1624
rect 9640 1612 9646 1624
rect 11238 1612 11244 1624
rect 9640 1584 11244 1612
rect 9640 1572 9646 1584
rect 11238 1572 11244 1584
rect 11296 1572 11302 1624
rect 14366 1436 14372 1488
rect 14424 1476 14430 1488
rect 15746 1476 15752 1488
rect 14424 1448 15752 1476
rect 14424 1436 14430 1448
rect 15746 1436 15752 1448
rect 15804 1436 15810 1488
rect 13998 1368 14004 1420
rect 14056 1408 14062 1420
rect 15378 1408 15384 1420
rect 14056 1380 15384 1408
rect 14056 1368 14062 1380
rect 15378 1368 15384 1380
rect 15436 1368 15442 1420
<< via1 >>
rect 2872 21904 2924 21956
rect 3148 21904 3200 21956
rect 7104 20748 7156 20800
rect 8852 20748 8904 20800
rect 18052 20748 18104 20800
rect 19340 20748 19392 20800
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 1860 20587 1912 20596
rect 1860 20553 1869 20587
rect 1869 20553 1903 20587
rect 1903 20553 1912 20587
rect 1860 20544 1912 20553
rect 2228 20587 2280 20596
rect 2228 20553 2237 20587
rect 2237 20553 2271 20587
rect 2271 20553 2280 20587
rect 2228 20544 2280 20553
rect 2780 20544 2832 20596
rect 2872 20519 2924 20528
rect 2872 20485 2881 20519
rect 2881 20485 2915 20519
rect 2915 20485 2924 20519
rect 2872 20476 2924 20485
rect 940 20408 992 20460
rect 2688 20408 2740 20460
rect 572 20340 624 20392
rect 2412 20340 2464 20392
rect 5080 20476 5132 20528
rect 5264 20476 5316 20528
rect 9864 20544 9916 20596
rect 18144 20544 18196 20596
rect 21640 20544 21692 20596
rect 4436 20408 4488 20460
rect 3240 20340 3292 20392
rect 3700 20340 3752 20392
rect 1584 20315 1636 20324
rect 1584 20281 1593 20315
rect 1593 20281 1627 20315
rect 1627 20281 1636 20315
rect 1584 20272 1636 20281
rect 2136 20272 2188 20324
rect 2320 20315 2372 20324
rect 2320 20281 2329 20315
rect 2329 20281 2363 20315
rect 2363 20281 2372 20315
rect 2320 20272 2372 20281
rect 2596 20272 2648 20324
rect 9036 20476 9088 20528
rect 10692 20476 10744 20528
rect 10876 20519 10928 20528
rect 10876 20485 10885 20519
rect 10885 20485 10919 20519
rect 10919 20485 10928 20519
rect 10876 20476 10928 20485
rect 11244 20519 11296 20528
rect 11244 20485 11253 20519
rect 11253 20485 11287 20519
rect 11287 20485 11296 20519
rect 11244 20476 11296 20485
rect 11704 20476 11756 20528
rect 12072 20476 12124 20528
rect 12440 20476 12492 20528
rect 12808 20476 12860 20528
rect 13176 20476 13228 20528
rect 13544 20476 13596 20528
rect 14004 20476 14056 20528
rect 14740 20519 14792 20528
rect 14740 20485 14749 20519
rect 14749 20485 14783 20519
rect 14783 20485 14792 20519
rect 14740 20476 14792 20485
rect 15108 20519 15160 20528
rect 15108 20485 15117 20519
rect 15117 20485 15151 20519
rect 15151 20485 15160 20519
rect 15108 20476 15160 20485
rect 15476 20519 15528 20528
rect 15476 20485 15485 20519
rect 15485 20485 15519 20519
rect 15519 20485 15528 20519
rect 15476 20476 15528 20485
rect 15844 20519 15896 20528
rect 15844 20485 15853 20519
rect 15853 20485 15887 20519
rect 15887 20485 15896 20519
rect 15844 20476 15896 20485
rect 16304 20519 16356 20528
rect 16304 20485 16313 20519
rect 16313 20485 16347 20519
rect 16347 20485 16356 20519
rect 16304 20476 16356 20485
rect 16672 20519 16724 20528
rect 16672 20485 16681 20519
rect 16681 20485 16715 20519
rect 16715 20485 16724 20519
rect 16672 20476 16724 20485
rect 17040 20476 17092 20528
rect 17408 20476 17460 20528
rect 17960 20519 18012 20528
rect 17960 20485 17969 20519
rect 17969 20485 18003 20519
rect 18003 20485 18012 20519
rect 17960 20476 18012 20485
rect 18604 20519 18656 20528
rect 18604 20485 18613 20519
rect 18613 20485 18647 20519
rect 18647 20485 18656 20519
rect 18604 20476 18656 20485
rect 20444 20519 20496 20528
rect 20444 20485 20453 20519
rect 20453 20485 20487 20519
rect 20487 20485 20496 20519
rect 20444 20476 20496 20485
rect 20536 20476 20588 20528
rect 20812 20519 20864 20528
rect 20812 20485 20821 20519
rect 20821 20485 20855 20519
rect 20855 20485 20864 20519
rect 20812 20476 20864 20485
rect 4804 20340 4856 20392
rect 5172 20340 5224 20392
rect 5632 20340 5684 20392
rect 6000 20340 6052 20392
rect 6276 20340 6328 20392
rect 6368 20383 6420 20392
rect 6368 20349 6377 20383
rect 6377 20349 6411 20383
rect 6411 20349 6420 20383
rect 6368 20340 6420 20349
rect 1492 20247 1544 20256
rect 1492 20213 1501 20247
rect 1501 20213 1535 20247
rect 1535 20213 1544 20247
rect 1492 20204 1544 20213
rect 2504 20204 2556 20256
rect 3332 20204 3384 20256
rect 3976 20204 4028 20256
rect 4712 20204 4764 20256
rect 4896 20204 4948 20256
rect 5448 20272 5500 20324
rect 6736 20272 6788 20324
rect 7104 20340 7156 20392
rect 7840 20340 7892 20392
rect 8116 20340 8168 20392
rect 8300 20340 8352 20392
rect 8760 20383 8812 20392
rect 8760 20349 8769 20383
rect 8769 20349 8803 20383
rect 8803 20349 8812 20383
rect 8760 20340 8812 20349
rect 9404 20340 9456 20392
rect 9772 20340 9824 20392
rect 10140 20340 10192 20392
rect 10692 20383 10744 20392
rect 10692 20349 10701 20383
rect 10701 20349 10735 20383
rect 10735 20349 10744 20383
rect 10692 20340 10744 20349
rect 7288 20272 7340 20324
rect 8852 20272 8904 20324
rect 9680 20272 9732 20324
rect 6092 20204 6144 20256
rect 7196 20204 7248 20256
rect 7748 20204 7800 20256
rect 8484 20204 8536 20256
rect 8668 20247 8720 20256
rect 8668 20213 8677 20247
rect 8677 20213 8711 20247
rect 8711 20213 8720 20247
rect 8668 20204 8720 20213
rect 9496 20247 9548 20256
rect 9496 20213 9505 20247
rect 9505 20213 9539 20247
rect 9539 20213 9548 20247
rect 9496 20204 9548 20213
rect 9956 20204 10008 20256
rect 10784 20204 10836 20256
rect 18144 20408 18196 20460
rect 19708 20408 19760 20460
rect 17868 20340 17920 20392
rect 18972 20340 19024 20392
rect 19156 20383 19208 20392
rect 19156 20349 19165 20383
rect 19165 20349 19199 20383
rect 19199 20349 19208 20383
rect 19156 20340 19208 20349
rect 19340 20340 19392 20392
rect 20260 20383 20312 20392
rect 20260 20349 20269 20383
rect 20269 20349 20303 20383
rect 20303 20349 20312 20383
rect 20260 20340 20312 20349
rect 21180 20451 21232 20460
rect 21180 20417 21189 20451
rect 21189 20417 21223 20451
rect 21223 20417 21232 20451
rect 21180 20408 21232 20417
rect 20996 20383 21048 20392
rect 20996 20349 21005 20383
rect 21005 20349 21039 20383
rect 21039 20349 21048 20383
rect 20996 20340 21048 20349
rect 11060 20315 11112 20324
rect 11060 20281 11069 20315
rect 11069 20281 11103 20315
rect 11103 20281 11112 20315
rect 11060 20272 11112 20281
rect 11428 20315 11480 20324
rect 11428 20281 11437 20315
rect 11437 20281 11471 20315
rect 11471 20281 11480 20315
rect 11428 20272 11480 20281
rect 12072 20315 12124 20324
rect 12072 20281 12081 20315
rect 12081 20281 12115 20315
rect 12115 20281 12124 20315
rect 12072 20272 12124 20281
rect 12440 20315 12492 20324
rect 12440 20281 12449 20315
rect 12449 20281 12483 20315
rect 12483 20281 12492 20315
rect 12808 20315 12860 20324
rect 12440 20272 12492 20281
rect 12808 20281 12817 20315
rect 12817 20281 12851 20315
rect 12851 20281 12860 20315
rect 12808 20272 12860 20281
rect 13176 20315 13228 20324
rect 13176 20281 13185 20315
rect 13185 20281 13219 20315
rect 13219 20281 13228 20315
rect 13176 20272 13228 20281
rect 13544 20315 13596 20324
rect 13544 20281 13553 20315
rect 13553 20281 13587 20315
rect 13587 20281 13596 20315
rect 13544 20272 13596 20281
rect 13820 20272 13872 20324
rect 14280 20315 14332 20324
rect 14280 20281 14289 20315
rect 14289 20281 14323 20315
rect 14323 20281 14332 20315
rect 14280 20272 14332 20281
rect 14648 20272 14700 20324
rect 15200 20272 15252 20324
rect 15660 20315 15712 20324
rect 15660 20281 15669 20315
rect 15669 20281 15703 20315
rect 15703 20281 15712 20315
rect 15660 20272 15712 20281
rect 16028 20315 16080 20324
rect 16028 20281 16037 20315
rect 16037 20281 16071 20315
rect 16071 20281 16080 20315
rect 16028 20272 16080 20281
rect 16488 20315 16540 20324
rect 16488 20281 16497 20315
rect 16497 20281 16531 20315
rect 16531 20281 16540 20315
rect 16488 20272 16540 20281
rect 16856 20315 16908 20324
rect 16856 20281 16865 20315
rect 16865 20281 16899 20315
rect 16899 20281 16908 20315
rect 16856 20272 16908 20281
rect 17408 20315 17460 20324
rect 17408 20281 17417 20315
rect 17417 20281 17451 20315
rect 17451 20281 17460 20315
rect 17408 20272 17460 20281
rect 17776 20315 17828 20324
rect 17776 20281 17785 20315
rect 17785 20281 17819 20315
rect 17819 20281 17828 20315
rect 17776 20272 17828 20281
rect 17960 20272 18012 20324
rect 15936 20204 15988 20256
rect 17224 20204 17276 20256
rect 18512 20247 18564 20256
rect 18512 20213 18521 20247
rect 18521 20213 18555 20247
rect 18555 20213 18564 20247
rect 18512 20204 18564 20213
rect 18880 20272 18932 20324
rect 19524 20315 19576 20324
rect 19524 20281 19533 20315
rect 19533 20281 19567 20315
rect 19567 20281 19576 20315
rect 19524 20272 19576 20281
rect 22376 20340 22428 20392
rect 21548 20315 21600 20324
rect 20076 20247 20128 20256
rect 20076 20213 20085 20247
rect 20085 20213 20119 20247
rect 20119 20213 20128 20247
rect 20076 20204 20128 20213
rect 20168 20204 20220 20256
rect 21548 20281 21557 20315
rect 21557 20281 21591 20315
rect 21591 20281 21600 20315
rect 21548 20272 21600 20281
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 1400 20000 1452 20052
rect 2044 20000 2096 20052
rect 3056 20000 3108 20052
rect 3240 20000 3292 20052
rect 5448 20000 5500 20052
rect 7012 20000 7064 20052
rect 7288 20000 7340 20052
rect 8760 20000 8812 20052
rect 9404 20000 9456 20052
rect 11428 20000 11480 20052
rect 12808 20000 12860 20052
rect 16948 20043 17000 20052
rect 16948 20009 16957 20043
rect 16957 20009 16991 20043
rect 16991 20009 17000 20043
rect 16948 20000 17000 20009
rect 17224 20043 17276 20052
rect 17224 20009 17233 20043
rect 17233 20009 17267 20043
rect 17267 20009 17276 20043
rect 17224 20000 17276 20009
rect 2228 19932 2280 19984
rect 2044 19864 2096 19916
rect 2412 19907 2464 19916
rect 204 19796 256 19848
rect 1768 19796 1820 19848
rect 2412 19873 2421 19907
rect 2421 19873 2455 19907
rect 2455 19873 2464 19907
rect 2412 19864 2464 19873
rect 3884 19932 3936 19984
rect 3976 19932 4028 19984
rect 2688 19907 2740 19916
rect 2688 19873 2697 19907
rect 2697 19873 2731 19907
rect 2731 19873 2740 19907
rect 2688 19864 2740 19873
rect 3056 19864 3108 19916
rect 3332 19864 3384 19916
rect 3700 19864 3752 19916
rect 4068 19864 4120 19916
rect 5264 19864 5316 19916
rect 5540 19932 5592 19984
rect 6000 19932 6052 19984
rect 6644 19932 6696 19984
rect 7104 19932 7156 19984
rect 7472 19932 7524 19984
rect 6552 19864 6604 19916
rect 6828 19864 6880 19916
rect 8300 19932 8352 19984
rect 5724 19796 5776 19848
rect 7380 19796 7432 19848
rect 9772 19864 9824 19916
rect 10324 19907 10376 19916
rect 10324 19873 10333 19907
rect 10333 19873 10367 19907
rect 10367 19873 10376 19907
rect 10324 19864 10376 19873
rect 10508 19864 10560 19916
rect 14372 19975 14424 19984
rect 14372 19941 14381 19975
rect 14381 19941 14415 19975
rect 14415 19941 14424 19975
rect 14372 19932 14424 19941
rect 11244 19864 11296 19916
rect 12532 19864 12584 19916
rect 14556 19907 14608 19916
rect 14556 19873 14565 19907
rect 14565 19873 14599 19907
rect 14599 19873 14608 19907
rect 14556 19864 14608 19873
rect 17040 19907 17092 19916
rect 17040 19873 17049 19907
rect 17049 19873 17083 19907
rect 17083 19873 17092 19907
rect 17040 19864 17092 19873
rect 17316 19907 17368 19916
rect 17316 19873 17325 19907
rect 17325 19873 17359 19907
rect 17359 19873 17368 19907
rect 17316 19864 17368 19873
rect 8116 19796 8168 19848
rect 17684 19864 17736 19916
rect 17868 19907 17920 19916
rect 17868 19873 17877 19907
rect 17877 19873 17911 19907
rect 17911 19873 17920 19907
rect 17868 19864 17920 19873
rect 18052 19864 18104 19916
rect 4068 19728 4120 19780
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 2872 19703 2924 19712
rect 2872 19669 2881 19703
rect 2881 19669 2915 19703
rect 2915 19669 2924 19703
rect 2872 19660 2924 19669
rect 3240 19660 3292 19712
rect 3424 19703 3476 19712
rect 3424 19669 3433 19703
rect 3433 19669 3467 19703
rect 3467 19669 3476 19703
rect 3424 19660 3476 19669
rect 3792 19660 3844 19712
rect 4988 19660 5040 19712
rect 6184 19660 6236 19712
rect 10140 19728 10192 19780
rect 17500 19771 17552 19780
rect 17500 19737 17509 19771
rect 17509 19737 17543 19771
rect 17543 19737 17552 19771
rect 17500 19728 17552 19737
rect 19248 20000 19300 20052
rect 19064 19932 19116 19984
rect 20076 19975 20128 19984
rect 19432 19864 19484 19916
rect 19708 19907 19760 19916
rect 19708 19873 19717 19907
rect 19717 19873 19751 19907
rect 19751 19873 19760 19907
rect 19708 19864 19760 19873
rect 20076 19941 20085 19975
rect 20085 19941 20119 19975
rect 20119 19941 20128 19975
rect 20076 19932 20128 19941
rect 20444 19975 20496 19984
rect 20444 19941 20453 19975
rect 20453 19941 20487 19975
rect 20487 19941 20496 19975
rect 20444 19932 20496 19941
rect 20720 19932 20772 19984
rect 20996 19864 21048 19916
rect 18696 19796 18748 19848
rect 19064 19796 19116 19848
rect 19892 19839 19944 19848
rect 19892 19805 19901 19839
rect 19901 19805 19935 19839
rect 19935 19805 19944 19839
rect 19892 19796 19944 19805
rect 22008 19932 22060 19984
rect 20536 19728 20588 19780
rect 6920 19660 6972 19712
rect 7288 19660 7340 19712
rect 7656 19703 7708 19712
rect 7656 19669 7665 19703
rect 7665 19669 7699 19703
rect 7699 19669 7708 19703
rect 7656 19660 7708 19669
rect 7748 19660 7800 19712
rect 8300 19660 8352 19712
rect 9404 19660 9456 19712
rect 10232 19660 10284 19712
rect 10692 19660 10744 19712
rect 11796 19703 11848 19712
rect 11796 19669 11805 19703
rect 11805 19669 11839 19703
rect 11839 19669 11848 19703
rect 11796 19660 11848 19669
rect 13636 19660 13688 19712
rect 17868 19660 17920 19712
rect 18604 19660 18656 19712
rect 19340 19660 19392 19712
rect 19800 19660 19852 19712
rect 21456 19703 21508 19712
rect 21456 19669 21465 19703
rect 21465 19669 21499 19703
rect 21499 19669 21508 19703
rect 21456 19660 21508 19669
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 1584 19456 1636 19508
rect 2412 19456 2464 19508
rect 3700 19499 3752 19508
rect 3700 19465 3709 19499
rect 3709 19465 3743 19499
rect 3743 19465 3752 19499
rect 3700 19456 3752 19465
rect 3976 19499 4028 19508
rect 3976 19465 3985 19499
rect 3985 19465 4019 19499
rect 4019 19465 4028 19499
rect 3976 19456 4028 19465
rect 2320 19388 2372 19440
rect 6184 19456 6236 19508
rect 6276 19456 6328 19508
rect 7012 19456 7064 19508
rect 6000 19388 6052 19440
rect 10324 19456 10376 19508
rect 11244 19456 11296 19508
rect 12440 19456 12492 19508
rect 13176 19456 13228 19508
rect 13544 19456 13596 19508
rect 14280 19456 14332 19508
rect 14648 19456 14700 19508
rect 16488 19456 16540 19508
rect 16856 19456 16908 19508
rect 17776 19456 17828 19508
rect 19156 19456 19208 19508
rect 21364 19499 21416 19508
rect 21364 19465 21373 19499
rect 21373 19465 21407 19499
rect 21407 19465 21416 19499
rect 21364 19456 21416 19465
rect 12072 19388 12124 19440
rect 16028 19388 16080 19440
rect 17316 19388 17368 19440
rect 1400 19295 1452 19304
rect 1400 19261 1409 19295
rect 1409 19261 1443 19295
rect 1443 19261 1452 19295
rect 1400 19252 1452 19261
rect 1952 19295 2004 19304
rect 1308 19184 1360 19236
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2688 19320 2740 19372
rect 1860 19184 1912 19236
rect 1676 19116 1728 19168
rect 2504 19252 2556 19304
rect 2780 19295 2832 19304
rect 2780 19261 2789 19295
rect 2789 19261 2823 19295
rect 2823 19261 2832 19295
rect 2780 19252 2832 19261
rect 5632 19320 5684 19372
rect 6552 19320 6604 19372
rect 2412 19116 2464 19168
rect 2688 19184 2740 19236
rect 4896 19252 4948 19304
rect 4988 19252 5040 19304
rect 5448 19252 5500 19304
rect 5724 19252 5776 19304
rect 5908 19295 5960 19304
rect 5908 19261 5917 19295
rect 5917 19261 5951 19295
rect 5951 19261 5960 19295
rect 5908 19252 5960 19261
rect 10600 19320 10652 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 3148 19184 3200 19236
rect 4620 19184 4672 19236
rect 2964 19116 3016 19168
rect 3792 19116 3844 19168
rect 4160 19159 4212 19168
rect 4160 19125 4169 19159
rect 4169 19125 4203 19159
rect 4203 19125 4212 19159
rect 4160 19116 4212 19125
rect 5172 19116 5224 19168
rect 7472 19184 7524 19236
rect 8116 19227 8168 19236
rect 8116 19193 8134 19227
rect 8134 19193 8168 19227
rect 9312 19295 9364 19304
rect 9312 19261 9321 19295
rect 9321 19261 9355 19295
rect 9355 19261 9364 19295
rect 9312 19252 9364 19261
rect 8116 19184 8168 19193
rect 8852 19227 8904 19236
rect 8852 19193 8861 19227
rect 8861 19193 8895 19227
rect 8895 19193 8904 19227
rect 8852 19184 8904 19193
rect 9036 19184 9088 19236
rect 6000 19116 6052 19168
rect 6828 19116 6880 19168
rect 7564 19116 7616 19168
rect 8944 19159 8996 19168
rect 8944 19125 8953 19159
rect 8953 19125 8987 19159
rect 8987 19125 8996 19159
rect 8944 19116 8996 19125
rect 9864 19252 9916 19304
rect 11060 19252 11112 19304
rect 11244 19295 11296 19304
rect 11244 19261 11253 19295
rect 11253 19261 11287 19295
rect 11287 19261 11296 19295
rect 11244 19252 11296 19261
rect 12256 19252 12308 19304
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 13636 19295 13688 19304
rect 11796 19184 11848 19236
rect 12900 19184 12952 19236
rect 13636 19261 13645 19295
rect 13645 19261 13679 19295
rect 13679 19261 13688 19295
rect 13636 19252 13688 19261
rect 14004 19252 14056 19304
rect 14464 19252 14516 19304
rect 10416 19159 10468 19168
rect 10416 19125 10425 19159
rect 10425 19125 10459 19159
rect 10459 19125 10468 19159
rect 10416 19116 10468 19125
rect 10876 19159 10928 19168
rect 10876 19125 10885 19159
rect 10885 19125 10919 19159
rect 10919 19125 10928 19159
rect 10876 19116 10928 19125
rect 11060 19116 11112 19168
rect 12072 19159 12124 19168
rect 12072 19125 12081 19159
rect 12081 19125 12115 19159
rect 12115 19125 12124 19159
rect 12072 19116 12124 19125
rect 12532 19116 12584 19168
rect 13728 19116 13780 19168
rect 17776 19320 17828 19372
rect 18972 19388 19024 19440
rect 19064 19388 19116 19440
rect 20536 19388 20588 19440
rect 15476 19252 15528 19304
rect 16120 19295 16172 19304
rect 16120 19261 16129 19295
rect 16129 19261 16163 19295
rect 16163 19261 16172 19295
rect 16120 19252 16172 19261
rect 17224 19295 17276 19304
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 17224 19252 17276 19261
rect 17500 19252 17552 19304
rect 18052 19184 18104 19236
rect 18788 19252 18840 19304
rect 19156 19252 19208 19304
rect 20720 19252 20772 19304
rect 20904 19252 20956 19304
rect 14464 19116 14516 19168
rect 14740 19159 14792 19168
rect 14740 19125 14749 19159
rect 14749 19125 14783 19159
rect 14783 19125 14792 19159
rect 14740 19116 14792 19125
rect 15200 19116 15252 19168
rect 15936 19159 15988 19168
rect 15936 19125 15945 19159
rect 15945 19125 15979 19159
rect 15979 19125 15988 19159
rect 15936 19116 15988 19125
rect 17040 19159 17092 19168
rect 17040 19125 17049 19159
rect 17049 19125 17083 19159
rect 17083 19125 17092 19159
rect 17040 19116 17092 19125
rect 17592 19116 17644 19168
rect 17960 19116 18012 19168
rect 18696 19159 18748 19168
rect 18696 19125 18705 19159
rect 18705 19125 18739 19159
rect 18739 19125 18748 19159
rect 18696 19116 18748 19125
rect 19248 19184 19300 19236
rect 19892 19116 19944 19168
rect 20076 19116 20128 19168
rect 20720 19116 20772 19168
rect 21088 19116 21140 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 1400 18887 1452 18896
rect 1400 18853 1409 18887
rect 1409 18853 1443 18887
rect 1443 18853 1452 18887
rect 1400 18844 1452 18853
rect 1860 18912 1912 18964
rect 2228 18912 2280 18964
rect 2504 18912 2556 18964
rect 3148 18912 3200 18964
rect 4068 18912 4120 18964
rect 5264 18912 5316 18964
rect 6460 18912 6512 18964
rect 6920 18912 6972 18964
rect 7104 18955 7156 18964
rect 7104 18921 7113 18955
rect 7113 18921 7147 18955
rect 7147 18921 7156 18955
rect 7104 18912 7156 18921
rect 7656 18955 7708 18964
rect 7656 18921 7665 18955
rect 7665 18921 7699 18955
rect 7699 18921 7708 18955
rect 7656 18912 7708 18921
rect 10416 18912 10468 18964
rect 11060 18912 11112 18964
rect 11888 18912 11940 18964
rect 12808 18912 12860 18964
rect 14556 18912 14608 18964
rect 18144 18955 18196 18964
rect 18144 18921 18153 18955
rect 18153 18921 18187 18955
rect 18187 18921 18196 18955
rect 18144 18912 18196 18921
rect 18420 18955 18472 18964
rect 18420 18921 18429 18955
rect 18429 18921 18463 18955
rect 18463 18921 18472 18955
rect 18420 18912 18472 18921
rect 19248 18955 19300 18964
rect 19248 18921 19257 18955
rect 19257 18921 19291 18955
rect 19291 18921 19300 18955
rect 19248 18912 19300 18921
rect 19708 18955 19760 18964
rect 19708 18921 19717 18955
rect 19717 18921 19751 18955
rect 19751 18921 19760 18955
rect 19708 18912 19760 18921
rect 19984 18912 20036 18964
rect 20444 18912 20496 18964
rect 22744 18912 22796 18964
rect 3332 18887 3384 18896
rect 3332 18853 3341 18887
rect 3341 18853 3375 18887
rect 3375 18853 3384 18887
rect 3332 18844 3384 18853
rect 3884 18844 3936 18896
rect 5632 18844 5684 18896
rect 1768 18776 1820 18828
rect 1952 18819 2004 18828
rect 1952 18785 1961 18819
rect 1961 18785 1995 18819
rect 1995 18785 2004 18819
rect 1952 18776 2004 18785
rect 2504 18819 2556 18828
rect 2504 18785 2513 18819
rect 2513 18785 2547 18819
rect 2547 18785 2556 18819
rect 2504 18776 2556 18785
rect 3056 18776 3108 18828
rect 3976 18776 4028 18828
rect 3516 18708 3568 18760
rect 1308 18572 1360 18624
rect 4252 18708 4304 18760
rect 5448 18776 5500 18828
rect 4436 18683 4488 18692
rect 4436 18649 4445 18683
rect 4445 18649 4479 18683
rect 4479 18649 4488 18683
rect 10968 18844 11020 18896
rect 6184 18776 6236 18828
rect 6460 18819 6512 18828
rect 6460 18785 6478 18819
rect 6478 18785 6512 18819
rect 6460 18776 6512 18785
rect 6644 18776 6696 18828
rect 8208 18776 8260 18828
rect 7564 18751 7616 18760
rect 4436 18640 4488 18649
rect 2688 18572 2740 18624
rect 3884 18572 3936 18624
rect 5724 18572 5776 18624
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 11152 18776 11204 18828
rect 11980 18776 12032 18828
rect 12256 18776 12308 18828
rect 18604 18844 18656 18896
rect 16120 18776 16172 18828
rect 19616 18844 19668 18896
rect 10048 18751 10100 18760
rect 7196 18640 7248 18692
rect 6828 18572 6880 18624
rect 6920 18572 6972 18624
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 9036 18640 9088 18692
rect 11796 18708 11848 18760
rect 17500 18751 17552 18760
rect 17500 18717 17509 18751
rect 17509 18717 17543 18751
rect 17543 18717 17552 18751
rect 17500 18708 17552 18717
rect 18604 18708 18656 18760
rect 9772 18572 9824 18624
rect 12808 18640 12860 18692
rect 14648 18640 14700 18692
rect 17592 18640 17644 18692
rect 18696 18683 18748 18692
rect 18696 18649 18705 18683
rect 18705 18649 18739 18683
rect 18739 18649 18748 18683
rect 18696 18640 18748 18649
rect 18972 18683 19024 18692
rect 18972 18649 18981 18683
rect 18981 18649 19015 18683
rect 19015 18649 19024 18683
rect 18972 18640 19024 18649
rect 19892 18819 19944 18828
rect 19892 18785 19901 18819
rect 19901 18785 19935 18819
rect 19935 18785 19944 18819
rect 19892 18776 19944 18785
rect 19984 18819 20036 18828
rect 19984 18785 19993 18819
rect 19993 18785 20027 18819
rect 20027 18785 20036 18819
rect 20536 18844 20588 18896
rect 21272 18844 21324 18896
rect 19984 18776 20036 18785
rect 20628 18819 20680 18828
rect 20628 18785 20637 18819
rect 20637 18785 20671 18819
rect 20671 18785 20680 18819
rect 20628 18776 20680 18785
rect 20996 18819 21048 18828
rect 20996 18785 21005 18819
rect 21005 18785 21039 18819
rect 21039 18785 21048 18819
rect 20996 18776 21048 18785
rect 21364 18819 21416 18828
rect 21364 18785 21373 18819
rect 21373 18785 21407 18819
rect 21407 18785 21416 18819
rect 21364 18776 21416 18785
rect 21548 18819 21600 18828
rect 21548 18785 21557 18819
rect 21557 18785 21591 18819
rect 21591 18785 21600 18819
rect 21548 18776 21600 18785
rect 19340 18708 19392 18760
rect 20352 18708 20404 18760
rect 12900 18615 12952 18624
rect 12900 18581 12909 18615
rect 12909 18581 12943 18615
rect 12943 18581 12952 18615
rect 12900 18572 12952 18581
rect 16580 18572 16632 18624
rect 17224 18572 17276 18624
rect 17960 18615 18012 18624
rect 17960 18581 17969 18615
rect 17969 18581 18003 18615
rect 18003 18581 18012 18615
rect 17960 18572 18012 18581
rect 19156 18572 19208 18624
rect 19524 18640 19576 18692
rect 19984 18572 20036 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 1860 18411 1912 18420
rect 1860 18377 1869 18411
rect 1869 18377 1903 18411
rect 1903 18377 1912 18411
rect 1860 18368 1912 18377
rect 1952 18368 2004 18420
rect 2872 18368 2924 18420
rect 5172 18368 5224 18420
rect 6460 18368 6512 18420
rect 8208 18411 8260 18420
rect 8208 18377 8217 18411
rect 8217 18377 8251 18411
rect 8251 18377 8260 18411
rect 8208 18368 8260 18377
rect 3240 18232 3292 18284
rect 4160 18300 4212 18352
rect 4344 18232 4396 18284
rect 4988 18232 5040 18284
rect 6644 18232 6696 18284
rect 13820 18368 13872 18420
rect 15660 18368 15712 18420
rect 17408 18368 17460 18420
rect 19340 18411 19392 18420
rect 19340 18377 19349 18411
rect 19349 18377 19383 18411
rect 19383 18377 19392 18411
rect 19340 18368 19392 18377
rect 19616 18411 19668 18420
rect 19616 18377 19625 18411
rect 19625 18377 19659 18411
rect 19659 18377 19668 18411
rect 19616 18368 19668 18377
rect 20168 18368 20220 18420
rect 20628 18368 20680 18420
rect 11152 18300 11204 18352
rect 11704 18300 11756 18352
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 5356 18164 5408 18216
rect 6276 18164 6328 18216
rect 6460 18164 6512 18216
rect 8852 18232 8904 18284
rect 7748 18164 7800 18216
rect 8576 18164 8628 18216
rect 9036 18164 9088 18216
rect 9588 18164 9640 18216
rect 11612 18164 11664 18216
rect 12440 18164 12492 18216
rect 14464 18207 14516 18216
rect 14464 18173 14473 18207
rect 14473 18173 14507 18207
rect 14507 18173 14516 18207
rect 14464 18164 14516 18173
rect 15844 18207 15896 18216
rect 15844 18173 15853 18207
rect 15853 18173 15887 18207
rect 15887 18173 15896 18207
rect 15844 18164 15896 18173
rect 19800 18300 19852 18352
rect 20996 18300 21048 18352
rect 21180 18343 21232 18352
rect 21180 18309 21189 18343
rect 21189 18309 21223 18343
rect 21223 18309 21232 18343
rect 21180 18300 21232 18309
rect 18972 18232 19024 18284
rect 19708 18207 19760 18216
rect 3608 18096 3660 18148
rect 4068 18096 4120 18148
rect 2964 18071 3016 18080
rect 2964 18037 2973 18071
rect 2973 18037 3007 18071
rect 3007 18037 3016 18071
rect 2964 18028 3016 18037
rect 3148 18071 3200 18080
rect 3148 18037 3157 18071
rect 3157 18037 3191 18071
rect 3191 18037 3200 18071
rect 3148 18028 3200 18037
rect 3424 18028 3476 18080
rect 3700 18028 3752 18080
rect 3976 18071 4028 18080
rect 3976 18037 3985 18071
rect 3985 18037 4019 18071
rect 4019 18037 4028 18071
rect 3976 18028 4028 18037
rect 5172 18028 5224 18080
rect 6092 18028 6144 18080
rect 6276 18071 6328 18080
rect 6276 18037 6285 18071
rect 6285 18037 6319 18071
rect 6319 18037 6328 18071
rect 6276 18028 6328 18037
rect 6460 18071 6512 18080
rect 6460 18037 6469 18071
rect 6469 18037 6503 18071
rect 6503 18037 6512 18071
rect 6460 18028 6512 18037
rect 6920 18071 6972 18080
rect 6920 18037 6929 18071
rect 6929 18037 6963 18071
rect 6963 18037 6972 18071
rect 6920 18028 6972 18037
rect 7656 18028 7708 18080
rect 8944 18096 8996 18148
rect 10600 18096 10652 18148
rect 11888 18096 11940 18148
rect 19708 18173 19717 18207
rect 19717 18173 19751 18207
rect 19751 18173 19760 18207
rect 19708 18164 19760 18173
rect 19892 18164 19944 18216
rect 20444 18232 20496 18284
rect 18972 18096 19024 18148
rect 19984 18096 20036 18148
rect 21548 18139 21600 18148
rect 21548 18105 21557 18139
rect 21557 18105 21591 18139
rect 21591 18105 21600 18139
rect 21548 18096 21600 18105
rect 10416 18028 10468 18080
rect 10968 18071 11020 18080
rect 10968 18037 10977 18071
rect 10977 18037 11011 18071
rect 11011 18037 11020 18071
rect 10968 18028 11020 18037
rect 12532 18028 12584 18080
rect 20628 18028 20680 18080
rect 21272 18028 21324 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 3148 17824 3200 17876
rect 4252 17824 4304 17876
rect 3240 17756 3292 17808
rect 3976 17756 4028 17808
rect 4528 17867 4580 17876
rect 4528 17833 4537 17867
rect 4537 17833 4571 17867
rect 4571 17833 4580 17867
rect 4896 17867 4948 17876
rect 4528 17824 4580 17833
rect 4896 17833 4905 17867
rect 4905 17833 4939 17867
rect 4939 17833 4948 17867
rect 4896 17824 4948 17833
rect 5264 17867 5316 17876
rect 5264 17833 5273 17867
rect 5273 17833 5307 17867
rect 5307 17833 5316 17867
rect 5264 17824 5316 17833
rect 6460 17824 6512 17876
rect 6736 17824 6788 17876
rect 6920 17824 6972 17876
rect 7196 17824 7248 17876
rect 7564 17824 7616 17876
rect 7748 17824 7800 17876
rect 8208 17867 8260 17876
rect 8208 17833 8217 17867
rect 8217 17833 8251 17867
rect 8251 17833 8260 17867
rect 8208 17824 8260 17833
rect 9772 17824 9824 17876
rect 10048 17824 10100 17876
rect 10416 17867 10468 17876
rect 10416 17833 10425 17867
rect 10425 17833 10459 17867
rect 10459 17833 10468 17867
rect 10416 17824 10468 17833
rect 10876 17824 10928 17876
rect 5540 17756 5592 17808
rect 6000 17756 6052 17808
rect 8760 17756 8812 17808
rect 11980 17824 12032 17876
rect 12072 17824 12124 17876
rect 14464 17824 14516 17876
rect 19708 17824 19760 17876
rect 20444 17824 20496 17876
rect 20628 17867 20680 17876
rect 20628 17833 20637 17867
rect 20637 17833 20671 17867
rect 20671 17833 20680 17867
rect 20628 17824 20680 17833
rect 1952 17731 2004 17740
rect 1952 17697 1961 17731
rect 1961 17697 1995 17731
rect 1995 17697 2004 17731
rect 1952 17688 2004 17697
rect 4160 17688 4212 17740
rect 6276 17688 6328 17740
rect 9864 17731 9916 17740
rect 2412 17620 2464 17672
rect 1768 17595 1820 17604
rect 1768 17561 1777 17595
rect 1777 17561 1811 17595
rect 1811 17561 1820 17595
rect 1768 17552 1820 17561
rect 2596 17552 2648 17604
rect 3608 17620 3660 17672
rect 4068 17620 4120 17672
rect 4988 17620 5040 17672
rect 5448 17663 5500 17672
rect 5448 17629 5457 17663
rect 5457 17629 5491 17663
rect 5491 17629 5500 17663
rect 5448 17620 5500 17629
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 2228 17484 2280 17536
rect 2320 17484 2372 17536
rect 3700 17484 3752 17536
rect 6000 17620 6052 17672
rect 6184 17663 6236 17672
rect 6184 17629 6193 17663
rect 6193 17629 6227 17663
rect 6227 17629 6236 17663
rect 6184 17620 6236 17629
rect 7564 17663 7616 17672
rect 7564 17629 7573 17663
rect 7573 17629 7607 17663
rect 7607 17629 7616 17663
rect 7564 17620 7616 17629
rect 7748 17620 7800 17672
rect 9864 17697 9873 17731
rect 9873 17697 9907 17731
rect 9907 17697 9916 17731
rect 9864 17688 9916 17697
rect 10324 17731 10376 17740
rect 10324 17697 10333 17731
rect 10333 17697 10367 17731
rect 10367 17697 10376 17731
rect 10324 17688 10376 17697
rect 11980 17731 12032 17740
rect 9772 17620 9824 17672
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 11980 17697 11989 17731
rect 11989 17697 12023 17731
rect 12023 17697 12032 17731
rect 11980 17688 12032 17697
rect 13544 17688 13596 17740
rect 11152 17620 11204 17672
rect 11336 17663 11388 17672
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11704 17663 11756 17672
rect 11336 17620 11388 17629
rect 11704 17629 11713 17663
rect 11713 17629 11747 17663
rect 11747 17629 11756 17663
rect 11704 17620 11756 17629
rect 13084 17663 13136 17672
rect 7196 17484 7248 17536
rect 7380 17484 7432 17536
rect 10784 17552 10836 17604
rect 12348 17552 12400 17604
rect 13084 17629 13093 17663
rect 13093 17629 13127 17663
rect 13127 17629 13136 17663
rect 13084 17620 13136 17629
rect 15292 17688 15344 17740
rect 15568 17731 15620 17740
rect 15568 17697 15577 17731
rect 15577 17697 15611 17731
rect 15611 17697 15620 17731
rect 15568 17688 15620 17697
rect 16396 17731 16448 17740
rect 16396 17697 16405 17731
rect 16405 17697 16439 17731
rect 16439 17697 16448 17731
rect 16396 17688 16448 17697
rect 20168 17731 20220 17740
rect 13452 17552 13504 17604
rect 8576 17484 8628 17536
rect 9220 17484 9272 17536
rect 15752 17620 15804 17672
rect 16764 17620 16816 17672
rect 20168 17697 20177 17731
rect 20177 17697 20211 17731
rect 20211 17697 20220 17731
rect 20168 17688 20220 17697
rect 20536 17688 20588 17740
rect 20904 17688 20956 17740
rect 20352 17620 20404 17672
rect 15844 17552 15896 17604
rect 21548 17595 21600 17604
rect 21548 17561 21557 17595
rect 21557 17561 21591 17595
rect 21591 17561 21600 17595
rect 21548 17552 21600 17561
rect 22008 17552 22060 17604
rect 20076 17527 20128 17536
rect 20076 17493 20085 17527
rect 20085 17493 20119 17527
rect 20119 17493 20128 17527
rect 20076 17484 20128 17493
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 3332 17280 3384 17332
rect 4344 17280 4396 17332
rect 5448 17280 5500 17332
rect 2596 17255 2648 17264
rect 2596 17221 2605 17255
rect 2605 17221 2639 17255
rect 2639 17221 2648 17255
rect 2596 17212 2648 17221
rect 4160 17255 4212 17264
rect 4160 17221 4169 17255
rect 4169 17221 4203 17255
rect 4203 17221 4212 17255
rect 4160 17212 4212 17221
rect 7380 17280 7432 17332
rect 7656 17280 7708 17332
rect 1768 17008 1820 17060
rect 2320 17144 2372 17196
rect 3792 17144 3844 17196
rect 5724 17212 5776 17264
rect 8392 17212 8444 17264
rect 4988 17144 5040 17196
rect 5816 17144 5868 17196
rect 6184 17144 6236 17196
rect 7564 17144 7616 17196
rect 9036 17280 9088 17332
rect 11980 17280 12032 17332
rect 13452 17280 13504 17332
rect 16764 17323 16816 17332
rect 16764 17289 16773 17323
rect 16773 17289 16807 17323
rect 16807 17289 16816 17323
rect 16764 17280 16816 17289
rect 21364 17280 21416 17332
rect 10048 17144 10100 17196
rect 11152 17212 11204 17264
rect 12348 17212 12400 17264
rect 21640 17212 21692 17264
rect 10600 17187 10652 17196
rect 10600 17153 10609 17187
rect 10609 17153 10643 17187
rect 10643 17153 10652 17187
rect 10600 17144 10652 17153
rect 11796 17144 11848 17196
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12440 17144 12492 17153
rect 13452 17144 13504 17196
rect 2228 17119 2280 17128
rect 2228 17085 2237 17119
rect 2237 17085 2271 17119
rect 2271 17085 2280 17119
rect 2228 17076 2280 17085
rect 5632 17076 5684 17128
rect 6552 17076 6604 17128
rect 8576 17076 8628 17128
rect 8852 17076 8904 17128
rect 9588 17076 9640 17128
rect 10968 17076 11020 17128
rect 11704 17076 11756 17128
rect 13912 17119 13964 17128
rect 13912 17085 13921 17119
rect 13921 17085 13955 17119
rect 13955 17085 13964 17119
rect 13912 17076 13964 17085
rect 20904 17144 20956 17196
rect 21548 17187 21600 17196
rect 21548 17153 21557 17187
rect 21557 17153 21591 17187
rect 21591 17153 21600 17187
rect 21548 17144 21600 17153
rect 17408 17076 17460 17128
rect 19892 17076 19944 17128
rect 20812 17119 20864 17128
rect 20812 17085 20821 17119
rect 20821 17085 20855 17119
rect 20855 17085 20864 17119
rect 20812 17076 20864 17085
rect 3148 17008 3200 17060
rect 4436 17008 4488 17060
rect 5172 17008 5224 17060
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 5724 16940 5776 16992
rect 6920 17008 6972 17060
rect 11612 17008 11664 17060
rect 11888 17008 11940 17060
rect 13268 17008 13320 17060
rect 13820 17008 13872 17060
rect 8944 16940 8996 16992
rect 9220 16940 9272 16992
rect 9404 16940 9456 16992
rect 10600 16940 10652 16992
rect 10968 16940 11020 16992
rect 15292 16983 15344 16992
rect 15292 16949 15301 16983
rect 15301 16949 15335 16983
rect 15335 16949 15344 16983
rect 15292 16940 15344 16949
rect 15752 17008 15804 17060
rect 21364 17051 21416 17060
rect 21364 17017 21373 17051
rect 21373 17017 21407 17051
rect 21407 17017 21416 17051
rect 21364 17008 21416 17017
rect 20168 16940 20220 16992
rect 20536 16940 20588 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 1768 16779 1820 16788
rect 1768 16745 1777 16779
rect 1777 16745 1811 16779
rect 1811 16745 1820 16779
rect 1768 16736 1820 16745
rect 1952 16736 2004 16788
rect 3240 16668 3292 16720
rect 2320 16600 2372 16652
rect 3424 16643 3476 16652
rect 3424 16609 3433 16643
rect 3433 16609 3467 16643
rect 3467 16609 3476 16643
rect 3424 16600 3476 16609
rect 7288 16736 7340 16788
rect 7564 16736 7616 16788
rect 8576 16736 8628 16788
rect 10508 16736 10560 16788
rect 10784 16736 10836 16788
rect 10968 16736 11020 16788
rect 11612 16736 11664 16788
rect 15752 16779 15804 16788
rect 15752 16745 15761 16779
rect 15761 16745 15795 16779
rect 15795 16745 15804 16779
rect 15752 16736 15804 16745
rect 4344 16711 4396 16720
rect 4344 16677 4378 16711
rect 4378 16677 4396 16711
rect 4344 16668 4396 16677
rect 3148 16575 3200 16584
rect 3148 16541 3157 16575
rect 3157 16541 3191 16575
rect 3191 16541 3200 16575
rect 5632 16600 5684 16652
rect 6000 16668 6052 16720
rect 8392 16668 8444 16720
rect 6184 16600 6236 16652
rect 6276 16600 6328 16652
rect 9588 16668 9640 16720
rect 10416 16668 10468 16720
rect 11704 16668 11756 16720
rect 15292 16668 15344 16720
rect 9864 16600 9916 16652
rect 10324 16600 10376 16652
rect 3148 16532 3200 16541
rect 9036 16532 9088 16584
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 10048 16532 10100 16541
rect 10416 16532 10468 16584
rect 11152 16600 11204 16652
rect 3516 16464 3568 16516
rect 3700 16464 3752 16516
rect 8944 16507 8996 16516
rect 8944 16473 8953 16507
rect 8953 16473 8987 16507
rect 8987 16473 8996 16507
rect 8944 16464 8996 16473
rect 11060 16532 11112 16584
rect 12532 16600 12584 16652
rect 12716 16643 12768 16652
rect 12716 16609 12725 16643
rect 12725 16609 12759 16643
rect 12759 16609 12768 16643
rect 12716 16600 12768 16609
rect 13084 16600 13136 16652
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 12440 16532 12492 16541
rect 13820 16600 13872 16652
rect 13912 16600 13964 16652
rect 20812 16736 20864 16788
rect 16764 16668 16816 16720
rect 19892 16668 19944 16720
rect 17408 16643 17460 16652
rect 13268 16532 13320 16584
rect 14280 16532 14332 16584
rect 17408 16609 17417 16643
rect 17417 16609 17451 16643
rect 17451 16609 17460 16643
rect 17408 16600 17460 16609
rect 19340 16600 19392 16652
rect 21548 16711 21600 16720
rect 21548 16677 21557 16711
rect 21557 16677 21591 16711
rect 21591 16677 21600 16711
rect 21548 16668 21600 16677
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 2412 16396 2464 16448
rect 5264 16396 5316 16448
rect 6184 16396 6236 16448
rect 6920 16439 6972 16448
rect 6920 16405 6929 16439
rect 6929 16405 6963 16439
rect 6963 16405 6972 16439
rect 6920 16396 6972 16405
rect 13728 16396 13780 16448
rect 15384 16396 15436 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 2412 16192 2464 16244
rect 3240 16235 3292 16244
rect 3240 16201 3249 16235
rect 3249 16201 3283 16235
rect 3283 16201 3292 16235
rect 3240 16192 3292 16201
rect 3332 16192 3384 16244
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 2320 16056 2372 16108
rect 9312 16192 9364 16244
rect 9588 16192 9640 16244
rect 10324 16192 10376 16244
rect 12256 16192 12308 16244
rect 13268 16235 13320 16244
rect 13268 16201 13277 16235
rect 13277 16201 13311 16235
rect 13311 16201 13320 16235
rect 13268 16192 13320 16201
rect 13544 16192 13596 16244
rect 15568 16192 15620 16244
rect 21364 16192 21416 16244
rect 5540 16099 5592 16108
rect 5540 16065 5549 16099
rect 5549 16065 5583 16099
rect 5583 16065 5592 16099
rect 5540 16056 5592 16065
rect 6460 16056 6512 16108
rect 6920 16056 6972 16108
rect 8392 16099 8444 16108
rect 8392 16065 8401 16099
rect 8401 16065 8435 16099
rect 8435 16065 8444 16099
rect 8392 16056 8444 16065
rect 9864 16124 9916 16176
rect 21548 16167 21600 16176
rect 11796 16056 11848 16108
rect 21548 16133 21557 16167
rect 21557 16133 21591 16167
rect 21591 16133 21600 16167
rect 21548 16124 21600 16133
rect 2872 15963 2924 15972
rect 2872 15929 2881 15963
rect 2881 15929 2915 15963
rect 2915 15929 2924 15963
rect 2872 15920 2924 15929
rect 5816 15988 5868 16040
rect 3792 15920 3844 15972
rect 4436 15920 4488 15972
rect 5540 15920 5592 15972
rect 6276 15988 6328 16040
rect 9956 15988 10008 16040
rect 10232 15988 10284 16040
rect 6644 15920 6696 15972
rect 7656 15963 7708 15972
rect 7656 15929 7665 15963
rect 7665 15929 7699 15963
rect 7699 15929 7708 15963
rect 7656 15920 7708 15929
rect 2780 15895 2832 15904
rect 2780 15861 2789 15895
rect 2789 15861 2823 15895
rect 2823 15861 2832 15895
rect 4252 15895 4304 15904
rect 2780 15852 2832 15861
rect 4252 15861 4261 15895
rect 4261 15861 4295 15895
rect 4295 15861 4304 15895
rect 4252 15852 4304 15861
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 6000 15895 6052 15904
rect 6000 15861 6009 15895
rect 6009 15861 6043 15895
rect 6043 15861 6052 15895
rect 6000 15852 6052 15861
rect 6276 15852 6328 15904
rect 6920 15895 6972 15904
rect 6920 15861 6929 15895
rect 6929 15861 6963 15895
rect 6963 15861 6972 15895
rect 7748 15895 7800 15904
rect 6920 15852 6972 15861
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 9036 15920 9088 15972
rect 12440 15988 12492 16040
rect 13176 15988 13228 16040
rect 15292 16056 15344 16108
rect 13728 15988 13780 16040
rect 20628 16031 20680 16040
rect 10784 15963 10836 15972
rect 10784 15929 10802 15963
rect 10802 15929 10836 15963
rect 10784 15920 10836 15929
rect 20628 15997 20637 16031
rect 20637 15997 20671 16031
rect 20671 15997 20680 16031
rect 20628 15988 20680 15997
rect 8392 15852 8444 15904
rect 9496 15852 9548 15904
rect 9864 15852 9916 15904
rect 11704 15895 11756 15904
rect 11704 15861 11713 15895
rect 11713 15861 11747 15895
rect 11747 15861 11756 15895
rect 11704 15852 11756 15861
rect 13912 15852 13964 15904
rect 20720 15920 20772 15972
rect 21180 15963 21232 15972
rect 21180 15929 21189 15963
rect 21189 15929 21223 15963
rect 21223 15929 21232 15963
rect 21180 15920 21232 15929
rect 14280 15852 14332 15904
rect 15844 15852 15896 15904
rect 16120 15895 16172 15904
rect 16120 15861 16129 15895
rect 16129 15861 16163 15895
rect 16163 15861 16172 15895
rect 16120 15852 16172 15861
rect 16304 15852 16356 15904
rect 20904 15852 20956 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 1860 15691 1912 15700
rect 1860 15657 1869 15691
rect 1869 15657 1903 15691
rect 1903 15657 1912 15691
rect 1860 15648 1912 15657
rect 2320 15691 2372 15700
rect 2320 15657 2329 15691
rect 2329 15657 2363 15691
rect 2363 15657 2372 15691
rect 2320 15648 2372 15657
rect 3424 15648 3476 15700
rect 4436 15691 4488 15700
rect 4436 15657 4445 15691
rect 4445 15657 4479 15691
rect 4479 15657 4488 15691
rect 4436 15648 4488 15657
rect 6000 15648 6052 15700
rect 6460 15691 6512 15700
rect 6460 15657 6469 15691
rect 6469 15657 6503 15691
rect 6503 15657 6512 15691
rect 6460 15648 6512 15657
rect 7748 15648 7800 15700
rect 8944 15648 8996 15700
rect 11152 15648 11204 15700
rect 11244 15648 11296 15700
rect 11888 15648 11940 15700
rect 12716 15648 12768 15700
rect 13912 15691 13964 15700
rect 13912 15657 13921 15691
rect 13921 15657 13955 15691
rect 13955 15657 13964 15691
rect 13912 15648 13964 15657
rect 14372 15648 14424 15700
rect 16120 15648 16172 15700
rect 3240 15580 3292 15632
rect 5172 15580 5224 15632
rect 5724 15580 5776 15632
rect 6552 15580 6604 15632
rect 1584 15555 1636 15564
rect 1584 15521 1593 15555
rect 1593 15521 1627 15555
rect 1627 15521 1636 15555
rect 1584 15512 1636 15521
rect 1952 15555 2004 15564
rect 1952 15521 1961 15555
rect 1961 15521 1995 15555
rect 1995 15521 2004 15555
rect 1952 15512 2004 15521
rect 4712 15512 4764 15564
rect 5908 15512 5960 15564
rect 9496 15580 9548 15632
rect 3700 15487 3752 15496
rect 3700 15453 3709 15487
rect 3709 15453 3743 15487
rect 3743 15453 3752 15487
rect 3700 15444 3752 15453
rect 4160 15444 4212 15496
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 5632 15444 5684 15496
rect 8576 15512 8628 15564
rect 9036 15512 9088 15564
rect 6184 15487 6236 15496
rect 1400 15419 1452 15428
rect 1400 15385 1409 15419
rect 1409 15385 1443 15419
rect 1443 15385 1452 15419
rect 1400 15376 1452 15385
rect 3792 15376 3844 15428
rect 6184 15453 6193 15487
rect 6193 15453 6227 15487
rect 6227 15453 6236 15487
rect 6184 15444 6236 15453
rect 6736 15444 6788 15496
rect 7196 15487 7248 15496
rect 7196 15453 7205 15487
rect 7205 15453 7239 15487
rect 7239 15453 7248 15487
rect 10232 15512 10284 15564
rect 11152 15512 11204 15564
rect 13268 15512 13320 15564
rect 13452 15555 13504 15564
rect 13452 15521 13461 15555
rect 13461 15521 13495 15555
rect 13495 15521 13504 15555
rect 13452 15512 13504 15521
rect 14096 15512 14148 15564
rect 10784 15487 10836 15496
rect 7196 15444 7248 15453
rect 6276 15376 6328 15428
rect 10784 15453 10793 15487
rect 10793 15453 10827 15487
rect 10827 15453 10836 15487
rect 10784 15444 10836 15453
rect 10876 15487 10928 15496
rect 10876 15453 10885 15487
rect 10885 15453 10919 15487
rect 10919 15453 10928 15487
rect 11980 15487 12032 15496
rect 10876 15444 10928 15453
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 12440 15487 12492 15496
rect 12440 15453 12449 15487
rect 12449 15453 12483 15487
rect 12483 15453 12492 15487
rect 12440 15444 12492 15453
rect 2044 15308 2096 15360
rect 5172 15308 5224 15360
rect 5448 15308 5500 15360
rect 8208 15308 8260 15360
rect 12900 15444 12952 15496
rect 13176 15487 13228 15496
rect 13176 15453 13185 15487
rect 13185 15453 13219 15487
rect 13219 15453 13228 15487
rect 13176 15444 13228 15453
rect 11888 15308 11940 15360
rect 11980 15308 12032 15360
rect 14280 15376 14332 15428
rect 15292 15580 15344 15632
rect 14832 15487 14884 15496
rect 14832 15453 14841 15487
rect 14841 15453 14875 15487
rect 14875 15453 14884 15487
rect 15384 15512 15436 15564
rect 14832 15444 14884 15453
rect 19892 15648 19944 15700
rect 20260 15648 20312 15700
rect 20720 15691 20772 15700
rect 17500 15580 17552 15632
rect 20720 15657 20729 15691
rect 20729 15657 20763 15691
rect 20763 15657 20772 15691
rect 20720 15648 20772 15657
rect 19616 15512 19668 15564
rect 20904 15580 20956 15632
rect 17960 15487 18012 15496
rect 17960 15453 17969 15487
rect 17969 15453 18003 15487
rect 18003 15453 18012 15487
rect 17960 15444 18012 15453
rect 18052 15444 18104 15496
rect 20444 15512 20496 15564
rect 20168 15444 20220 15496
rect 21548 15419 21600 15428
rect 15200 15308 15252 15360
rect 15936 15308 15988 15360
rect 16120 15351 16172 15360
rect 16120 15317 16129 15351
rect 16129 15317 16163 15351
rect 16163 15317 16172 15351
rect 16120 15308 16172 15317
rect 16212 15308 16264 15360
rect 21548 15385 21557 15419
rect 21557 15385 21591 15419
rect 21591 15385 21600 15419
rect 21548 15376 21600 15385
rect 19524 15308 19576 15360
rect 20444 15308 20496 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 1952 15104 2004 15156
rect 2872 15104 2924 15156
rect 4252 15104 4304 15156
rect 5632 15104 5684 15156
rect 6736 15104 6788 15156
rect 1584 15036 1636 15088
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 2044 14900 2096 14952
rect 2228 14943 2280 14952
rect 2228 14909 2237 14943
rect 2237 14909 2271 14943
rect 2271 14909 2280 14943
rect 2228 14900 2280 14909
rect 3976 15036 4028 15088
rect 6552 15036 6604 15088
rect 7196 15104 7248 15156
rect 10876 15104 10928 15156
rect 8208 15036 8260 15088
rect 3240 15011 3292 15020
rect 3240 14977 3249 15011
rect 3249 14977 3283 15011
rect 3283 14977 3292 15011
rect 3240 14968 3292 14977
rect 2504 14764 2556 14816
rect 4160 14900 4212 14952
rect 4988 14900 5040 14952
rect 5540 14900 5592 14952
rect 7748 14968 7800 15020
rect 9496 14968 9548 15020
rect 7012 14900 7064 14952
rect 11060 14968 11112 15020
rect 12348 15104 12400 15156
rect 13820 15104 13872 15156
rect 14096 15104 14148 15156
rect 16212 15104 16264 15156
rect 16396 15147 16448 15156
rect 16396 15113 16405 15147
rect 16405 15113 16439 15147
rect 16439 15113 16448 15147
rect 16396 15104 16448 15113
rect 20168 15147 20220 15156
rect 13084 15036 13136 15088
rect 20168 15113 20177 15147
rect 20177 15113 20211 15147
rect 20211 15113 20220 15147
rect 20168 15104 20220 15113
rect 20628 15104 20680 15156
rect 13176 14968 13228 15020
rect 11336 14900 11388 14952
rect 11796 14900 11848 14952
rect 12440 14900 12492 14952
rect 12992 14900 13044 14952
rect 13544 14968 13596 15020
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 15752 15011 15804 15020
rect 15752 14977 15761 15011
rect 15761 14977 15795 15011
rect 15795 14977 15804 15011
rect 15752 14968 15804 14977
rect 15936 15011 15988 15020
rect 15936 14977 15945 15011
rect 15945 14977 15979 15011
rect 15979 14977 15988 15011
rect 15936 14968 15988 14977
rect 17408 14968 17460 15020
rect 14648 14900 14700 14952
rect 16120 14900 16172 14952
rect 19524 14900 19576 14952
rect 21548 15011 21600 15020
rect 21548 14977 21557 15011
rect 21557 14977 21591 15011
rect 21591 14977 21600 15011
rect 21548 14968 21600 14977
rect 7840 14832 7892 14884
rect 9588 14832 9640 14884
rect 10324 14832 10376 14884
rect 10600 14832 10652 14884
rect 3516 14807 3568 14816
rect 3516 14773 3525 14807
rect 3525 14773 3559 14807
rect 3559 14773 3568 14807
rect 3516 14764 3568 14773
rect 3792 14807 3844 14816
rect 3792 14773 3801 14807
rect 3801 14773 3835 14807
rect 3835 14773 3844 14807
rect 3792 14764 3844 14773
rect 4068 14764 4120 14816
rect 4436 14807 4488 14816
rect 4436 14773 4445 14807
rect 4445 14773 4479 14807
rect 4479 14773 4488 14807
rect 4436 14764 4488 14773
rect 5264 14764 5316 14816
rect 6000 14764 6052 14816
rect 6644 14764 6696 14816
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 7380 14764 7432 14816
rect 8576 14807 8628 14816
rect 8576 14773 8585 14807
rect 8585 14773 8619 14807
rect 8619 14773 8628 14807
rect 8576 14764 8628 14773
rect 9864 14807 9916 14816
rect 9864 14773 9873 14807
rect 9873 14773 9907 14807
rect 9907 14773 9916 14807
rect 9864 14764 9916 14773
rect 10784 14807 10836 14816
rect 10784 14773 10793 14807
rect 10793 14773 10827 14807
rect 10827 14773 10836 14807
rect 10784 14764 10836 14773
rect 11152 14832 11204 14884
rect 12164 14832 12216 14884
rect 14096 14832 14148 14884
rect 14832 14832 14884 14884
rect 16948 14832 17000 14884
rect 17224 14832 17276 14884
rect 12348 14764 12400 14816
rect 13176 14764 13228 14816
rect 13268 14764 13320 14816
rect 13912 14764 13964 14816
rect 14188 14807 14240 14816
rect 14188 14773 14197 14807
rect 14197 14773 14231 14807
rect 14231 14773 14240 14807
rect 14188 14764 14240 14773
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 15936 14764 15988 14816
rect 17960 14764 18012 14816
rect 20812 14764 20864 14816
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 2780 14560 2832 14612
rect 3516 14560 3568 14612
rect 4160 14560 4212 14612
rect 6920 14560 6972 14612
rect 7288 14560 7340 14612
rect 2044 14492 2096 14544
rect 2872 14492 2924 14544
rect 3148 14492 3200 14544
rect 3700 14492 3752 14544
rect 4344 14492 4396 14544
rect 6276 14492 6328 14544
rect 11152 14560 11204 14612
rect 7564 14492 7616 14544
rect 4252 14467 4304 14476
rect 4252 14433 4261 14467
rect 4261 14433 4295 14467
rect 4295 14433 4304 14467
rect 4252 14424 4304 14433
rect 6460 14424 6512 14476
rect 7012 14424 7064 14476
rect 8852 14492 8904 14544
rect 9588 14492 9640 14544
rect 11060 14492 11112 14544
rect 12164 14560 12216 14612
rect 12532 14560 12584 14612
rect 14004 14560 14056 14612
rect 2412 14356 2464 14408
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 3976 14356 4028 14408
rect 4344 14399 4396 14408
rect 4344 14365 4353 14399
rect 4353 14365 4387 14399
rect 4387 14365 4396 14399
rect 4344 14356 4396 14365
rect 5724 14356 5776 14408
rect 6184 14356 6236 14408
rect 7196 14399 7248 14408
rect 7196 14365 7205 14399
rect 7205 14365 7239 14399
rect 7239 14365 7248 14399
rect 7196 14356 7248 14365
rect 2872 14288 2924 14340
rect 4436 14288 4488 14340
rect 5540 14288 5592 14340
rect 6736 14288 6788 14340
rect 7472 14288 7524 14340
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2504 14263 2556 14272
rect 2504 14229 2513 14263
rect 2513 14229 2547 14263
rect 2547 14229 2556 14263
rect 2504 14220 2556 14229
rect 4988 14263 5040 14272
rect 4988 14229 4997 14263
rect 4997 14229 5031 14263
rect 5031 14229 5040 14263
rect 4988 14220 5040 14229
rect 5172 14263 5224 14272
rect 5172 14229 5181 14263
rect 5181 14229 5215 14263
rect 5215 14229 5224 14263
rect 5172 14220 5224 14229
rect 8852 14288 8904 14340
rect 8576 14220 8628 14272
rect 9404 14288 9456 14340
rect 9496 14220 9548 14272
rect 10692 14356 10744 14408
rect 11428 14424 11480 14476
rect 12624 14492 12676 14544
rect 13636 14492 13688 14544
rect 15476 14535 15528 14544
rect 15476 14501 15494 14535
rect 15494 14501 15528 14535
rect 15476 14492 15528 14501
rect 10784 14288 10836 14340
rect 10692 14220 10744 14272
rect 11980 14424 12032 14476
rect 12164 14356 12216 14408
rect 12440 14356 12492 14408
rect 12808 14399 12860 14408
rect 12808 14365 12817 14399
rect 12817 14365 12851 14399
rect 12851 14365 12860 14399
rect 12808 14356 12860 14365
rect 12992 14356 13044 14408
rect 14556 14424 14608 14476
rect 18972 14560 19024 14612
rect 19616 14603 19668 14612
rect 19616 14569 19625 14603
rect 19625 14569 19659 14603
rect 19659 14569 19668 14603
rect 19616 14560 19668 14569
rect 17960 14492 18012 14544
rect 21180 14535 21232 14544
rect 21180 14501 21189 14535
rect 21189 14501 21223 14535
rect 21223 14501 21232 14535
rect 21180 14492 21232 14501
rect 16856 14424 16908 14476
rect 17408 14424 17460 14476
rect 18144 14424 18196 14476
rect 19524 14424 19576 14476
rect 20628 14467 20680 14476
rect 20628 14433 20637 14467
rect 20637 14433 20671 14467
rect 20671 14433 20680 14467
rect 20628 14424 20680 14433
rect 21364 14467 21416 14476
rect 21364 14433 21373 14467
rect 21373 14433 21407 14467
rect 21407 14433 21416 14467
rect 21364 14424 21416 14433
rect 19064 14399 19116 14408
rect 19064 14365 19073 14399
rect 19073 14365 19107 14399
rect 19107 14365 19116 14399
rect 19064 14356 19116 14365
rect 19156 14356 19208 14408
rect 21548 14331 21600 14340
rect 11060 14220 11112 14272
rect 11796 14220 11848 14272
rect 11888 14220 11940 14272
rect 13360 14263 13412 14272
rect 13360 14229 13369 14263
rect 13369 14229 13403 14263
rect 13403 14229 13412 14263
rect 13360 14220 13412 14229
rect 13452 14220 13504 14272
rect 14740 14220 14792 14272
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 17224 14220 17276 14272
rect 21548 14297 21557 14331
rect 21557 14297 21591 14331
rect 21591 14297 21600 14331
rect 21548 14288 21600 14297
rect 20628 14220 20680 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 2228 14016 2280 14068
rect 2964 14016 3016 14068
rect 5816 14016 5868 14068
rect 7656 14016 7708 14068
rect 9864 14016 9916 14068
rect 12532 14059 12584 14068
rect 2412 13991 2464 14000
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 1768 13855 1820 13864
rect 1768 13821 1777 13855
rect 1777 13821 1811 13855
rect 1811 13821 1820 13855
rect 1768 13812 1820 13821
rect 2412 13957 2421 13991
rect 2421 13957 2455 13991
rect 2455 13957 2464 13991
rect 2412 13948 2464 13957
rect 3884 13948 3936 14000
rect 4896 13948 4948 14000
rect 2320 13855 2372 13864
rect 2320 13821 2329 13855
rect 2329 13821 2363 13855
rect 2363 13821 2372 13855
rect 2320 13812 2372 13821
rect 5632 13880 5684 13932
rect 6184 13923 6236 13932
rect 6184 13889 6193 13923
rect 6193 13889 6227 13923
rect 6227 13889 6236 13923
rect 6184 13880 6236 13889
rect 6644 13880 6696 13932
rect 5356 13812 5408 13864
rect 5908 13812 5960 13864
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 9220 13948 9272 14000
rect 12532 14025 12541 14059
rect 12541 14025 12575 14059
rect 12575 14025 12584 14059
rect 12532 14016 12584 14025
rect 13360 14016 13412 14068
rect 16488 14059 16540 14068
rect 10692 13948 10744 14000
rect 9588 13923 9640 13932
rect 9588 13889 9597 13923
rect 9597 13889 9631 13923
rect 9631 13889 9640 13923
rect 9588 13880 9640 13889
rect 11980 13948 12032 14000
rect 13636 13948 13688 14000
rect 11888 13923 11940 13932
rect 11888 13889 11897 13923
rect 11897 13889 11931 13923
rect 11931 13889 11940 13923
rect 11888 13880 11940 13889
rect 13452 13880 13504 13932
rect 16488 14025 16497 14059
rect 16497 14025 16531 14059
rect 16531 14025 16540 14059
rect 16948 14059 17000 14068
rect 16488 14016 16540 14025
rect 16948 14025 16957 14059
rect 16957 14025 16991 14059
rect 16991 14025 17000 14059
rect 16948 14016 17000 14025
rect 19156 14016 19208 14068
rect 19524 14059 19576 14068
rect 19524 14025 19533 14059
rect 19533 14025 19567 14059
rect 19567 14025 19576 14059
rect 19524 14016 19576 14025
rect 21364 14016 21416 14068
rect 16672 13948 16724 14000
rect 18144 13923 18196 13932
rect 18144 13889 18153 13923
rect 18153 13889 18187 13923
rect 18187 13889 18196 13923
rect 18880 13923 18932 13932
rect 18144 13880 18196 13889
rect 18880 13889 18889 13923
rect 18889 13889 18923 13923
rect 18923 13889 18932 13923
rect 18880 13880 18932 13889
rect 7288 13812 7340 13864
rect 7748 13812 7800 13864
rect 2136 13744 2188 13796
rect 3148 13744 3200 13796
rect 2412 13676 2464 13728
rect 3240 13676 3292 13728
rect 4712 13744 4764 13796
rect 9588 13744 9640 13796
rect 10324 13744 10376 13796
rect 11336 13812 11388 13864
rect 13084 13787 13136 13796
rect 13084 13753 13093 13787
rect 13093 13753 13127 13787
rect 13127 13753 13136 13787
rect 13084 13744 13136 13753
rect 5908 13719 5960 13728
rect 5908 13685 5917 13719
rect 5917 13685 5951 13719
rect 5951 13685 5960 13719
rect 5908 13676 5960 13685
rect 7564 13676 7616 13728
rect 8208 13719 8260 13728
rect 8208 13685 8217 13719
rect 8217 13685 8251 13719
rect 8251 13685 8260 13719
rect 8208 13676 8260 13685
rect 9864 13676 9916 13728
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 10416 13676 10468 13728
rect 11980 13719 12032 13728
rect 11980 13685 11989 13719
rect 11989 13685 12023 13719
rect 12023 13685 12032 13719
rect 11980 13676 12032 13685
rect 12164 13676 12216 13728
rect 12808 13676 12860 13728
rect 12992 13719 13044 13728
rect 12992 13685 13001 13719
rect 13001 13685 13035 13719
rect 13035 13685 13044 13719
rect 12992 13676 13044 13685
rect 13544 13812 13596 13864
rect 13820 13812 13872 13864
rect 14372 13812 14424 13864
rect 16856 13812 16908 13864
rect 17408 13855 17460 13864
rect 17408 13821 17417 13855
rect 17417 13821 17451 13855
rect 17451 13821 17460 13855
rect 17408 13812 17460 13821
rect 17960 13812 18012 13864
rect 18696 13812 18748 13864
rect 19064 13812 19116 13864
rect 15108 13744 15160 13796
rect 15200 13744 15252 13796
rect 16120 13744 16172 13796
rect 18328 13787 18380 13796
rect 13912 13676 13964 13728
rect 15568 13676 15620 13728
rect 15660 13676 15712 13728
rect 18328 13753 18337 13787
rect 18337 13753 18371 13787
rect 18371 13753 18380 13787
rect 18328 13744 18380 13753
rect 18788 13676 18840 13728
rect 19708 13812 19760 13864
rect 21548 13855 21600 13864
rect 21548 13821 21557 13855
rect 21557 13821 21591 13855
rect 21591 13821 21600 13855
rect 21548 13812 21600 13821
rect 21364 13787 21416 13796
rect 21364 13753 21373 13787
rect 21373 13753 21407 13787
rect 21407 13753 21416 13787
rect 21364 13744 21416 13753
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 2136 13515 2188 13524
rect 2136 13481 2145 13515
rect 2145 13481 2179 13515
rect 2179 13481 2188 13515
rect 2136 13472 2188 13481
rect 2320 13472 2372 13524
rect 3332 13515 3384 13524
rect 3332 13481 3341 13515
rect 3341 13481 3375 13515
rect 3375 13481 3384 13515
rect 3332 13472 3384 13481
rect 4344 13472 4396 13524
rect 5264 13515 5316 13524
rect 5264 13481 5273 13515
rect 5273 13481 5307 13515
rect 5307 13481 5316 13515
rect 5264 13472 5316 13481
rect 5908 13515 5960 13524
rect 5908 13481 5917 13515
rect 5917 13481 5951 13515
rect 5951 13481 5960 13515
rect 5908 13472 5960 13481
rect 3056 13404 3108 13456
rect 4896 13404 4948 13456
rect 4988 13404 5040 13456
rect 5356 13447 5408 13456
rect 5356 13413 5365 13447
rect 5365 13413 5399 13447
rect 5399 13413 5408 13447
rect 5356 13404 5408 13413
rect 6920 13404 6972 13456
rect 7196 13472 7248 13524
rect 8576 13515 8628 13524
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 9036 13472 9088 13524
rect 1952 13379 2004 13388
rect 1952 13345 1961 13379
rect 1961 13345 1995 13379
rect 1995 13345 2004 13379
rect 1952 13336 2004 13345
rect 2412 13336 2464 13388
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 2872 13379 2924 13388
rect 2872 13345 2881 13379
rect 2881 13345 2915 13379
rect 2915 13345 2924 13379
rect 2872 13336 2924 13345
rect 2964 13336 3016 13388
rect 3976 13336 4028 13388
rect 4436 13336 4488 13388
rect 1768 13200 1820 13252
rect 1400 13132 1452 13184
rect 1860 13175 1912 13184
rect 1860 13141 1869 13175
rect 1869 13141 1903 13175
rect 1903 13141 1912 13175
rect 1860 13132 1912 13141
rect 3240 13268 3292 13320
rect 5816 13336 5868 13388
rect 6184 13336 6236 13388
rect 6828 13336 6880 13388
rect 7656 13404 7708 13456
rect 8392 13336 8444 13388
rect 5908 13268 5960 13320
rect 8852 13404 8904 13456
rect 10140 13472 10192 13524
rect 11796 13472 11848 13524
rect 11888 13472 11940 13524
rect 12164 13472 12216 13524
rect 12348 13472 12400 13524
rect 12992 13472 13044 13524
rect 13636 13472 13688 13524
rect 14556 13515 14608 13524
rect 14556 13481 14565 13515
rect 14565 13481 14599 13515
rect 14599 13481 14608 13515
rect 14556 13472 14608 13481
rect 11060 13404 11112 13456
rect 13544 13404 13596 13456
rect 6644 13200 6696 13252
rect 5540 13132 5592 13184
rect 8576 13200 8628 13252
rect 9312 13336 9364 13388
rect 9404 13336 9456 13388
rect 10876 13379 10928 13388
rect 10876 13345 10910 13379
rect 10910 13345 10928 13379
rect 10876 13336 10928 13345
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 12716 13336 12768 13388
rect 15016 13404 15068 13456
rect 15936 13472 15988 13524
rect 16212 13515 16264 13524
rect 16212 13481 16221 13515
rect 16221 13481 16255 13515
rect 16255 13481 16264 13515
rect 16212 13472 16264 13481
rect 16856 13515 16908 13524
rect 16856 13481 16865 13515
rect 16865 13481 16899 13515
rect 16899 13481 16908 13515
rect 16856 13472 16908 13481
rect 18328 13472 18380 13524
rect 16028 13404 16080 13456
rect 16120 13404 16172 13456
rect 18788 13447 18840 13456
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 14556 13336 14608 13388
rect 18788 13413 18797 13447
rect 18797 13413 18831 13447
rect 18831 13413 18840 13447
rect 18788 13404 18840 13413
rect 19432 13472 19484 13524
rect 20444 13404 20496 13456
rect 17868 13336 17920 13388
rect 18144 13336 18196 13388
rect 18696 13336 18748 13388
rect 20260 13336 20312 13388
rect 21548 13379 21600 13388
rect 8300 13132 8352 13184
rect 10232 13200 10284 13252
rect 13268 13243 13320 13252
rect 13268 13209 13277 13243
rect 13277 13209 13311 13243
rect 13311 13209 13320 13243
rect 13268 13200 13320 13209
rect 14832 13268 14884 13320
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 16488 13311 16540 13320
rect 16488 13277 16497 13311
rect 16497 13277 16531 13311
rect 16531 13277 16540 13311
rect 16488 13268 16540 13277
rect 17224 13311 17276 13320
rect 17224 13277 17233 13311
rect 17233 13277 17267 13311
rect 17267 13277 17276 13311
rect 17224 13268 17276 13277
rect 17776 13268 17828 13320
rect 18880 13268 18932 13320
rect 15752 13200 15804 13252
rect 17408 13200 17460 13252
rect 11704 13132 11756 13184
rect 12256 13132 12308 13184
rect 12624 13132 12676 13184
rect 16212 13132 16264 13184
rect 18052 13132 18104 13184
rect 21548 13345 21557 13379
rect 21557 13345 21591 13379
rect 21591 13345 21600 13379
rect 21548 13336 21600 13345
rect 20904 13132 20956 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 1952 12971 2004 12980
rect 1952 12937 1961 12971
rect 1961 12937 1995 12971
rect 1995 12937 2004 12971
rect 1952 12928 2004 12937
rect 4344 12928 4396 12980
rect 5724 12928 5776 12980
rect 6460 12971 6512 12980
rect 6460 12937 6469 12971
rect 6469 12937 6503 12971
rect 6503 12937 6512 12971
rect 6460 12928 6512 12937
rect 7012 12928 7064 12980
rect 8668 12928 8720 12980
rect 9036 12928 9088 12980
rect 9864 12928 9916 12980
rect 10692 12928 10744 12980
rect 11980 12928 12032 12980
rect 14004 12928 14056 12980
rect 15752 12971 15804 12980
rect 9588 12860 9640 12912
rect 4068 12792 4120 12844
rect 5724 12792 5776 12844
rect 5816 12792 5868 12844
rect 6644 12792 6696 12844
rect 7564 12835 7616 12844
rect 7564 12801 7573 12835
rect 7573 12801 7607 12835
rect 7607 12801 7616 12835
rect 7564 12792 7616 12801
rect 10140 12792 10192 12844
rect 10876 12835 10928 12844
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 1952 12656 2004 12708
rect 2780 12724 2832 12776
rect 3976 12724 4028 12776
rect 5080 12724 5132 12776
rect 5908 12724 5960 12776
rect 6184 12724 6236 12776
rect 7840 12724 7892 12776
rect 8300 12724 8352 12776
rect 9496 12724 9548 12776
rect 9588 12724 9640 12776
rect 2872 12656 2924 12708
rect 3240 12656 3292 12708
rect 4988 12656 5040 12708
rect 7104 12656 7156 12708
rect 7748 12656 7800 12708
rect 9312 12656 9364 12708
rect 10508 12767 10560 12776
rect 10508 12733 10517 12767
rect 10517 12733 10551 12767
rect 10551 12733 10560 12767
rect 10508 12724 10560 12733
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 11244 12792 11296 12844
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 12716 12792 12768 12844
rect 13636 12792 13688 12844
rect 15752 12937 15761 12971
rect 15761 12937 15795 12971
rect 15795 12937 15804 12971
rect 15752 12928 15804 12937
rect 17776 12971 17828 12980
rect 17776 12937 17785 12971
rect 17785 12937 17819 12971
rect 17819 12937 17828 12971
rect 17776 12928 17828 12937
rect 17868 12928 17920 12980
rect 21364 12928 21416 12980
rect 15200 12860 15252 12912
rect 14832 12792 14884 12844
rect 16488 12860 16540 12912
rect 18880 12860 18932 12912
rect 16028 12792 16080 12844
rect 16396 12835 16448 12844
rect 16396 12801 16405 12835
rect 16405 12801 16439 12835
rect 16439 12801 16448 12835
rect 16396 12792 16448 12801
rect 11888 12656 11940 12708
rect 16028 12656 16080 12708
rect 16396 12656 16448 12708
rect 2964 12588 3016 12640
rect 3976 12631 4028 12640
rect 3976 12597 3985 12631
rect 3985 12597 4019 12631
rect 4019 12597 4028 12631
rect 4344 12631 4396 12640
rect 3976 12588 4028 12597
rect 4344 12597 4353 12631
rect 4353 12597 4387 12631
rect 4387 12597 4396 12631
rect 4344 12588 4396 12597
rect 4896 12588 4948 12640
rect 5264 12588 5316 12640
rect 5540 12588 5592 12640
rect 6184 12588 6236 12640
rect 6644 12588 6696 12640
rect 8208 12588 8260 12640
rect 8576 12588 8628 12640
rect 10968 12588 11020 12640
rect 13084 12631 13136 12640
rect 13084 12597 13093 12631
rect 13093 12597 13127 12631
rect 13127 12597 13136 12631
rect 13084 12588 13136 12597
rect 13268 12588 13320 12640
rect 13636 12588 13688 12640
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 14004 12588 14056 12640
rect 16948 12724 17000 12776
rect 17408 12767 17460 12776
rect 17408 12733 17417 12767
rect 17417 12733 17451 12767
rect 17451 12733 17460 12767
rect 17408 12724 17460 12733
rect 21548 12835 21600 12844
rect 21548 12801 21557 12835
rect 21557 12801 21591 12835
rect 21591 12801 21600 12835
rect 21548 12792 21600 12801
rect 16856 12656 16908 12708
rect 17500 12656 17552 12708
rect 18880 12724 18932 12776
rect 19064 12724 19116 12776
rect 20168 12724 20220 12776
rect 19432 12656 19484 12708
rect 20720 12656 20772 12708
rect 19248 12588 19300 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 2596 12427 2648 12436
rect 2596 12393 2605 12427
rect 2605 12393 2639 12427
rect 2639 12393 2648 12427
rect 2596 12384 2648 12393
rect 3976 12427 4028 12436
rect 3976 12393 3985 12427
rect 3985 12393 4019 12427
rect 4019 12393 4028 12427
rect 3976 12384 4028 12393
rect 1400 12248 1452 12300
rect 2228 12291 2280 12300
rect 2228 12257 2237 12291
rect 2237 12257 2271 12291
rect 2271 12257 2280 12291
rect 2228 12248 2280 12257
rect 3608 12248 3660 12300
rect 4068 12316 4120 12368
rect 4160 12248 4212 12300
rect 4896 12316 4948 12368
rect 5080 12316 5132 12368
rect 5356 12316 5408 12368
rect 5724 12384 5776 12436
rect 9220 12384 9272 12436
rect 9588 12427 9640 12436
rect 9588 12393 9597 12427
rect 9597 12393 9631 12427
rect 9631 12393 9640 12427
rect 9588 12384 9640 12393
rect 10048 12427 10100 12436
rect 10048 12393 10057 12427
rect 10057 12393 10091 12427
rect 10091 12393 10100 12427
rect 10048 12384 10100 12393
rect 10140 12384 10192 12436
rect 10876 12384 10928 12436
rect 11796 12384 11848 12436
rect 12072 12384 12124 12436
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 12900 12384 12952 12436
rect 13360 12384 13412 12436
rect 13452 12384 13504 12436
rect 15200 12384 15252 12436
rect 16396 12384 16448 12436
rect 16856 12384 16908 12436
rect 17592 12384 17644 12436
rect 19248 12427 19300 12436
rect 19248 12393 19257 12427
rect 19257 12393 19291 12427
rect 19291 12393 19300 12427
rect 19248 12384 19300 12393
rect 19984 12384 20036 12436
rect 20168 12427 20220 12436
rect 20168 12393 20177 12427
rect 20177 12393 20211 12427
rect 20211 12393 20220 12427
rect 20168 12384 20220 12393
rect 6460 12316 6512 12368
rect 1952 12223 2004 12232
rect 1952 12189 1961 12223
rect 1961 12189 1995 12223
rect 1995 12189 2004 12223
rect 1952 12180 2004 12189
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 5264 12248 5316 12300
rect 5448 12248 5500 12300
rect 6828 12248 6880 12300
rect 7380 12248 7432 12300
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 7564 12248 7616 12257
rect 8024 12316 8076 12368
rect 10508 12316 10560 12368
rect 11336 12316 11388 12368
rect 8300 12248 8352 12300
rect 2596 12044 2648 12096
rect 8024 12180 8076 12232
rect 8208 12180 8260 12232
rect 9036 12248 9088 12300
rect 10876 12248 10928 12300
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 12164 12291 12216 12300
rect 11704 12248 11756 12257
rect 12164 12257 12173 12291
rect 12173 12257 12207 12291
rect 12207 12257 12216 12291
rect 12164 12248 12216 12257
rect 12716 12316 12768 12368
rect 13084 12359 13136 12368
rect 13084 12325 13096 12359
rect 13096 12325 13136 12359
rect 13084 12316 13136 12325
rect 13268 12316 13320 12368
rect 13636 12316 13688 12368
rect 14004 12316 14056 12368
rect 14556 12359 14608 12368
rect 14556 12325 14565 12359
rect 14565 12325 14599 12359
rect 14599 12325 14608 12359
rect 14556 12316 14608 12325
rect 14740 12316 14792 12368
rect 16488 12316 16540 12368
rect 16764 12316 16816 12368
rect 9772 12180 9824 12232
rect 10048 12180 10100 12232
rect 5356 12155 5408 12164
rect 5356 12121 5365 12155
rect 5365 12121 5399 12155
rect 5399 12121 5408 12155
rect 5356 12112 5408 12121
rect 7104 12112 7156 12164
rect 9864 12112 9916 12164
rect 4896 12044 4948 12096
rect 5540 12087 5592 12096
rect 5540 12053 5549 12087
rect 5549 12053 5583 12087
rect 5583 12053 5592 12087
rect 5540 12044 5592 12053
rect 7196 12087 7248 12096
rect 7196 12053 7205 12087
rect 7205 12053 7239 12087
rect 7239 12053 7248 12087
rect 7196 12044 7248 12053
rect 7748 12044 7800 12096
rect 8760 12044 8812 12096
rect 10232 12180 10284 12232
rect 10416 12180 10468 12232
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 14740 12223 14792 12232
rect 12072 12180 12124 12189
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 14740 12180 14792 12189
rect 16580 12180 16632 12232
rect 17500 12291 17552 12300
rect 17500 12257 17509 12291
rect 17509 12257 17543 12291
rect 17543 12257 17552 12291
rect 17500 12248 17552 12257
rect 18052 12248 18104 12300
rect 18788 12316 18840 12368
rect 21180 12359 21232 12368
rect 21180 12325 21189 12359
rect 21189 12325 21223 12359
rect 21223 12325 21232 12359
rect 21180 12316 21232 12325
rect 19708 12248 19760 12300
rect 19984 12291 20036 12300
rect 19984 12257 19993 12291
rect 19993 12257 20027 12291
rect 20027 12257 20036 12291
rect 19984 12248 20036 12257
rect 20996 12291 21048 12300
rect 20996 12257 21005 12291
rect 21005 12257 21039 12291
rect 21039 12257 21048 12291
rect 20996 12248 21048 12257
rect 16764 12223 16816 12232
rect 16764 12189 16773 12223
rect 16773 12189 16807 12223
rect 16807 12189 16816 12223
rect 16764 12180 16816 12189
rect 18604 12180 18656 12232
rect 20812 12180 20864 12232
rect 16028 12112 16080 12164
rect 16948 12112 17000 12164
rect 18512 12112 18564 12164
rect 20260 12112 20312 12164
rect 21548 12155 21600 12164
rect 21548 12121 21557 12155
rect 21557 12121 21591 12155
rect 21591 12121 21600 12155
rect 21548 12112 21600 12121
rect 11980 12044 12032 12096
rect 12348 12044 12400 12096
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 14280 12044 14332 12096
rect 15844 12044 15896 12096
rect 17132 12044 17184 12096
rect 17684 12044 17736 12096
rect 18604 12044 18656 12096
rect 18696 12044 18748 12096
rect 18880 12087 18932 12096
rect 18880 12053 18889 12087
rect 18889 12053 18923 12087
rect 18923 12053 18932 12087
rect 18880 12044 18932 12053
rect 19156 12044 19208 12096
rect 20168 12044 20220 12096
rect 20628 12044 20680 12096
rect 21456 12044 21508 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 1952 11840 2004 11892
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 3056 11840 3108 11892
rect 3608 11883 3660 11892
rect 3608 11849 3617 11883
rect 3617 11849 3651 11883
rect 3651 11849 3660 11883
rect 3608 11840 3660 11849
rect 4252 11840 4304 11892
rect 5632 11840 5684 11892
rect 6460 11883 6512 11892
rect 6460 11849 6469 11883
rect 6469 11849 6503 11883
rect 6503 11849 6512 11883
rect 6460 11840 6512 11849
rect 7932 11840 7984 11892
rect 9220 11840 9272 11892
rect 10600 11840 10652 11892
rect 12072 11840 12124 11892
rect 14464 11840 14516 11892
rect 14740 11840 14792 11892
rect 7840 11772 7892 11824
rect 2872 11747 2924 11756
rect 2872 11713 2881 11747
rect 2881 11713 2915 11747
rect 2915 11713 2924 11747
rect 2872 11704 2924 11713
rect 3700 11704 3752 11756
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 5540 11704 5592 11756
rect 6552 11704 6604 11756
rect 8300 11704 8352 11756
rect 8852 11772 8904 11824
rect 2596 11679 2648 11688
rect 2596 11645 2614 11679
rect 2614 11645 2648 11679
rect 2596 11636 2648 11645
rect 4896 11679 4948 11688
rect 2044 11568 2096 11620
rect 2964 11500 3016 11552
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 7196 11636 7248 11688
rect 8576 11636 8628 11688
rect 9036 11704 9088 11756
rect 9772 11704 9824 11756
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 12532 11772 12584 11824
rect 15568 11840 15620 11892
rect 11152 11704 11204 11756
rect 11244 11704 11296 11756
rect 12716 11747 12768 11756
rect 12716 11713 12725 11747
rect 12725 11713 12759 11747
rect 12759 11713 12768 11747
rect 12716 11704 12768 11713
rect 10508 11636 10560 11688
rect 3608 11500 3660 11552
rect 3884 11500 3936 11552
rect 4160 11500 4212 11552
rect 4344 11568 4396 11620
rect 5632 11568 5684 11620
rect 7472 11568 7524 11620
rect 8024 11568 8076 11620
rect 5540 11500 5592 11552
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 6644 11500 6696 11552
rect 6828 11500 6880 11552
rect 8300 11543 8352 11552
rect 8300 11509 8309 11543
rect 8309 11509 8343 11543
rect 8343 11509 8352 11543
rect 8300 11500 8352 11509
rect 8576 11500 8628 11552
rect 8760 11500 8812 11552
rect 8852 11500 8904 11552
rect 9496 11500 9548 11552
rect 10692 11500 10744 11552
rect 11060 11568 11112 11620
rect 11980 11568 12032 11620
rect 14280 11636 14332 11688
rect 16304 11636 16356 11688
rect 16028 11568 16080 11620
rect 16672 11568 16724 11620
rect 18144 11840 18196 11892
rect 19984 11883 20036 11892
rect 18052 11772 18104 11824
rect 16948 11679 17000 11688
rect 16948 11645 16957 11679
rect 16957 11645 16991 11679
rect 16991 11645 17000 11679
rect 16948 11636 17000 11645
rect 17500 11636 17552 11688
rect 18052 11636 18104 11688
rect 18880 11747 18932 11756
rect 18880 11713 18889 11747
rect 18889 11713 18923 11747
rect 18923 11713 18932 11747
rect 18880 11704 18932 11713
rect 19064 11747 19116 11756
rect 19064 11713 19073 11747
rect 19073 11713 19107 11747
rect 19107 11713 19116 11747
rect 19064 11704 19116 11713
rect 19524 11772 19576 11824
rect 19984 11849 19993 11883
rect 19993 11849 20027 11883
rect 20027 11849 20036 11883
rect 19984 11840 20036 11849
rect 20260 11883 20312 11892
rect 20260 11849 20269 11883
rect 20269 11849 20303 11883
rect 20303 11849 20312 11883
rect 20260 11840 20312 11849
rect 20720 11883 20772 11892
rect 20720 11849 20729 11883
rect 20729 11849 20763 11883
rect 20763 11849 20772 11883
rect 20720 11840 20772 11849
rect 20996 11883 21048 11892
rect 20996 11849 21005 11883
rect 21005 11849 21039 11883
rect 21039 11849 21048 11883
rect 20996 11840 21048 11849
rect 21456 11704 21508 11756
rect 19800 11636 19852 11688
rect 20444 11679 20496 11688
rect 20444 11645 20453 11679
rect 20453 11645 20487 11679
rect 20487 11645 20496 11679
rect 20444 11636 20496 11645
rect 20720 11636 20772 11688
rect 17408 11568 17460 11620
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 12808 11500 12860 11552
rect 13544 11543 13596 11552
rect 13544 11509 13553 11543
rect 13553 11509 13587 11543
rect 13587 11509 13596 11543
rect 13544 11500 13596 11509
rect 13636 11500 13688 11552
rect 16304 11543 16356 11552
rect 16304 11509 16313 11543
rect 16313 11509 16347 11543
rect 16347 11509 16356 11543
rect 16304 11500 16356 11509
rect 16396 11543 16448 11552
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16396 11500 16448 11509
rect 20628 11568 20680 11620
rect 21548 11568 21600 11620
rect 19156 11500 19208 11552
rect 20812 11500 20864 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 1676 11296 1728 11348
rect 2596 11296 2648 11348
rect 3240 11296 3292 11348
rect 3976 11296 4028 11348
rect 4068 11228 4120 11280
rect 1492 11203 1544 11212
rect 1492 11169 1501 11203
rect 1501 11169 1535 11203
rect 1535 11169 1544 11203
rect 1492 11160 1544 11169
rect 2872 11203 2924 11212
rect 2872 11169 2890 11203
rect 2890 11169 2924 11203
rect 3332 11203 3384 11212
rect 2872 11160 2924 11169
rect 3332 11169 3341 11203
rect 3341 11169 3375 11203
rect 3375 11169 3384 11203
rect 3332 11160 3384 11169
rect 4252 11203 4304 11212
rect 4252 11169 4261 11203
rect 4261 11169 4295 11203
rect 4295 11169 4304 11203
rect 4252 11160 4304 11169
rect 4896 11228 4948 11280
rect 5540 11228 5592 11280
rect 7380 11296 7432 11348
rect 7564 11296 7616 11348
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 9036 11296 9088 11348
rect 10600 11339 10652 11348
rect 6552 11228 6604 11280
rect 7104 11228 7156 11280
rect 4988 11160 5040 11212
rect 3884 11092 3936 11144
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 7472 11160 7524 11212
rect 9956 11228 10008 11280
rect 10600 11305 10609 11339
rect 10609 11305 10643 11339
rect 10643 11305 10652 11339
rect 10600 11296 10652 11305
rect 10876 11296 10928 11348
rect 6644 11135 6696 11144
rect 3700 11024 3752 11076
rect 6644 11101 6653 11135
rect 6653 11101 6687 11135
rect 6687 11101 6696 11135
rect 6644 11092 6696 11101
rect 9864 11092 9916 11144
rect 10048 11092 10100 11144
rect 10140 11092 10192 11144
rect 13176 11271 13228 11280
rect 10508 11160 10560 11212
rect 10692 11092 10744 11144
rect 11980 11160 12032 11212
rect 12440 11160 12492 11212
rect 11244 11135 11296 11144
rect 11244 11101 11253 11135
rect 11253 11101 11287 11135
rect 11287 11101 11296 11135
rect 11244 11092 11296 11101
rect 11612 11092 11664 11144
rect 11888 11092 11940 11144
rect 6092 11024 6144 11076
rect 8300 11024 8352 11076
rect 8576 11024 8628 11076
rect 9220 11024 9272 11076
rect 12164 11024 12216 11076
rect 13176 11237 13185 11271
rect 13185 11237 13219 11271
rect 13219 11237 13228 11271
rect 13176 11228 13228 11237
rect 13544 11296 13596 11348
rect 13728 11271 13780 11280
rect 13728 11237 13737 11271
rect 13737 11237 13771 11271
rect 13771 11237 13780 11271
rect 13728 11228 13780 11237
rect 15200 11228 15252 11280
rect 17684 11296 17736 11348
rect 17776 11339 17828 11348
rect 17776 11305 17785 11339
rect 17785 11305 17819 11339
rect 17819 11305 17828 11339
rect 17776 11296 17828 11305
rect 18052 11296 18104 11348
rect 18880 11296 18932 11348
rect 19156 11296 19208 11348
rect 19432 11296 19484 11348
rect 19800 11296 19852 11348
rect 12900 11160 12952 11212
rect 14924 11160 14976 11212
rect 16948 11228 17000 11280
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 14556 11092 14608 11144
rect 14832 11092 14884 11144
rect 13452 11024 13504 11076
rect 16028 11024 16080 11076
rect 5264 10956 5316 11008
rect 5724 10999 5776 11008
rect 5724 10965 5733 10999
rect 5733 10965 5767 10999
rect 5767 10965 5776 10999
rect 5724 10956 5776 10965
rect 6552 10999 6604 11008
rect 6552 10965 6561 10999
rect 6561 10965 6595 10999
rect 6595 10965 6604 10999
rect 6552 10956 6604 10965
rect 8024 10999 8076 11008
rect 8024 10965 8033 10999
rect 8033 10965 8067 10999
rect 8067 10965 8076 10999
rect 8024 10956 8076 10965
rect 13912 10956 13964 11008
rect 15200 10999 15252 11008
rect 15200 10965 15209 10999
rect 15209 10965 15243 10999
rect 15243 10965 15252 10999
rect 15200 10956 15252 10965
rect 15292 10956 15344 11008
rect 19616 11160 19668 11212
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 20444 11160 20496 11212
rect 21456 11203 21508 11212
rect 21456 11169 21465 11203
rect 21465 11169 21499 11203
rect 21499 11169 21508 11203
rect 21456 11160 21508 11169
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 19340 11092 19392 11144
rect 17408 11067 17460 11076
rect 17408 11033 17417 11067
rect 17417 11033 17451 11067
rect 17451 11033 17460 11067
rect 21088 11092 21140 11144
rect 21364 11092 21416 11144
rect 17408 11024 17460 11033
rect 20260 11024 20312 11076
rect 19156 10956 19208 11008
rect 19708 10956 19760 11008
rect 20812 10956 20864 11008
rect 22192 10956 22244 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 2228 10795 2280 10804
rect 2228 10761 2237 10795
rect 2237 10761 2271 10795
rect 2271 10761 2280 10795
rect 2228 10752 2280 10761
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 3884 10752 3936 10804
rect 4252 10752 4304 10804
rect 4160 10684 4212 10736
rect 5264 10752 5316 10804
rect 5632 10752 5684 10804
rect 5908 10752 5960 10804
rect 7380 10795 7432 10804
rect 7380 10761 7389 10795
rect 7389 10761 7423 10795
rect 7423 10761 7432 10795
rect 7380 10752 7432 10761
rect 4068 10548 4120 10600
rect 7104 10684 7156 10736
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 5632 10548 5684 10600
rect 5724 10548 5776 10600
rect 6552 10616 6604 10668
rect 2596 10523 2648 10532
rect 2596 10489 2630 10523
rect 2630 10489 2648 10523
rect 2596 10480 2648 10489
rect 3792 10480 3844 10532
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 2228 10412 2280 10464
rect 2872 10412 2924 10464
rect 3700 10455 3752 10464
rect 3700 10421 3709 10455
rect 3709 10421 3743 10455
rect 3743 10421 3752 10455
rect 3700 10412 3752 10421
rect 4528 10480 4580 10532
rect 5540 10480 5592 10532
rect 6460 10480 6512 10532
rect 4252 10455 4304 10464
rect 4252 10421 4261 10455
rect 4261 10421 4295 10455
rect 4295 10421 4304 10455
rect 4252 10412 4304 10421
rect 5356 10412 5408 10464
rect 6000 10455 6052 10464
rect 6000 10421 6009 10455
rect 6009 10421 6043 10455
rect 6043 10421 6052 10455
rect 7564 10727 7616 10736
rect 7564 10693 7573 10727
rect 7573 10693 7607 10727
rect 7607 10693 7616 10727
rect 7564 10684 7616 10693
rect 7656 10616 7708 10668
rect 8024 10616 8076 10668
rect 8760 10684 8812 10736
rect 9680 10684 9732 10736
rect 8852 10548 8904 10600
rect 9496 10616 9548 10668
rect 9772 10616 9824 10668
rect 11244 10752 11296 10804
rect 11980 10752 12032 10804
rect 13268 10752 13320 10804
rect 11060 10684 11112 10736
rect 9680 10548 9732 10600
rect 9956 10591 10008 10600
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 9956 10548 10008 10557
rect 11612 10616 11664 10668
rect 12072 10616 12124 10668
rect 13636 10684 13688 10736
rect 14372 10752 14424 10804
rect 14740 10752 14792 10804
rect 14924 10684 14976 10736
rect 14556 10616 14608 10668
rect 7748 10480 7800 10532
rect 6000 10412 6052 10421
rect 7564 10412 7616 10464
rect 9128 10480 9180 10532
rect 10508 10480 10560 10532
rect 11152 10480 11204 10532
rect 12348 10480 12400 10532
rect 12716 10548 12768 10600
rect 13268 10591 13320 10600
rect 13268 10557 13286 10591
rect 13286 10557 13320 10591
rect 13268 10548 13320 10557
rect 13452 10548 13504 10600
rect 13912 10548 13964 10600
rect 14096 10548 14148 10600
rect 14740 10548 14792 10600
rect 16304 10752 16356 10804
rect 16764 10752 16816 10804
rect 16396 10684 16448 10736
rect 19248 10752 19300 10804
rect 19984 10752 20036 10804
rect 20444 10795 20496 10804
rect 20444 10761 20453 10795
rect 20453 10761 20487 10795
rect 20487 10761 20496 10795
rect 20444 10752 20496 10761
rect 20720 10795 20772 10804
rect 20720 10761 20729 10795
rect 20729 10761 20763 10795
rect 20763 10761 20772 10795
rect 20720 10752 20772 10761
rect 16028 10616 16080 10668
rect 17592 10659 17644 10668
rect 17592 10625 17601 10659
rect 17601 10625 17635 10659
rect 17635 10625 17644 10659
rect 17592 10616 17644 10625
rect 17960 10659 18012 10668
rect 17960 10625 17969 10659
rect 17969 10625 18003 10659
rect 18003 10625 18012 10659
rect 17960 10616 18012 10625
rect 19892 10616 19944 10668
rect 16948 10548 17000 10600
rect 17316 10591 17368 10600
rect 17316 10557 17325 10591
rect 17325 10557 17359 10591
rect 17359 10557 17368 10591
rect 17316 10548 17368 10557
rect 17684 10548 17736 10600
rect 18880 10548 18932 10600
rect 19156 10548 19208 10600
rect 15292 10480 15344 10532
rect 8852 10412 8904 10464
rect 9312 10412 9364 10464
rect 10968 10412 11020 10464
rect 12808 10412 12860 10464
rect 13728 10412 13780 10464
rect 14096 10455 14148 10464
rect 14096 10421 14105 10455
rect 14105 10421 14139 10455
rect 14139 10421 14148 10455
rect 14096 10412 14148 10421
rect 14556 10455 14608 10464
rect 14556 10421 14565 10455
rect 14565 10421 14599 10455
rect 14599 10421 14608 10455
rect 14556 10412 14608 10421
rect 16488 10455 16540 10464
rect 16488 10421 16497 10455
rect 16497 10421 16531 10455
rect 16531 10421 16540 10455
rect 17776 10480 17828 10532
rect 21088 10523 21140 10532
rect 16488 10412 16540 10421
rect 17224 10412 17276 10464
rect 18972 10412 19024 10464
rect 19708 10455 19760 10464
rect 19708 10421 19717 10455
rect 19717 10421 19751 10455
rect 19751 10421 19760 10455
rect 19708 10412 19760 10421
rect 19800 10455 19852 10464
rect 19800 10421 19809 10455
rect 19809 10421 19843 10455
rect 19843 10421 19852 10455
rect 21088 10489 21097 10523
rect 21097 10489 21131 10523
rect 21131 10489 21140 10523
rect 21088 10480 21140 10489
rect 21180 10480 21232 10532
rect 21456 10523 21508 10532
rect 21456 10489 21465 10523
rect 21465 10489 21499 10523
rect 21499 10489 21508 10523
rect 21456 10480 21508 10489
rect 19800 10412 19852 10421
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 3332 10208 3384 10260
rect 4068 10208 4120 10260
rect 4344 10208 4396 10260
rect 2872 10140 2924 10192
rect 3792 10140 3844 10192
rect 4988 10140 5040 10192
rect 6460 10208 6512 10260
rect 8208 10208 8260 10260
rect 8300 10208 8352 10260
rect 9588 10208 9640 10260
rect 10968 10251 11020 10260
rect 10968 10217 10977 10251
rect 10977 10217 11011 10251
rect 11011 10217 11020 10251
rect 10968 10208 11020 10217
rect 6000 10140 6052 10192
rect 6920 10140 6972 10192
rect 11796 10208 11848 10260
rect 14096 10208 14148 10260
rect 14556 10208 14608 10260
rect 15292 10251 15344 10260
rect 15292 10217 15301 10251
rect 15301 10217 15335 10251
rect 15335 10217 15344 10251
rect 15292 10208 15344 10217
rect 15660 10251 15712 10260
rect 15660 10217 15669 10251
rect 15669 10217 15703 10251
rect 15703 10217 15712 10251
rect 15660 10208 15712 10217
rect 16488 10208 16540 10260
rect 17316 10208 17368 10260
rect 17960 10208 18012 10260
rect 18972 10251 19024 10260
rect 18972 10217 18981 10251
rect 18981 10217 19015 10251
rect 19015 10217 19024 10251
rect 18972 10208 19024 10217
rect 19064 10208 19116 10260
rect 3148 10072 3200 10124
rect 3424 10072 3476 10124
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2136 10004 2188 10056
rect 2504 10004 2556 10056
rect 2228 9979 2280 9988
rect 2228 9945 2237 9979
rect 2237 9945 2271 9979
rect 2271 9945 2280 9979
rect 2228 9936 2280 9945
rect 2596 9936 2648 9988
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 4528 10004 4580 10056
rect 5264 10004 5316 10056
rect 5540 10072 5592 10124
rect 6276 10072 6328 10124
rect 7104 10115 7156 10124
rect 7104 10081 7113 10115
rect 7113 10081 7147 10115
rect 7147 10081 7156 10115
rect 7104 10072 7156 10081
rect 5816 10004 5868 10056
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 7196 10004 7248 10056
rect 7656 10004 7708 10056
rect 8208 10004 8260 10056
rect 4252 9936 4304 9988
rect 9220 10004 9272 10056
rect 8484 9936 8536 9988
rect 9312 9936 9364 9988
rect 7012 9868 7064 9920
rect 7564 9868 7616 9920
rect 8024 9868 8076 9920
rect 8300 9868 8352 9920
rect 9220 9868 9272 9920
rect 9772 10072 9824 10124
rect 10600 10004 10652 10056
rect 10968 10004 11020 10056
rect 12164 10140 12216 10192
rect 12532 10140 12584 10192
rect 17592 10140 17644 10192
rect 13268 10072 13320 10124
rect 13544 10115 13596 10124
rect 13544 10081 13562 10115
rect 13562 10081 13596 10115
rect 13544 10072 13596 10081
rect 13728 10072 13780 10124
rect 13912 10072 13964 10124
rect 15476 10072 15528 10124
rect 15752 10115 15804 10124
rect 15752 10081 15761 10115
rect 15761 10081 15795 10115
rect 15795 10081 15804 10115
rect 15752 10072 15804 10081
rect 11244 9936 11296 9988
rect 10968 9868 11020 9920
rect 14004 10004 14056 10056
rect 14740 10004 14792 10056
rect 16304 10072 16356 10124
rect 19340 10072 19392 10124
rect 19892 10115 19944 10124
rect 19892 10081 19926 10115
rect 19926 10081 19944 10115
rect 19892 10072 19944 10081
rect 20444 10072 20496 10124
rect 21640 10072 21692 10124
rect 12716 9868 12768 9920
rect 14280 9936 14332 9988
rect 17592 10004 17644 10056
rect 19064 10004 19116 10056
rect 21364 9979 21416 9988
rect 21364 9945 21373 9979
rect 21373 9945 21407 9979
rect 21407 9945 21416 9979
rect 21364 9936 21416 9945
rect 14832 9868 14884 9920
rect 15660 9868 15712 9920
rect 19248 9868 19300 9920
rect 19432 9911 19484 9920
rect 19432 9877 19441 9911
rect 19441 9877 19475 9911
rect 19475 9877 19484 9911
rect 19432 9868 19484 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 1768 9664 1820 9716
rect 3792 9664 3844 9716
rect 6552 9664 6604 9716
rect 10508 9707 10560 9716
rect 2688 9596 2740 9648
rect 3976 9596 4028 9648
rect 6644 9596 6696 9648
rect 8944 9639 8996 9648
rect 8944 9605 8953 9639
rect 8953 9605 8987 9639
rect 8987 9605 8996 9639
rect 8944 9596 8996 9605
rect 10508 9673 10517 9707
rect 10517 9673 10551 9707
rect 10551 9673 10560 9707
rect 10508 9664 10560 9673
rect 1676 9528 1728 9580
rect 2596 9528 2648 9580
rect 4160 9571 4212 9580
rect 4160 9537 4169 9571
rect 4169 9537 4203 9571
rect 4203 9537 4212 9571
rect 4160 9528 4212 9537
rect 5080 9528 5132 9580
rect 7472 9528 7524 9580
rect 11244 9596 11296 9648
rect 12164 9664 12216 9716
rect 12440 9664 12492 9716
rect 13176 9664 13228 9716
rect 14004 9596 14056 9648
rect 2872 9460 2924 9512
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 5448 9460 5500 9512
rect 6092 9460 6144 9512
rect 6644 9503 6696 9512
rect 1492 9367 1544 9376
rect 1492 9333 1501 9367
rect 1501 9333 1535 9367
rect 1535 9333 1544 9367
rect 1492 9324 1544 9333
rect 2320 9324 2372 9376
rect 3056 9324 3108 9376
rect 3516 9392 3568 9444
rect 4068 9392 4120 9444
rect 4896 9392 4948 9444
rect 5264 9392 5316 9444
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 7012 9460 7064 9512
rect 3608 9367 3660 9376
rect 3608 9333 3617 9367
rect 3617 9333 3651 9367
rect 3651 9333 3660 9367
rect 3608 9324 3660 9333
rect 5632 9324 5684 9376
rect 5908 9324 5960 9376
rect 6092 9324 6144 9376
rect 7012 9367 7064 9376
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 7012 9324 7064 9333
rect 7196 9324 7248 9376
rect 8208 9435 8260 9444
rect 8208 9401 8237 9435
rect 8237 9401 8260 9435
rect 8208 9392 8260 9401
rect 9036 9460 9088 9512
rect 9956 9460 10008 9512
rect 10600 9460 10652 9512
rect 9220 9392 9272 9444
rect 11980 9528 12032 9580
rect 13176 9528 13228 9580
rect 13728 9528 13780 9580
rect 14280 9596 14332 9648
rect 14556 9596 14608 9648
rect 15568 9596 15620 9648
rect 15660 9596 15712 9648
rect 16580 9596 16632 9648
rect 16948 9639 17000 9648
rect 16948 9605 16957 9639
rect 16957 9605 16991 9639
rect 16991 9605 17000 9639
rect 16948 9596 17000 9605
rect 17960 9664 18012 9716
rect 18604 9664 18656 9716
rect 18972 9664 19024 9716
rect 19708 9664 19760 9716
rect 18788 9596 18840 9648
rect 20444 9639 20496 9648
rect 20444 9605 20453 9639
rect 20453 9605 20487 9639
rect 20487 9605 20496 9639
rect 20444 9596 20496 9605
rect 10968 9503 11020 9512
rect 10968 9469 10977 9503
rect 10977 9469 11011 9503
rect 11011 9469 11020 9503
rect 10968 9460 11020 9469
rect 11612 9460 11664 9512
rect 12992 9460 13044 9512
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 12532 9392 12584 9444
rect 12808 9435 12860 9444
rect 12808 9401 12848 9435
rect 12848 9401 12860 9435
rect 14280 9460 14332 9512
rect 14648 9460 14700 9512
rect 15200 9460 15252 9512
rect 16672 9528 16724 9580
rect 17592 9571 17644 9580
rect 17592 9537 17601 9571
rect 17601 9537 17635 9571
rect 17635 9537 17644 9571
rect 17592 9528 17644 9537
rect 16120 9460 16172 9512
rect 16764 9503 16816 9512
rect 16764 9469 16773 9503
rect 16773 9469 16807 9503
rect 16807 9469 16816 9503
rect 16764 9460 16816 9469
rect 18696 9460 18748 9512
rect 19064 9503 19116 9512
rect 19064 9469 19073 9503
rect 19073 9469 19107 9503
rect 19107 9469 19116 9503
rect 19064 9460 19116 9469
rect 21088 9528 21140 9580
rect 21548 9503 21600 9512
rect 21548 9469 21557 9503
rect 21557 9469 21591 9503
rect 21591 9469 21600 9503
rect 21548 9460 21600 9469
rect 12808 9392 12860 9401
rect 10968 9324 11020 9376
rect 11152 9324 11204 9376
rect 11704 9367 11756 9376
rect 11704 9333 11713 9367
rect 11713 9333 11747 9367
rect 11747 9333 11756 9367
rect 11704 9324 11756 9333
rect 13084 9324 13136 9376
rect 13360 9367 13412 9376
rect 13360 9333 13369 9367
rect 13369 9333 13403 9367
rect 13403 9333 13412 9367
rect 14556 9392 14608 9444
rect 14832 9435 14884 9444
rect 14832 9401 14841 9435
rect 14841 9401 14875 9435
rect 14875 9401 14884 9435
rect 14832 9392 14884 9401
rect 17960 9435 18012 9444
rect 13360 9324 13412 9333
rect 13728 9324 13780 9376
rect 14648 9324 14700 9376
rect 15476 9324 15528 9376
rect 17960 9401 17969 9435
rect 17969 9401 18003 9435
rect 18003 9401 18012 9435
rect 17960 9392 18012 9401
rect 20260 9392 20312 9444
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 18512 9367 18564 9376
rect 18512 9333 18521 9367
rect 18521 9333 18555 9367
rect 18555 9333 18564 9367
rect 18512 9324 18564 9333
rect 19800 9324 19852 9376
rect 20904 9367 20956 9376
rect 20904 9333 20913 9367
rect 20913 9333 20947 9367
rect 20947 9333 20956 9367
rect 20904 9324 20956 9333
rect 20996 9367 21048 9376
rect 20996 9333 21005 9367
rect 21005 9333 21039 9367
rect 21039 9333 21048 9367
rect 21364 9367 21416 9376
rect 20996 9324 21048 9333
rect 21364 9333 21373 9367
rect 21373 9333 21407 9367
rect 21407 9333 21416 9367
rect 21364 9324 21416 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 3148 9120 3200 9172
rect 3700 9052 3752 9104
rect 2320 8984 2372 9036
rect 2688 9027 2740 9036
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 2688 8984 2740 8993
rect 3148 9027 3200 9036
rect 3148 8993 3157 9027
rect 3157 8993 3191 9027
rect 3191 8993 3200 9027
rect 3148 8984 3200 8993
rect 3608 8984 3660 9036
rect 2596 8916 2648 8968
rect 3240 8916 3292 8968
rect 5724 9120 5776 9172
rect 3884 9027 3936 9036
rect 3884 8993 3893 9027
rect 3893 8993 3927 9027
rect 3927 8993 3936 9027
rect 4160 9027 4212 9036
rect 3884 8984 3936 8993
rect 4160 8993 4194 9027
rect 4194 8993 4212 9027
rect 4160 8984 4212 8993
rect 5908 9027 5960 9036
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 6184 9027 6236 9036
rect 6184 8993 6218 9027
rect 6218 8993 6236 9027
rect 6184 8984 6236 8993
rect 7104 9120 7156 9172
rect 8944 9120 8996 9172
rect 6920 9052 6972 9104
rect 8760 9052 8812 9104
rect 10140 9120 10192 9172
rect 10324 9120 10376 9172
rect 10968 9120 11020 9172
rect 11152 9163 11204 9172
rect 11152 9129 11161 9163
rect 11161 9129 11195 9163
rect 11195 9129 11204 9163
rect 11152 9120 11204 9129
rect 11520 9120 11572 9172
rect 12440 9120 12492 9172
rect 12532 9120 12584 9172
rect 7932 8984 7984 9036
rect 8116 8984 8168 9036
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 8208 8916 8260 8968
rect 8576 8916 8628 8968
rect 8760 8916 8812 8968
rect 2136 8848 2188 8900
rect 3332 8891 3384 8900
rect 3332 8857 3341 8891
rect 3341 8857 3375 8891
rect 3375 8857 3384 8891
rect 3332 8848 3384 8857
rect 4896 8848 4948 8900
rect 7472 8848 7524 8900
rect 9496 9027 9548 9036
rect 9496 8993 9505 9027
rect 9505 8993 9539 9027
rect 9539 8993 9548 9027
rect 9496 8984 9548 8993
rect 8944 8916 8996 8968
rect 9772 8959 9824 8968
rect 9772 8925 9781 8959
rect 9781 8925 9815 8959
rect 9815 8925 9824 8959
rect 9772 8916 9824 8925
rect 2688 8780 2740 8832
rect 6828 8780 6880 8832
rect 6920 8780 6972 8832
rect 8208 8780 8260 8832
rect 9128 8823 9180 8832
rect 9128 8789 9137 8823
rect 9137 8789 9171 8823
rect 9171 8789 9180 8823
rect 9128 8780 9180 8789
rect 9772 8780 9824 8832
rect 10416 9052 10468 9104
rect 11612 9095 11664 9104
rect 11612 9061 11621 9095
rect 11621 9061 11655 9095
rect 11655 9061 11664 9095
rect 11612 9052 11664 9061
rect 11980 9052 12032 9104
rect 12992 9120 13044 9172
rect 13268 9163 13320 9172
rect 13268 9129 13277 9163
rect 13277 9129 13311 9163
rect 13311 9129 13320 9163
rect 13268 9120 13320 9129
rect 13728 9163 13780 9172
rect 13728 9129 13737 9163
rect 13737 9129 13771 9163
rect 13771 9129 13780 9163
rect 13728 9120 13780 9129
rect 15568 9120 15620 9172
rect 17776 9120 17828 9172
rect 10600 8984 10652 9036
rect 11152 8984 11204 9036
rect 11520 8984 11572 9036
rect 11888 8984 11940 9036
rect 12164 9027 12216 9036
rect 12164 8993 12173 9027
rect 12173 8993 12207 9027
rect 12207 8993 12216 9027
rect 12164 8984 12216 8993
rect 10416 8916 10468 8968
rect 10508 8916 10560 8968
rect 11888 8848 11940 8900
rect 12808 8984 12860 9036
rect 13360 8984 13412 9036
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 13728 8984 13780 9036
rect 15660 9052 15712 9104
rect 18512 9120 18564 9172
rect 18788 9120 18840 9172
rect 14372 9027 14424 9036
rect 14372 8993 14381 9027
rect 14381 8993 14415 9027
rect 14415 8993 14424 9027
rect 14372 8984 14424 8993
rect 14556 8984 14608 9036
rect 13544 8916 13596 8968
rect 14004 8916 14056 8968
rect 15752 8984 15804 9036
rect 13084 8848 13136 8900
rect 15476 8848 15528 8900
rect 16764 9027 16816 9036
rect 21088 9120 21140 9172
rect 21364 9052 21416 9104
rect 16764 8993 16782 9027
rect 16782 8993 16816 9027
rect 16764 8984 16816 8993
rect 18052 9027 18104 9036
rect 17408 8959 17460 8968
rect 10140 8780 10192 8832
rect 12716 8780 12768 8832
rect 14556 8823 14608 8832
rect 14556 8789 14565 8823
rect 14565 8789 14599 8823
rect 14599 8789 14608 8823
rect 14556 8780 14608 8789
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 15200 8823 15252 8832
rect 15200 8789 15209 8823
rect 15209 8789 15243 8823
rect 15243 8789 15252 8823
rect 15200 8780 15252 8789
rect 15660 8823 15712 8832
rect 15660 8789 15669 8823
rect 15669 8789 15703 8823
rect 15703 8789 15712 8823
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 18052 8993 18061 9027
rect 18061 8993 18095 9027
rect 18095 8993 18104 9027
rect 18052 8984 18104 8993
rect 18788 8984 18840 9036
rect 19064 9027 19116 9036
rect 19064 8993 19073 9027
rect 19073 8993 19107 9027
rect 19107 8993 19116 9027
rect 19064 8984 19116 8993
rect 19432 8984 19484 9036
rect 19892 9027 19944 9036
rect 17960 8916 18012 8968
rect 19892 8993 19926 9027
rect 19926 8993 19944 9027
rect 19892 8984 19944 8993
rect 21548 9027 21600 9036
rect 21548 8993 21557 9027
rect 21557 8993 21591 9027
rect 21591 8993 21600 9027
rect 21548 8984 21600 8993
rect 18236 8891 18288 8900
rect 18236 8857 18245 8891
rect 18245 8857 18279 8891
rect 18279 8857 18288 8891
rect 18236 8848 18288 8857
rect 18972 8848 19024 8900
rect 15660 8780 15712 8789
rect 18144 8780 18196 8832
rect 19340 8780 19392 8832
rect 19616 8780 19668 8832
rect 20536 8780 20588 8832
rect 20812 8780 20864 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 1768 8576 1820 8628
rect 1860 8508 1912 8560
rect 1952 8551 2004 8560
rect 1952 8517 1961 8551
rect 1961 8517 1995 8551
rect 1995 8517 2004 8551
rect 4160 8576 4212 8628
rect 4804 8576 4856 8628
rect 5632 8576 5684 8628
rect 6000 8576 6052 8628
rect 8944 8576 8996 8628
rect 10140 8576 10192 8628
rect 10600 8576 10652 8628
rect 1952 8508 2004 8517
rect 6276 8551 6328 8560
rect 6276 8517 6285 8551
rect 6285 8517 6319 8551
rect 6319 8517 6328 8551
rect 6276 8508 6328 8517
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 6184 8440 6236 8492
rect 7104 8483 7156 8492
rect 7104 8449 7113 8483
rect 7113 8449 7147 8483
rect 7147 8449 7156 8483
rect 7104 8440 7156 8449
rect 7196 8440 7248 8492
rect 7380 8440 7432 8492
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 8300 8483 8352 8492
rect 8300 8449 8309 8483
rect 8309 8449 8343 8483
rect 8343 8449 8352 8483
rect 8300 8440 8352 8449
rect 2780 8372 2832 8424
rect 3792 8372 3844 8424
rect 5540 8372 5592 8424
rect 5816 8372 5868 8424
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 7012 8372 7064 8424
rect 9128 8372 9180 8424
rect 9220 8372 9272 8424
rect 9588 8372 9640 8424
rect 10508 8508 10560 8560
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 2136 8279 2188 8288
rect 2136 8245 2145 8279
rect 2145 8245 2179 8279
rect 2179 8245 2188 8279
rect 2136 8236 2188 8245
rect 2872 8304 2924 8356
rect 3056 8304 3108 8356
rect 3332 8304 3384 8356
rect 7104 8304 7156 8356
rect 10048 8304 10100 8356
rect 10876 8576 10928 8628
rect 11060 8576 11112 8628
rect 11244 8576 11296 8628
rect 12532 8576 12584 8628
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 13268 8576 13320 8628
rect 11244 8440 11296 8492
rect 12716 8508 12768 8560
rect 12256 8483 12308 8492
rect 12256 8449 12265 8483
rect 12265 8449 12299 8483
rect 12299 8449 12308 8483
rect 12256 8440 12308 8449
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 15660 8576 15712 8628
rect 15752 8576 15804 8628
rect 17776 8619 17828 8628
rect 16764 8551 16816 8560
rect 16764 8517 16773 8551
rect 16773 8517 16807 8551
rect 16807 8517 16816 8551
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 16764 8508 16816 8517
rect 12164 8415 12216 8424
rect 12164 8381 12173 8415
rect 12173 8381 12207 8415
rect 12207 8381 12216 8415
rect 12164 8372 12216 8381
rect 13728 8372 13780 8424
rect 18052 8508 18104 8560
rect 15476 8372 15528 8424
rect 18972 8440 19024 8492
rect 17684 8372 17736 8424
rect 20168 8576 20220 8628
rect 20904 8576 20956 8628
rect 19892 8483 19944 8492
rect 10876 8304 10928 8356
rect 12440 8304 12492 8356
rect 12808 8304 12860 8356
rect 12900 8304 12952 8356
rect 14832 8304 14884 8356
rect 3424 8236 3476 8288
rect 4896 8236 4948 8288
rect 4988 8236 5040 8288
rect 5448 8236 5500 8288
rect 5816 8279 5868 8288
rect 5816 8245 5825 8279
rect 5825 8245 5859 8279
rect 5859 8245 5868 8279
rect 5816 8236 5868 8245
rect 7288 8279 7340 8288
rect 7288 8245 7297 8279
rect 7297 8245 7331 8279
rect 7331 8245 7340 8279
rect 7288 8236 7340 8245
rect 8392 8279 8444 8288
rect 8392 8245 8401 8279
rect 8401 8245 8435 8279
rect 8435 8245 8444 8279
rect 8392 8236 8444 8245
rect 8944 8279 8996 8288
rect 8944 8245 8953 8279
rect 8953 8245 8987 8279
rect 8987 8245 8996 8279
rect 8944 8236 8996 8245
rect 9312 8236 9364 8288
rect 10140 8279 10192 8288
rect 10140 8245 10149 8279
rect 10149 8245 10183 8279
rect 10183 8245 10192 8279
rect 10140 8236 10192 8245
rect 12164 8236 12216 8288
rect 13360 8279 13412 8288
rect 13360 8245 13369 8279
rect 13369 8245 13403 8279
rect 13403 8245 13412 8279
rect 13360 8236 13412 8245
rect 13728 8236 13780 8288
rect 14004 8236 14056 8288
rect 15844 8304 15896 8356
rect 16028 8304 16080 8356
rect 15936 8236 15988 8288
rect 17132 8304 17184 8356
rect 17592 8304 17644 8356
rect 18328 8304 18380 8356
rect 18420 8236 18472 8288
rect 19892 8449 19901 8483
rect 19901 8449 19935 8483
rect 19935 8449 19944 8483
rect 19892 8440 19944 8449
rect 20720 8440 20772 8492
rect 19340 8372 19392 8424
rect 19708 8372 19760 8424
rect 20536 8372 20588 8424
rect 21180 8372 21232 8424
rect 21548 8415 21600 8424
rect 21548 8381 21557 8415
rect 21557 8381 21591 8415
rect 21591 8381 21600 8415
rect 21548 8372 21600 8381
rect 21088 8304 21140 8356
rect 19984 8279 20036 8288
rect 19984 8245 19993 8279
rect 19993 8245 20027 8279
rect 20027 8245 20036 8279
rect 19984 8236 20036 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 3056 8075 3108 8084
rect 2136 7964 2188 8016
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 2964 7964 3016 8016
rect 1952 7939 2004 7948
rect 1952 7905 1986 7939
rect 1986 7905 2004 7939
rect 4068 7964 4120 8016
rect 5172 8032 5224 8084
rect 6828 8032 6880 8084
rect 7104 8075 7156 8084
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 7288 8032 7340 8084
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 3240 7939 3292 7948
rect 1952 7896 2004 7905
rect 3240 7905 3249 7939
rect 3249 7905 3283 7939
rect 3283 7905 3292 7939
rect 3240 7896 3292 7905
rect 3516 7939 3568 7948
rect 3516 7905 3525 7939
rect 3525 7905 3559 7939
rect 3559 7905 3568 7939
rect 3516 7896 3568 7905
rect 4252 7939 4304 7948
rect 4252 7905 4261 7939
rect 4261 7905 4295 7939
rect 4295 7905 4304 7939
rect 4252 7896 4304 7905
rect 4160 7828 4212 7880
rect 4896 7896 4948 7948
rect 5632 7964 5684 8016
rect 7748 7964 7800 8016
rect 8392 8032 8444 8084
rect 8944 8032 8996 8084
rect 9956 8032 10008 8084
rect 10784 8032 10836 8084
rect 10968 8075 11020 8084
rect 10968 8041 10977 8075
rect 10977 8041 11011 8075
rect 11011 8041 11020 8075
rect 10968 8032 11020 8041
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 2872 7760 2924 7812
rect 3332 7692 3384 7744
rect 3424 7692 3476 7744
rect 3976 7692 4028 7744
rect 6828 7692 6880 7744
rect 8576 7939 8628 7948
rect 8576 7905 8585 7939
rect 8585 7905 8619 7939
rect 8619 7905 8628 7939
rect 8576 7896 8628 7905
rect 9220 7964 9272 8016
rect 9588 7964 9640 8016
rect 10416 7964 10468 8016
rect 10600 7964 10652 8016
rect 7472 7828 7524 7880
rect 12164 8032 12216 8084
rect 13360 8032 13412 8084
rect 13728 8032 13780 8084
rect 15568 8032 15620 8084
rect 7748 7692 7800 7744
rect 10416 7828 10468 7880
rect 12256 7896 12308 7948
rect 12624 7964 12676 8016
rect 15108 7964 15160 8016
rect 15292 7964 15344 8016
rect 19340 8032 19392 8084
rect 19984 8032 20036 8084
rect 21548 8075 21600 8084
rect 21548 8041 21557 8075
rect 21557 8041 21591 8075
rect 21591 8041 21600 8075
rect 21548 8032 21600 8041
rect 17592 7964 17644 8016
rect 13176 7896 13228 7948
rect 13268 7896 13320 7948
rect 13820 7939 13872 7948
rect 13820 7905 13829 7939
rect 13829 7905 13863 7939
rect 13863 7905 13872 7939
rect 13820 7896 13872 7905
rect 14740 7939 14792 7948
rect 14740 7905 14749 7939
rect 14749 7905 14783 7939
rect 14783 7905 14792 7939
rect 14740 7896 14792 7905
rect 12808 7828 12860 7880
rect 12440 7803 12492 7812
rect 12440 7769 12449 7803
rect 12449 7769 12483 7803
rect 12483 7769 12492 7803
rect 13084 7828 13136 7880
rect 13728 7828 13780 7880
rect 14004 7871 14056 7880
rect 14004 7837 14013 7871
rect 14013 7837 14047 7871
rect 14047 7837 14056 7871
rect 14004 7828 14056 7837
rect 15752 7896 15804 7948
rect 16580 7896 16632 7948
rect 15660 7828 15712 7880
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 16764 7828 16816 7880
rect 19708 7896 19760 7948
rect 17960 7871 18012 7880
rect 12440 7760 12492 7769
rect 9772 7692 9824 7744
rect 10600 7735 10652 7744
rect 10600 7701 10609 7735
rect 10609 7701 10643 7735
rect 10643 7701 10652 7735
rect 15844 7760 15896 7812
rect 10600 7692 10652 7701
rect 13084 7692 13136 7744
rect 13360 7692 13412 7744
rect 13912 7692 13964 7744
rect 15200 7692 15252 7744
rect 16028 7692 16080 7744
rect 16396 7692 16448 7744
rect 16764 7692 16816 7744
rect 17408 7760 17460 7812
rect 17960 7837 17969 7871
rect 17969 7837 18003 7871
rect 18003 7837 18012 7871
rect 17960 7828 18012 7837
rect 18972 7828 19024 7880
rect 20168 7896 20220 7948
rect 20536 7896 20588 7948
rect 20444 7828 20496 7880
rect 20812 7828 20864 7880
rect 20720 7760 20772 7812
rect 21272 7828 21324 7880
rect 19892 7692 19944 7744
rect 20444 7735 20496 7744
rect 20444 7701 20453 7735
rect 20453 7701 20487 7735
rect 20487 7701 20496 7735
rect 20444 7692 20496 7701
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 1952 7488 2004 7540
rect 2872 7488 2924 7540
rect 3424 7488 3476 7540
rect 3792 7488 3844 7540
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 4160 7488 4212 7497
rect 4988 7531 5040 7540
rect 4988 7497 4997 7531
rect 4997 7497 5031 7531
rect 5031 7497 5040 7531
rect 4988 7488 5040 7497
rect 5080 7488 5132 7540
rect 6736 7488 6788 7540
rect 8392 7488 8444 7540
rect 8576 7488 8628 7540
rect 1492 7327 1544 7336
rect 1492 7293 1501 7327
rect 1501 7293 1535 7327
rect 1535 7293 1544 7327
rect 4068 7352 4120 7404
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 5356 7352 5408 7404
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 9220 7420 9272 7472
rect 7104 7352 7156 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 9312 7352 9364 7404
rect 1492 7284 1544 7293
rect 3332 7284 3384 7336
rect 4160 7284 4212 7336
rect 6092 7284 6144 7336
rect 2872 7216 2924 7268
rect 4068 7216 4120 7268
rect 5908 7216 5960 7268
rect 3240 7148 3292 7200
rect 3332 7148 3384 7200
rect 3700 7191 3752 7200
rect 3700 7157 3709 7191
rect 3709 7157 3743 7191
rect 3743 7157 3752 7191
rect 3700 7148 3752 7157
rect 4528 7191 4580 7200
rect 4528 7157 4537 7191
rect 4537 7157 4571 7191
rect 4571 7157 4580 7191
rect 4528 7148 4580 7157
rect 4620 7148 4672 7200
rect 5540 7148 5592 7200
rect 5632 7148 5684 7200
rect 6276 7148 6328 7200
rect 7012 7216 7064 7268
rect 10232 7488 10284 7540
rect 9956 7420 10008 7472
rect 11244 7420 11296 7472
rect 13360 7420 13412 7472
rect 13544 7420 13596 7472
rect 12900 7352 12952 7404
rect 13084 7352 13136 7404
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 15108 7420 15160 7472
rect 17776 7420 17828 7472
rect 19064 7488 19116 7540
rect 19248 7488 19300 7540
rect 19432 7488 19484 7540
rect 18512 7420 18564 7472
rect 19984 7420 20036 7472
rect 16396 7352 16448 7404
rect 17132 7395 17184 7404
rect 17132 7361 17141 7395
rect 17141 7361 17175 7395
rect 17175 7361 17184 7395
rect 17132 7352 17184 7361
rect 18972 7352 19024 7404
rect 21824 7420 21876 7472
rect 12440 7284 12492 7336
rect 10416 7216 10468 7268
rect 10968 7216 11020 7268
rect 13544 7284 13596 7336
rect 13912 7284 13964 7336
rect 14096 7284 14148 7336
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 17592 7327 17644 7336
rect 17592 7293 17601 7327
rect 17601 7293 17635 7327
rect 17635 7293 17644 7327
rect 17592 7284 17644 7293
rect 17776 7284 17828 7336
rect 20720 7352 20772 7404
rect 19248 7284 19300 7336
rect 19524 7284 19576 7336
rect 19708 7284 19760 7336
rect 21548 7327 21600 7336
rect 21548 7293 21557 7327
rect 21557 7293 21591 7327
rect 21591 7293 21600 7327
rect 21548 7284 21600 7293
rect 7472 7191 7524 7200
rect 7472 7157 7481 7191
rect 7481 7157 7515 7191
rect 7515 7157 7524 7191
rect 7472 7148 7524 7157
rect 10324 7191 10376 7200
rect 10324 7157 10333 7191
rect 10333 7157 10367 7191
rect 10367 7157 10376 7191
rect 10324 7148 10376 7157
rect 10600 7191 10652 7200
rect 10600 7157 10609 7191
rect 10609 7157 10643 7191
rect 10643 7157 10652 7191
rect 10600 7148 10652 7157
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11428 7191 11480 7200
rect 11152 7148 11204 7157
rect 11428 7157 11437 7191
rect 11437 7157 11471 7191
rect 11471 7157 11480 7191
rect 11428 7148 11480 7157
rect 11520 7148 11572 7200
rect 13636 7216 13688 7268
rect 16948 7216 17000 7268
rect 12900 7148 12952 7200
rect 13360 7191 13412 7200
rect 13360 7157 13369 7191
rect 13369 7157 13403 7191
rect 13403 7157 13412 7191
rect 13360 7148 13412 7157
rect 14188 7191 14240 7200
rect 14188 7157 14197 7191
rect 14197 7157 14231 7191
rect 14231 7157 14240 7191
rect 14188 7148 14240 7157
rect 14372 7148 14424 7200
rect 15292 7148 15344 7200
rect 15660 7191 15712 7200
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 16120 7148 16172 7157
rect 17960 7216 18012 7268
rect 17684 7148 17736 7200
rect 19064 7216 19116 7268
rect 18328 7191 18380 7200
rect 18328 7157 18337 7191
rect 18337 7157 18371 7191
rect 18371 7157 18380 7191
rect 18328 7148 18380 7157
rect 18604 7148 18656 7200
rect 18788 7148 18840 7200
rect 19524 7148 19576 7200
rect 20168 7148 20220 7200
rect 20904 7191 20956 7200
rect 20904 7157 20913 7191
rect 20913 7157 20947 7191
rect 20947 7157 20956 7191
rect 20904 7148 20956 7157
rect 21456 7148 21508 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 3148 6987 3200 6996
rect 1676 6919 1728 6928
rect 1676 6885 1685 6919
rect 1685 6885 1719 6919
rect 1719 6885 1728 6919
rect 1676 6876 1728 6885
rect 3148 6953 3157 6987
rect 3157 6953 3191 6987
rect 3191 6953 3200 6987
rect 3148 6944 3200 6953
rect 4344 6944 4396 6996
rect 4528 6944 4580 6996
rect 6092 6987 6144 6996
rect 3332 6876 3384 6928
rect 3516 6876 3568 6928
rect 4160 6876 4212 6928
rect 6092 6953 6101 6987
rect 6101 6953 6135 6987
rect 6135 6953 6144 6987
rect 6092 6944 6144 6953
rect 6736 6944 6788 6996
rect 8208 6944 8260 6996
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 1400 6604 1452 6656
rect 2964 6740 3016 6792
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 4712 6808 4764 6860
rect 8576 6876 8628 6928
rect 9220 6944 9272 6996
rect 10324 6987 10376 6996
rect 10324 6953 10333 6987
rect 10333 6953 10367 6987
rect 10367 6953 10376 6987
rect 10324 6944 10376 6953
rect 12256 6944 12308 6996
rect 12440 6944 12492 6996
rect 13176 6944 13228 6996
rect 13360 6944 13412 6996
rect 14096 6987 14148 6996
rect 14096 6953 14105 6987
rect 14105 6953 14139 6987
rect 14139 6953 14148 6987
rect 14096 6944 14148 6953
rect 11152 6876 11204 6928
rect 12348 6876 12400 6928
rect 12992 6876 13044 6928
rect 5540 6851 5592 6860
rect 5540 6817 5557 6851
rect 5557 6817 5591 6851
rect 5591 6817 5592 6851
rect 5540 6808 5592 6817
rect 6092 6808 6144 6860
rect 9864 6808 9916 6860
rect 10324 6808 10376 6860
rect 10968 6808 11020 6860
rect 12900 6851 12952 6860
rect 12900 6817 12918 6851
rect 12918 6817 12952 6851
rect 13544 6876 13596 6928
rect 12900 6808 12952 6817
rect 3148 6672 3200 6724
rect 2228 6604 2280 6656
rect 3056 6604 3108 6656
rect 3792 6604 3844 6656
rect 4068 6604 4120 6656
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 7104 6740 7156 6792
rect 7656 6740 7708 6792
rect 8392 6740 8444 6792
rect 9312 6740 9364 6792
rect 9680 6740 9732 6792
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 11152 6783 11204 6792
rect 11152 6749 11161 6783
rect 11161 6749 11195 6783
rect 11195 6749 11204 6783
rect 13176 6783 13228 6792
rect 11152 6740 11204 6749
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 5365 6715 5417 6724
rect 5365 6681 5399 6715
rect 5399 6681 5417 6715
rect 5365 6672 5417 6681
rect 6736 6672 6788 6724
rect 8484 6715 8536 6724
rect 8484 6681 8493 6715
rect 8493 6681 8527 6715
rect 8527 6681 8536 6715
rect 8484 6672 8536 6681
rect 15476 6919 15528 6928
rect 15476 6885 15485 6919
rect 15485 6885 15519 6919
rect 15519 6885 15528 6919
rect 15476 6876 15528 6885
rect 16120 6944 16172 6996
rect 16948 6987 17000 6996
rect 16948 6953 16957 6987
rect 16957 6953 16991 6987
rect 16991 6953 17000 6987
rect 16948 6944 17000 6953
rect 17316 6944 17368 6996
rect 14556 6851 14608 6860
rect 14556 6817 14565 6851
rect 14565 6817 14599 6851
rect 14599 6817 14608 6851
rect 14556 6808 14608 6817
rect 18328 6944 18380 6996
rect 20168 6987 20220 6996
rect 20168 6953 20177 6987
rect 20177 6953 20211 6987
rect 20211 6953 20220 6987
rect 20168 6944 20220 6953
rect 20444 6944 20496 6996
rect 21548 6987 21600 6996
rect 21548 6953 21557 6987
rect 21557 6953 21591 6987
rect 21591 6953 21600 6987
rect 21548 6944 21600 6953
rect 20812 6876 20864 6928
rect 17316 6851 17368 6860
rect 17316 6817 17325 6851
rect 17325 6817 17359 6851
rect 17359 6817 17368 6851
rect 17316 6808 17368 6817
rect 18052 6808 18104 6860
rect 18420 6851 18472 6860
rect 18420 6817 18429 6851
rect 18429 6817 18463 6851
rect 18463 6817 18472 6851
rect 18420 6808 18472 6817
rect 19248 6808 19300 6860
rect 19984 6808 20036 6860
rect 21088 6851 21140 6860
rect 5540 6604 5592 6656
rect 5816 6604 5868 6656
rect 7104 6604 7156 6656
rect 7840 6604 7892 6656
rect 8208 6604 8260 6656
rect 9404 6647 9456 6656
rect 9404 6613 9413 6647
rect 9413 6613 9447 6647
rect 9447 6613 9456 6647
rect 9404 6604 9456 6613
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9956 6647 10008 6656
rect 9680 6604 9732 6613
rect 9956 6613 9965 6647
rect 9965 6613 9999 6647
rect 9999 6613 10008 6647
rect 9956 6604 10008 6613
rect 10324 6604 10376 6656
rect 10692 6604 10744 6656
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 11796 6647 11848 6656
rect 11796 6613 11805 6647
rect 11805 6613 11839 6647
rect 11839 6613 11848 6647
rect 11796 6604 11848 6613
rect 12808 6604 12860 6656
rect 13544 6604 13596 6656
rect 13912 6672 13964 6724
rect 14740 6672 14792 6724
rect 15752 6740 15804 6792
rect 16120 6740 16172 6792
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 17500 6783 17552 6792
rect 16672 6740 16724 6749
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 17592 6740 17644 6792
rect 18144 6783 18196 6792
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 18972 6740 19024 6792
rect 19892 6783 19944 6792
rect 19892 6749 19901 6783
rect 19901 6749 19935 6783
rect 19935 6749 19944 6783
rect 21088 6817 21097 6851
rect 21097 6817 21131 6851
rect 21131 6817 21140 6851
rect 21088 6808 21140 6817
rect 19892 6740 19944 6749
rect 18512 6672 18564 6724
rect 14556 6604 14608 6656
rect 14832 6604 14884 6656
rect 15568 6604 15620 6656
rect 16028 6604 16080 6656
rect 16212 6604 16264 6656
rect 17684 6604 17736 6656
rect 20444 6672 20496 6724
rect 20996 6672 21048 6724
rect 20168 6604 20220 6656
rect 20260 6604 20312 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 1952 6443 2004 6452
rect 1952 6409 1961 6443
rect 1961 6409 1995 6443
rect 1995 6409 2004 6443
rect 1952 6400 2004 6409
rect 3700 6400 3752 6452
rect 4252 6400 4304 6452
rect 5172 6400 5224 6452
rect 5724 6400 5776 6452
rect 6736 6400 6788 6452
rect 6828 6400 6880 6452
rect 2412 6332 2464 6384
rect 2872 6332 2924 6384
rect 3792 6332 3844 6384
rect 2228 6307 2280 6316
rect 2228 6273 2237 6307
rect 2237 6273 2271 6307
rect 2271 6273 2280 6307
rect 2228 6264 2280 6273
rect 2688 6264 2740 6316
rect 4436 6332 4488 6384
rect 4804 6332 4856 6384
rect 1768 6239 1820 6248
rect 1216 6128 1268 6180
rect 1768 6205 1777 6239
rect 1777 6205 1811 6239
rect 1811 6205 1820 6239
rect 1768 6196 1820 6205
rect 4068 6196 4120 6248
rect 4252 6196 4304 6248
rect 3516 6128 3568 6180
rect 4988 6264 5040 6316
rect 5540 6264 5592 6316
rect 6644 6264 6696 6316
rect 7380 6400 7432 6452
rect 7288 6332 7340 6384
rect 7840 6332 7892 6384
rect 7196 6264 7248 6316
rect 7472 6264 7524 6316
rect 7288 6196 7340 6248
rect 7748 6196 7800 6248
rect 4804 6128 4856 6180
rect 5080 6128 5132 6180
rect 5172 6128 5224 6180
rect 9496 6400 9548 6452
rect 8668 6332 8720 6384
rect 9680 6332 9732 6384
rect 10968 6400 11020 6452
rect 11060 6332 11112 6384
rect 11244 6400 11296 6452
rect 12256 6443 12308 6452
rect 8576 6264 8628 6316
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 9956 6239 10008 6248
rect 2504 6060 2556 6112
rect 2688 6060 2740 6112
rect 2964 6060 3016 6112
rect 3332 6103 3384 6112
rect 3332 6069 3341 6103
rect 3341 6069 3375 6103
rect 3375 6069 3384 6103
rect 3332 6060 3384 6069
rect 3700 6103 3752 6112
rect 3700 6069 3709 6103
rect 3709 6069 3743 6103
rect 3743 6069 3752 6103
rect 3700 6060 3752 6069
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 5816 6103 5868 6112
rect 3792 6060 3844 6069
rect 5816 6069 5825 6103
rect 5825 6069 5859 6103
rect 5859 6069 5868 6103
rect 5816 6060 5868 6069
rect 6552 6060 6604 6112
rect 8944 6128 8996 6180
rect 9312 6171 9364 6180
rect 9312 6137 9321 6171
rect 9321 6137 9355 6171
rect 9355 6137 9364 6171
rect 9312 6128 9364 6137
rect 9956 6205 9965 6239
rect 9965 6205 9999 6239
rect 9999 6205 10008 6239
rect 9956 6196 10008 6205
rect 11336 6264 11388 6316
rect 12256 6409 12265 6443
rect 12265 6409 12299 6443
rect 12299 6409 12308 6443
rect 12256 6400 12308 6409
rect 12348 6400 12400 6452
rect 13176 6400 13228 6452
rect 22008 6443 22060 6452
rect 22008 6409 22017 6443
rect 22017 6409 22051 6443
rect 22051 6409 22060 6443
rect 22008 6400 22060 6409
rect 12256 6264 12308 6316
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 12900 6332 12952 6384
rect 13912 6375 13964 6384
rect 13544 6307 13596 6316
rect 13544 6273 13553 6307
rect 13553 6273 13587 6307
rect 13587 6273 13596 6307
rect 13544 6264 13596 6273
rect 13912 6341 13921 6375
rect 13921 6341 13955 6375
rect 13955 6341 13964 6375
rect 13912 6332 13964 6341
rect 14096 6332 14148 6384
rect 14280 6307 14332 6316
rect 14280 6273 14289 6307
rect 14289 6273 14323 6307
rect 14323 6273 14332 6307
rect 14280 6264 14332 6273
rect 14832 6264 14884 6316
rect 15752 6264 15804 6316
rect 19156 6332 19208 6384
rect 20720 6332 20772 6384
rect 17316 6264 17368 6316
rect 17500 6307 17552 6316
rect 17500 6273 17509 6307
rect 17509 6273 17543 6307
rect 17543 6273 17552 6307
rect 17500 6264 17552 6273
rect 17868 6307 17920 6316
rect 17868 6273 17877 6307
rect 17877 6273 17911 6307
rect 17911 6273 17920 6307
rect 17868 6264 17920 6273
rect 18052 6264 18104 6316
rect 18880 6264 18932 6316
rect 19248 6307 19300 6316
rect 19248 6273 19257 6307
rect 19257 6273 19291 6307
rect 19291 6273 19300 6307
rect 19248 6264 19300 6273
rect 11520 6196 11572 6248
rect 13360 6196 13412 6248
rect 14188 6196 14240 6248
rect 14556 6239 14608 6248
rect 14556 6205 14565 6239
rect 14565 6205 14599 6239
rect 14599 6205 14608 6239
rect 14556 6196 14608 6205
rect 15476 6239 15528 6248
rect 8392 6103 8444 6112
rect 8392 6069 8401 6103
rect 8401 6069 8435 6103
rect 8435 6069 8444 6103
rect 8392 6060 8444 6069
rect 9128 6060 9180 6112
rect 9404 6103 9456 6112
rect 9404 6069 9413 6103
rect 9413 6069 9447 6103
rect 9447 6069 9456 6103
rect 9404 6060 9456 6069
rect 9864 6103 9916 6112
rect 9864 6069 9873 6103
rect 9873 6069 9907 6103
rect 9907 6069 9916 6103
rect 9864 6060 9916 6069
rect 11244 6128 11296 6180
rect 12624 6171 12676 6180
rect 10600 6060 10652 6112
rect 10968 6060 11020 6112
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 11428 6103 11480 6112
rect 11428 6069 11437 6103
rect 11437 6069 11471 6103
rect 11471 6069 11480 6103
rect 11428 6060 11480 6069
rect 11612 6060 11664 6112
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 12624 6137 12633 6171
rect 12633 6137 12667 6171
rect 12667 6137 12676 6171
rect 12624 6128 12676 6137
rect 12808 6128 12860 6180
rect 15476 6205 15485 6239
rect 15485 6205 15519 6239
rect 15519 6205 15528 6239
rect 15476 6196 15528 6205
rect 16028 6239 16080 6248
rect 16028 6205 16037 6239
rect 16037 6205 16071 6239
rect 16071 6205 16080 6239
rect 16028 6196 16080 6205
rect 18144 6196 18196 6248
rect 14832 6128 14884 6180
rect 14004 6060 14056 6112
rect 14372 6060 14424 6112
rect 17960 6128 18012 6180
rect 15384 6060 15436 6112
rect 16764 6060 16816 6112
rect 16948 6103 17000 6112
rect 16948 6069 16957 6103
rect 16957 6069 16991 6103
rect 16991 6069 17000 6103
rect 16948 6060 17000 6069
rect 17040 6060 17092 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 17684 6060 17736 6112
rect 18788 6103 18840 6112
rect 18788 6069 18797 6103
rect 18797 6069 18831 6103
rect 18831 6069 18840 6103
rect 18788 6060 18840 6069
rect 18972 6103 19024 6112
rect 18972 6069 18981 6103
rect 18981 6069 19015 6103
rect 19015 6069 19024 6103
rect 18972 6060 19024 6069
rect 20168 6128 20220 6180
rect 21088 6171 21140 6180
rect 21088 6137 21097 6171
rect 21097 6137 21131 6171
rect 21131 6137 21140 6171
rect 21088 6128 21140 6137
rect 21548 6128 21600 6180
rect 19984 6060 20036 6112
rect 20720 6060 20772 6112
rect 21180 6060 21232 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 2872 5856 2924 5908
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 3700 5856 3752 5908
rect 3976 5856 4028 5908
rect 5448 5856 5500 5908
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 5816 5856 5868 5908
rect 6736 5899 6788 5908
rect 6736 5865 6745 5899
rect 6745 5865 6779 5899
rect 6779 5865 6788 5899
rect 6736 5856 6788 5865
rect 1952 5788 2004 5840
rect 1308 5720 1360 5772
rect 7932 5788 7984 5840
rect 3240 5720 3292 5772
rect 3976 5720 4028 5772
rect 3148 5652 3200 5704
rect 4252 5720 4304 5772
rect 4804 5720 4856 5772
rect 5724 5720 5776 5772
rect 6184 5720 6236 5772
rect 7288 5720 7340 5772
rect 8024 5720 8076 5772
rect 8944 5788 8996 5840
rect 10324 5788 10376 5840
rect 10968 5856 11020 5908
rect 12348 5856 12400 5908
rect 12440 5856 12492 5908
rect 11244 5831 11296 5840
rect 11244 5797 11253 5831
rect 11253 5797 11287 5831
rect 11287 5797 11296 5831
rect 11244 5788 11296 5797
rect 11796 5788 11848 5840
rect 12900 5788 12952 5840
rect 13820 5788 13872 5840
rect 10508 5763 10560 5772
rect 10508 5729 10526 5763
rect 10526 5729 10560 5763
rect 10508 5720 10560 5729
rect 6828 5652 6880 5704
rect 2688 5516 2740 5568
rect 3700 5516 3752 5568
rect 3792 5516 3844 5568
rect 5172 5516 5224 5568
rect 5816 5516 5868 5568
rect 6184 5559 6236 5568
rect 6184 5525 6193 5559
rect 6193 5525 6227 5559
rect 6227 5525 6236 5559
rect 6184 5516 6236 5525
rect 6920 5516 6972 5568
rect 7656 5516 7708 5568
rect 8208 5516 8260 5568
rect 8576 5652 8628 5704
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 11612 5720 11664 5772
rect 11888 5720 11940 5772
rect 12348 5720 12400 5772
rect 13268 5720 13320 5772
rect 15476 5856 15528 5908
rect 17040 5856 17092 5908
rect 17408 5899 17460 5908
rect 17408 5865 17417 5899
rect 17417 5865 17451 5899
rect 17451 5865 17460 5899
rect 17408 5856 17460 5865
rect 18144 5856 18196 5908
rect 14280 5788 14332 5840
rect 8668 5584 8720 5636
rect 9772 5584 9824 5636
rect 11244 5584 11296 5636
rect 8484 5516 8536 5568
rect 9496 5516 9548 5568
rect 14004 5652 14056 5704
rect 11796 5584 11848 5636
rect 12072 5584 12124 5636
rect 12532 5584 12584 5636
rect 12256 5516 12308 5568
rect 12808 5516 12860 5568
rect 14096 5584 14148 5636
rect 15752 5627 15804 5636
rect 15752 5593 15761 5627
rect 15761 5593 15795 5627
rect 15795 5593 15804 5627
rect 15752 5584 15804 5593
rect 16672 5720 16724 5772
rect 16212 5652 16264 5704
rect 16856 5720 16908 5772
rect 17224 5720 17276 5772
rect 19984 5856 20036 5908
rect 20076 5856 20128 5908
rect 20628 5899 20680 5908
rect 20628 5865 20637 5899
rect 20637 5865 20671 5899
rect 20671 5865 20680 5899
rect 20628 5856 20680 5865
rect 19064 5788 19116 5840
rect 19156 5763 19208 5772
rect 19156 5729 19174 5763
rect 19174 5729 19208 5763
rect 19156 5720 19208 5729
rect 19432 5695 19484 5704
rect 19432 5661 19441 5695
rect 19441 5661 19475 5695
rect 19475 5661 19484 5695
rect 19432 5652 19484 5661
rect 17776 5584 17828 5636
rect 18144 5584 18196 5636
rect 13912 5559 13964 5568
rect 13912 5525 13921 5559
rect 13921 5525 13955 5559
rect 13955 5525 13964 5559
rect 13912 5516 13964 5525
rect 19984 5652 20036 5704
rect 20168 5584 20220 5636
rect 20076 5559 20128 5568
rect 20076 5525 20085 5559
rect 20085 5525 20119 5559
rect 20119 5525 20128 5559
rect 20076 5516 20128 5525
rect 21456 5763 21508 5772
rect 21456 5729 21465 5763
rect 21465 5729 21499 5763
rect 21499 5729 21508 5763
rect 21456 5720 21508 5729
rect 20444 5584 20496 5636
rect 21548 5516 21600 5568
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 1768 5312 1820 5364
rect 3792 5312 3844 5364
rect 4068 5355 4120 5364
rect 4068 5321 4077 5355
rect 4077 5321 4111 5355
rect 4111 5321 4120 5355
rect 4068 5312 4120 5321
rect 1952 5176 2004 5228
rect 2688 5219 2740 5228
rect 2688 5185 2697 5219
rect 2697 5185 2731 5219
rect 2731 5185 2740 5219
rect 2688 5176 2740 5185
rect 1308 5108 1360 5160
rect 3516 5108 3568 5160
rect 2872 5040 2924 5092
rect 3976 5176 4028 5228
rect 6920 5312 6972 5364
rect 4804 5219 4856 5228
rect 4804 5185 4813 5219
rect 4813 5185 4847 5219
rect 4847 5185 4856 5219
rect 4804 5176 4856 5185
rect 4988 5176 5040 5228
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 2320 4972 2372 4981
rect 2504 4972 2556 5024
rect 4252 5108 4304 5160
rect 5080 5108 5132 5160
rect 5264 5176 5316 5228
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 5908 5108 5960 5160
rect 7012 5219 7064 5228
rect 7012 5185 7021 5219
rect 7021 5185 7055 5219
rect 7055 5185 7064 5219
rect 7012 5176 7064 5185
rect 7564 5176 7616 5228
rect 8024 5151 8076 5160
rect 8024 5117 8033 5151
rect 8033 5117 8067 5151
rect 8067 5117 8076 5151
rect 8024 5108 8076 5117
rect 8208 5219 8260 5228
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 10416 5312 10468 5364
rect 8208 5176 8260 5185
rect 8668 5108 8720 5160
rect 8944 5108 8996 5160
rect 9220 5108 9272 5160
rect 9772 5108 9824 5160
rect 10692 5108 10744 5160
rect 3884 5040 3936 5092
rect 6184 5040 6236 5092
rect 3976 4972 4028 5024
rect 4712 4972 4764 5024
rect 5080 4972 5132 5024
rect 5448 5015 5500 5024
rect 5448 4981 5457 5015
rect 5457 4981 5491 5015
rect 5491 4981 5500 5015
rect 5448 4972 5500 4981
rect 7472 5040 7524 5092
rect 6736 4972 6788 5024
rect 6828 4972 6880 5024
rect 7196 5015 7248 5024
rect 7196 4981 7205 5015
rect 7205 4981 7239 5015
rect 7239 4981 7248 5015
rect 9128 5040 9180 5092
rect 11152 5176 11204 5228
rect 13176 5244 13228 5296
rect 12256 5176 12308 5228
rect 11060 5151 11112 5160
rect 11060 5117 11069 5151
rect 11069 5117 11103 5151
rect 11103 5117 11112 5151
rect 11060 5108 11112 5117
rect 11888 5108 11940 5160
rect 12808 5219 12860 5228
rect 12808 5185 12817 5219
rect 12817 5185 12851 5219
rect 12851 5185 12860 5219
rect 12808 5176 12860 5185
rect 13084 5176 13136 5228
rect 13544 5176 13596 5228
rect 13912 5219 13964 5228
rect 13912 5185 13921 5219
rect 13921 5185 13955 5219
rect 13955 5185 13964 5219
rect 13912 5176 13964 5185
rect 7196 4972 7248 4981
rect 7748 4972 7800 5024
rect 8300 4972 8352 5024
rect 8576 4972 8628 5024
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 12532 5040 12584 5092
rect 13820 5108 13872 5160
rect 14740 5312 14792 5364
rect 14280 5219 14332 5228
rect 14280 5185 14289 5219
rect 14289 5185 14323 5219
rect 14323 5185 14332 5219
rect 14280 5176 14332 5185
rect 15660 5312 15712 5364
rect 16396 5355 16448 5364
rect 16396 5321 16405 5355
rect 16405 5321 16439 5355
rect 16439 5321 16448 5355
rect 16396 5312 16448 5321
rect 17684 5355 17736 5364
rect 17684 5321 17693 5355
rect 17693 5321 17727 5355
rect 17727 5321 17736 5355
rect 17684 5312 17736 5321
rect 19248 5312 19300 5364
rect 19340 5312 19392 5364
rect 16396 5176 16448 5228
rect 18052 5219 18104 5228
rect 18052 5185 18061 5219
rect 18061 5185 18095 5219
rect 18095 5185 18104 5219
rect 18052 5176 18104 5185
rect 19616 5312 19668 5364
rect 20168 5312 20220 5364
rect 20444 5312 20496 5364
rect 19524 5244 19576 5296
rect 20812 5312 20864 5364
rect 21916 5312 21968 5364
rect 22284 5244 22336 5296
rect 21272 5219 21324 5228
rect 15752 5108 15804 5160
rect 16948 5108 17000 5160
rect 18788 5108 18840 5160
rect 20812 5108 20864 5160
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 21088 5108 21140 5160
rect 21732 5108 21784 5160
rect 13912 5040 13964 5092
rect 14740 5040 14792 5092
rect 16764 5040 16816 5092
rect 18236 5040 18288 5092
rect 18420 5040 18472 5092
rect 20076 5040 20128 5092
rect 21456 5083 21508 5092
rect 21456 5049 21465 5083
rect 21465 5049 21499 5083
rect 21499 5049 21508 5083
rect 21456 5040 21508 5049
rect 9220 4972 9272 4981
rect 11612 4972 11664 5024
rect 11888 4972 11940 5024
rect 12348 4972 12400 5024
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 13360 5015 13412 5024
rect 13360 4981 13369 5015
rect 13369 4981 13403 5015
rect 13403 4981 13412 5015
rect 13360 4972 13412 4981
rect 13544 4972 13596 5024
rect 13820 5015 13872 5024
rect 13820 4981 13829 5015
rect 13829 4981 13863 5015
rect 13863 4981 13872 5015
rect 13820 4972 13872 4981
rect 14096 4972 14148 5024
rect 14372 4972 14424 5024
rect 17040 4972 17092 5024
rect 17316 4972 17368 5024
rect 18144 4972 18196 5024
rect 18788 4972 18840 5024
rect 20168 4972 20220 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 1952 4768 2004 4820
rect 2320 4768 2372 4820
rect 6276 4768 6328 4820
rect 7288 4811 7340 4820
rect 7288 4777 7297 4811
rect 7297 4777 7331 4811
rect 7331 4777 7340 4811
rect 7288 4768 7340 4777
rect 7748 4811 7800 4820
rect 7748 4777 7757 4811
rect 7757 4777 7791 4811
rect 7791 4777 7800 4811
rect 7748 4768 7800 4777
rect 9680 4768 9732 4820
rect 9864 4768 9916 4820
rect 13084 4768 13136 4820
rect 13176 4768 13228 4820
rect 17224 4768 17276 4820
rect 17868 4768 17920 4820
rect 18420 4768 18472 4820
rect 18788 4811 18840 4820
rect 18788 4777 18797 4811
rect 18797 4777 18831 4811
rect 18831 4777 18840 4811
rect 18788 4768 18840 4777
rect 18880 4768 18932 4820
rect 19064 4768 19116 4820
rect 3056 4700 3108 4752
rect 2688 4632 2740 4684
rect 5632 4700 5684 4752
rect 3424 4607 3476 4616
rect 2596 4428 2648 4480
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 4712 4632 4764 4684
rect 5816 4632 5868 4684
rect 7104 4675 7156 4684
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 7656 4700 7708 4752
rect 9220 4700 9272 4752
rect 9128 4675 9180 4684
rect 9128 4641 9137 4675
rect 9137 4641 9171 4675
rect 9171 4641 9180 4675
rect 9128 4632 9180 4641
rect 10508 4700 10560 4752
rect 11612 4700 11664 4752
rect 4344 4564 4396 4616
rect 5264 4607 5316 4616
rect 5264 4573 5273 4607
rect 5273 4573 5307 4607
rect 5307 4573 5316 4607
rect 5264 4564 5316 4573
rect 3056 4496 3108 4548
rect 4988 4496 5040 4548
rect 3792 4428 3844 4480
rect 4252 4428 4304 4480
rect 5724 4428 5776 4480
rect 6736 4428 6788 4480
rect 7288 4564 7340 4616
rect 7380 4564 7432 4616
rect 8208 4564 8260 4616
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 9496 4564 9548 4616
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 10784 4564 10836 4616
rect 11060 4564 11112 4616
rect 11244 4564 11296 4616
rect 11888 4632 11940 4684
rect 12072 4675 12124 4684
rect 12072 4641 12081 4675
rect 12081 4641 12115 4675
rect 12115 4641 12124 4675
rect 12072 4632 12124 4641
rect 12256 4632 12308 4684
rect 12440 4632 12492 4684
rect 13820 4675 13872 4684
rect 13820 4641 13838 4675
rect 13838 4641 13872 4675
rect 13820 4632 13872 4641
rect 14004 4632 14056 4684
rect 14556 4632 14608 4684
rect 12164 4564 12216 4616
rect 14372 4564 14424 4616
rect 15660 4632 15712 4684
rect 16396 4700 16448 4752
rect 19984 4768 20036 4820
rect 20260 4768 20312 4820
rect 20720 4811 20772 4820
rect 20720 4777 20729 4811
rect 20729 4777 20763 4811
rect 20763 4777 20772 4811
rect 20720 4768 20772 4777
rect 21824 4768 21876 4820
rect 17316 4632 17368 4684
rect 17684 4632 17736 4684
rect 18788 4632 18840 4684
rect 19156 4675 19208 4684
rect 19156 4641 19165 4675
rect 19165 4641 19199 4675
rect 19199 4641 19208 4675
rect 19156 4632 19208 4641
rect 19248 4632 19300 4684
rect 19984 4675 20036 4684
rect 19984 4641 19993 4675
rect 19993 4641 20027 4675
rect 20027 4641 20036 4675
rect 19984 4632 20036 4641
rect 20904 4675 20956 4684
rect 18052 4564 18104 4616
rect 18236 4607 18288 4616
rect 18236 4573 18245 4607
rect 18245 4573 18279 4607
rect 18279 4573 18288 4607
rect 18236 4564 18288 4573
rect 19616 4564 19668 4616
rect 12624 4496 12676 4548
rect 7380 4471 7432 4480
rect 7380 4437 7389 4471
rect 7389 4437 7423 4471
rect 7423 4437 7432 4471
rect 7380 4428 7432 4437
rect 8760 4428 8812 4480
rect 9312 4471 9364 4480
rect 9312 4437 9321 4471
rect 9321 4437 9355 4471
rect 9355 4437 9364 4471
rect 9312 4428 9364 4437
rect 12348 4471 12400 4480
rect 12348 4437 12357 4471
rect 12357 4437 12391 4471
rect 12391 4437 12400 4471
rect 12348 4428 12400 4437
rect 14188 4428 14240 4480
rect 15292 4428 15344 4480
rect 18880 4496 18932 4548
rect 19156 4428 19208 4480
rect 19800 4496 19852 4548
rect 19340 4428 19392 4480
rect 20076 4428 20128 4480
rect 20168 4428 20220 4480
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 21456 4675 21508 4684
rect 21456 4641 21465 4675
rect 21465 4641 21499 4675
rect 21499 4641 21508 4675
rect 21456 4632 21508 4641
rect 21824 4564 21876 4616
rect 20996 4471 21048 4480
rect 20996 4437 21005 4471
rect 21005 4437 21039 4471
rect 21039 4437 21048 4471
rect 20996 4428 21048 4437
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 2688 4267 2740 4276
rect 2688 4233 2697 4267
rect 2697 4233 2731 4267
rect 2731 4233 2740 4267
rect 2688 4224 2740 4233
rect 7196 4224 7248 4276
rect 7564 4224 7616 4276
rect 8852 4224 8904 4276
rect 2872 4156 2924 4208
rect 1308 4020 1360 4072
rect 2964 4088 3016 4140
rect 4712 4156 4764 4208
rect 6736 4156 6788 4208
rect 3976 4020 4028 4072
rect 5080 4088 5132 4140
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 6000 4088 6052 4140
rect 4436 4020 4488 4072
rect 4620 4063 4672 4072
rect 4620 4029 4629 4063
rect 4629 4029 4663 4063
rect 4663 4029 4672 4063
rect 4620 4020 4672 4029
rect 3332 3952 3384 4004
rect 3608 3952 3660 4004
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 1860 3884 1912 3936
rect 3976 3884 4028 3936
rect 4160 3927 4212 3936
rect 4160 3893 4169 3927
rect 4169 3893 4203 3927
rect 4203 3893 4212 3927
rect 4160 3884 4212 3893
rect 4344 3884 4396 3936
rect 4436 3927 4488 3936
rect 4436 3893 4445 3927
rect 4445 3893 4479 3927
rect 4479 3893 4488 3927
rect 5724 3952 5776 4004
rect 7380 4020 7432 4072
rect 7472 4020 7524 4072
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 9312 4224 9364 4276
rect 14372 4224 14424 4276
rect 15292 4224 15344 4276
rect 15752 4267 15804 4276
rect 15752 4233 15761 4267
rect 15761 4233 15795 4267
rect 15795 4233 15804 4267
rect 15752 4224 15804 4233
rect 17684 4267 17736 4276
rect 17684 4233 17693 4267
rect 17693 4233 17727 4267
rect 17727 4233 17736 4267
rect 17684 4224 17736 4233
rect 18052 4224 18104 4276
rect 19340 4224 19392 4276
rect 20904 4224 20956 4276
rect 21456 4224 21508 4276
rect 9496 4199 9548 4208
rect 9496 4165 9505 4199
rect 9505 4165 9539 4199
rect 9539 4165 9548 4199
rect 9496 4156 9548 4165
rect 9864 4156 9916 4208
rect 8392 4020 8444 4072
rect 4436 3884 4488 3893
rect 4988 3884 5040 3936
rect 5356 3884 5408 3936
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 6644 3884 6696 3936
rect 6736 3884 6788 3936
rect 8208 3952 8260 4004
rect 9680 4088 9732 4140
rect 10876 4088 10928 4140
rect 12164 4131 12216 4140
rect 12164 4097 12173 4131
rect 12173 4097 12207 4131
rect 12207 4097 12216 4131
rect 12164 4088 12216 4097
rect 12532 4156 12584 4208
rect 16948 4156 17000 4208
rect 20536 4156 20588 4208
rect 20812 4199 20864 4208
rect 20812 4165 20821 4199
rect 20821 4165 20855 4199
rect 20855 4165 20864 4199
rect 20812 4156 20864 4165
rect 12624 4088 12676 4140
rect 13452 4088 13504 4140
rect 15292 4088 15344 4140
rect 8944 4020 8996 4072
rect 9404 3952 9456 4004
rect 10232 3952 10284 4004
rect 10600 4020 10652 4072
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 10968 3952 11020 4004
rect 9772 3884 9824 3936
rect 10048 3884 10100 3936
rect 10416 3884 10468 3936
rect 13084 4020 13136 4072
rect 13268 4020 13320 4072
rect 12532 3952 12584 4004
rect 14464 4020 14516 4072
rect 14648 4063 14700 4072
rect 14648 4029 14657 4063
rect 14657 4029 14691 4063
rect 14691 4029 14700 4063
rect 14648 4020 14700 4029
rect 17592 4088 17644 4140
rect 19156 4088 19208 4140
rect 19800 4131 19852 4140
rect 13728 3952 13780 4004
rect 12164 3884 12216 3936
rect 12716 3927 12768 3936
rect 12716 3893 12725 3927
rect 12725 3893 12759 3927
rect 12759 3893 12768 3927
rect 12716 3884 12768 3893
rect 12808 3927 12860 3936
rect 12808 3893 12817 3927
rect 12817 3893 12851 3927
rect 12851 3893 12860 3927
rect 12808 3884 12860 3893
rect 13360 3884 13412 3936
rect 14556 3927 14608 3936
rect 14556 3893 14565 3927
rect 14565 3893 14599 3927
rect 14599 3893 14608 3927
rect 14556 3884 14608 3893
rect 14648 3884 14700 3936
rect 15936 4063 15988 4072
rect 15936 4029 15945 4063
rect 15945 4029 15979 4063
rect 15979 4029 15988 4063
rect 15936 4020 15988 4029
rect 16396 4020 16448 4072
rect 16580 4063 16632 4072
rect 16580 4029 16589 4063
rect 16589 4029 16623 4063
rect 16623 4029 16632 4063
rect 16580 4020 16632 4029
rect 16948 4063 17000 4072
rect 16948 4029 16957 4063
rect 16957 4029 16991 4063
rect 16991 4029 17000 4063
rect 16948 4020 17000 4029
rect 17960 4020 18012 4072
rect 19800 4097 19809 4131
rect 19809 4097 19843 4131
rect 19843 4097 19852 4131
rect 19800 4088 19852 4097
rect 19984 4131 20036 4140
rect 19984 4097 19993 4131
rect 19993 4097 20027 4131
rect 20027 4097 20036 4131
rect 19984 4088 20036 4097
rect 20076 4088 20128 4140
rect 19340 4020 19392 4072
rect 15384 3952 15436 4004
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 16304 3884 16356 3936
rect 16488 3927 16540 3936
rect 16488 3893 16497 3927
rect 16497 3893 16531 3927
rect 16531 3893 16540 3927
rect 16488 3884 16540 3893
rect 16764 3927 16816 3936
rect 16764 3893 16773 3927
rect 16773 3893 16807 3927
rect 16807 3893 16816 3927
rect 16764 3884 16816 3893
rect 17132 3927 17184 3936
rect 17132 3893 17141 3927
rect 17141 3893 17175 3927
rect 17175 3893 17184 3927
rect 17132 3884 17184 3893
rect 18696 3884 18748 3936
rect 18880 3952 18932 4004
rect 20444 4020 20496 4072
rect 20720 4063 20772 4072
rect 20720 4029 20729 4063
rect 20729 4029 20763 4063
rect 20763 4029 20772 4063
rect 20720 4020 20772 4029
rect 21272 4063 21324 4072
rect 21272 4029 21281 4063
rect 21281 4029 21315 4063
rect 21315 4029 21324 4063
rect 21272 4020 21324 4029
rect 21548 4063 21600 4072
rect 21548 4029 21557 4063
rect 21557 4029 21591 4063
rect 21591 4029 21600 4063
rect 21548 4020 21600 4029
rect 19524 3927 19576 3936
rect 19524 3893 19533 3927
rect 19533 3893 19567 3927
rect 19567 3893 19576 3927
rect 19524 3884 19576 3893
rect 19708 3884 19760 3936
rect 20904 3884 20956 3936
rect 22100 3884 22152 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 2044 3680 2096 3732
rect 2228 3680 2280 3732
rect 3424 3680 3476 3732
rect 4344 3680 4396 3732
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 2780 3612 2832 3664
rect 5448 3680 5500 3732
rect 8300 3680 8352 3732
rect 8760 3680 8812 3732
rect 9036 3680 9088 3732
rect 9772 3680 9824 3732
rect 10324 3680 10376 3732
rect 11980 3680 12032 3732
rect 12532 3680 12584 3732
rect 12716 3723 12768 3732
rect 12716 3689 12725 3723
rect 12725 3689 12759 3723
rect 12759 3689 12768 3723
rect 12716 3680 12768 3689
rect 4712 3612 4764 3664
rect 2872 3544 2924 3596
rect 4528 3544 4580 3596
rect 2596 3519 2648 3528
rect 2596 3485 2605 3519
rect 2605 3485 2639 3519
rect 2639 3485 2648 3519
rect 2596 3476 2648 3485
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 3608 3519 3660 3528
rect 2688 3476 2740 3485
rect 3608 3485 3617 3519
rect 3617 3485 3651 3519
rect 3651 3485 3660 3519
rect 3608 3476 3660 3485
rect 3884 3519 3936 3528
rect 3884 3485 3893 3519
rect 3893 3485 3927 3519
rect 3927 3485 3936 3519
rect 3884 3476 3936 3485
rect 3976 3476 4028 3528
rect 4896 3544 4948 3596
rect 5264 3612 5316 3664
rect 5724 3612 5776 3664
rect 6092 3612 6144 3664
rect 7472 3612 7524 3664
rect 9220 3655 9272 3664
rect 7104 3544 7156 3596
rect 8208 3544 8260 3596
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 6092 3476 6144 3528
rect 6920 3476 6972 3528
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8576 3587 8628 3596
rect 8576 3553 8585 3587
rect 8585 3553 8619 3587
rect 8619 3553 8628 3587
rect 8576 3544 8628 3553
rect 9220 3621 9229 3655
rect 9229 3621 9263 3655
rect 9263 3621 9272 3655
rect 9220 3612 9272 3621
rect 10048 3612 10100 3664
rect 10784 3612 10836 3664
rect 12440 3612 12492 3664
rect 14188 3680 14240 3732
rect 14740 3680 14792 3732
rect 12900 3612 12952 3664
rect 8116 3476 8168 3485
rect 8484 3476 8536 3528
rect 2504 3408 2556 3460
rect 1676 3340 1728 3392
rect 2228 3340 2280 3392
rect 3240 3340 3292 3392
rect 3424 3340 3476 3392
rect 6828 3408 6880 3460
rect 8208 3408 8260 3460
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 7748 3340 7800 3392
rect 9220 3340 9272 3392
rect 9680 3340 9732 3392
rect 10692 3340 10744 3392
rect 11704 3544 11756 3596
rect 13360 3544 13412 3596
rect 13544 3544 13596 3596
rect 14096 3612 14148 3664
rect 14556 3612 14608 3664
rect 15108 3544 15160 3596
rect 17132 3612 17184 3664
rect 18788 3680 18840 3732
rect 12624 3519 12676 3528
rect 12624 3485 12633 3519
rect 12633 3485 12667 3519
rect 12667 3485 12676 3519
rect 12624 3476 12676 3485
rect 12900 3476 12952 3528
rect 17224 3587 17276 3596
rect 17224 3553 17242 3587
rect 17242 3553 17276 3587
rect 17592 3587 17644 3596
rect 17224 3544 17276 3553
rect 17592 3553 17601 3587
rect 17601 3553 17635 3587
rect 17635 3553 17644 3587
rect 17592 3544 17644 3553
rect 12992 3408 13044 3460
rect 16212 3476 16264 3528
rect 18236 3544 18288 3596
rect 18512 3544 18564 3596
rect 18144 3476 18196 3528
rect 20536 3612 20588 3664
rect 21364 3655 21416 3664
rect 21364 3621 21373 3655
rect 21373 3621 21407 3655
rect 21407 3621 21416 3655
rect 21364 3612 21416 3621
rect 19984 3587 20036 3596
rect 19984 3553 19993 3587
rect 19993 3553 20027 3587
rect 20027 3553 20036 3587
rect 19984 3544 20036 3553
rect 20628 3544 20680 3596
rect 21640 3544 21692 3596
rect 19524 3476 19576 3528
rect 15292 3408 15344 3460
rect 16396 3408 16448 3460
rect 17592 3408 17644 3460
rect 19616 3451 19668 3460
rect 11060 3340 11112 3392
rect 13176 3383 13228 3392
rect 13176 3349 13185 3383
rect 13185 3349 13219 3383
rect 13219 3349 13228 3383
rect 13176 3340 13228 3349
rect 13544 3340 13596 3392
rect 15844 3340 15896 3392
rect 15936 3383 15988 3392
rect 15936 3349 15945 3383
rect 15945 3349 15979 3383
rect 15979 3349 15988 3383
rect 15936 3340 15988 3349
rect 16304 3340 16356 3392
rect 17316 3340 17368 3392
rect 17684 3340 17736 3392
rect 18788 3340 18840 3392
rect 19064 3383 19116 3392
rect 19064 3349 19073 3383
rect 19073 3349 19107 3383
rect 19107 3349 19116 3383
rect 19064 3340 19116 3349
rect 19340 3383 19392 3392
rect 19340 3349 19349 3383
rect 19349 3349 19383 3383
rect 19383 3349 19392 3383
rect 19340 3340 19392 3349
rect 19616 3417 19625 3451
rect 19625 3417 19659 3451
rect 19659 3417 19668 3451
rect 19616 3408 19668 3417
rect 19800 3476 19852 3528
rect 21088 3476 21140 3528
rect 20260 3408 20312 3460
rect 20996 3408 21048 3460
rect 21916 3408 21968 3460
rect 20628 3383 20680 3392
rect 20628 3349 20637 3383
rect 20637 3349 20671 3383
rect 20671 3349 20680 3383
rect 20628 3340 20680 3349
rect 22744 3340 22796 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 2596 3136 2648 3188
rect 3700 3136 3752 3188
rect 5080 3136 5132 3188
rect 5724 3136 5776 3188
rect 5816 3136 5868 3188
rect 6644 3136 6696 3188
rect 8300 3136 8352 3188
rect 8484 3179 8536 3188
rect 8484 3145 8493 3179
rect 8493 3145 8527 3179
rect 8527 3145 8536 3179
rect 8484 3136 8536 3145
rect 1308 2932 1360 2984
rect 2136 3000 2188 3052
rect 1860 2975 1912 2984
rect 1860 2941 1869 2975
rect 1869 2941 1903 2975
rect 1903 2941 1912 2975
rect 1860 2932 1912 2941
rect 2228 2975 2280 2984
rect 2228 2941 2237 2975
rect 2237 2941 2271 2975
rect 2271 2941 2280 2975
rect 2228 2932 2280 2941
rect 2688 2975 2740 2984
rect 2688 2941 2697 2975
rect 2697 2941 2731 2975
rect 2731 2941 2740 2975
rect 2688 2932 2740 2941
rect 3148 2932 3200 2984
rect 204 2864 256 2916
rect 1492 2864 1544 2916
rect 2412 2839 2464 2848
rect 2412 2805 2421 2839
rect 2421 2805 2455 2839
rect 2455 2805 2464 2839
rect 2412 2796 2464 2805
rect 2504 2839 2556 2848
rect 2504 2805 2513 2839
rect 2513 2805 2547 2839
rect 2547 2805 2556 2839
rect 3240 2864 3292 2916
rect 3516 3068 3568 3120
rect 5448 3068 5500 3120
rect 6092 3068 6144 3120
rect 6368 3068 6420 3120
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 3792 3000 3844 3052
rect 7104 3068 7156 3120
rect 8208 3068 8260 3120
rect 9404 3068 9456 3120
rect 4160 2975 4212 2984
rect 4160 2941 4194 2975
rect 4194 2941 4212 2975
rect 4160 2932 4212 2941
rect 4712 2932 4764 2984
rect 5172 2932 5224 2984
rect 7656 2932 7708 2984
rect 8760 3000 8812 3052
rect 8852 2975 8904 2984
rect 4896 2864 4948 2916
rect 6644 2907 6696 2916
rect 2504 2796 2556 2805
rect 3424 2839 3476 2848
rect 3424 2805 3433 2839
rect 3433 2805 3467 2839
rect 3467 2805 3476 2839
rect 3424 2796 3476 2805
rect 4160 2796 4212 2848
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 6644 2873 6653 2907
rect 6653 2873 6687 2907
rect 6687 2873 6696 2907
rect 6644 2864 6696 2873
rect 8116 2864 8168 2916
rect 8852 2941 8861 2975
rect 8861 2941 8895 2975
rect 8895 2941 8904 2975
rect 9772 3136 9824 3188
rect 11152 3136 11204 3188
rect 11704 3179 11756 3188
rect 11704 3145 11713 3179
rect 11713 3145 11747 3179
rect 11747 3145 11756 3179
rect 11704 3136 11756 3145
rect 10784 3068 10836 3120
rect 15200 3136 15252 3188
rect 13084 3068 13136 3120
rect 13176 3000 13228 3052
rect 8852 2932 8904 2941
rect 9680 2932 9732 2984
rect 10692 2932 10744 2984
rect 10968 2932 11020 2984
rect 10140 2864 10192 2916
rect 10232 2864 10284 2916
rect 8760 2796 8812 2848
rect 9772 2796 9824 2848
rect 10876 2796 10928 2848
rect 11152 2864 11204 2916
rect 12992 2932 13044 2984
rect 13360 2932 13412 2984
rect 13544 2975 13596 2984
rect 13544 2941 13553 2975
rect 13553 2941 13587 2975
rect 13587 2941 13596 2975
rect 13544 2932 13596 2941
rect 12716 2864 12768 2916
rect 12900 2864 12952 2916
rect 16580 3068 16632 3120
rect 17592 3136 17644 3188
rect 18880 3136 18932 3188
rect 19984 3136 20036 3188
rect 19248 3068 19300 3120
rect 19616 3068 19668 3120
rect 20812 3068 20864 3120
rect 18052 3000 18104 3052
rect 18236 3000 18288 3052
rect 19340 3000 19392 3052
rect 14372 2932 14424 2984
rect 14648 2932 14700 2984
rect 15108 2975 15160 2984
rect 15108 2941 15117 2975
rect 15117 2941 15151 2975
rect 15151 2941 15160 2975
rect 15108 2932 15160 2941
rect 15384 2975 15436 2984
rect 15384 2941 15393 2975
rect 15393 2941 15427 2975
rect 15427 2941 15436 2975
rect 15384 2932 15436 2941
rect 15844 2975 15896 2984
rect 15844 2941 15853 2975
rect 15853 2941 15887 2975
rect 15887 2941 15896 2975
rect 15844 2932 15896 2941
rect 15936 2932 15988 2984
rect 16488 2932 16540 2984
rect 18420 2932 18472 2984
rect 19524 2975 19576 2984
rect 19524 2941 19533 2975
rect 19533 2941 19567 2975
rect 19567 2941 19576 2975
rect 19524 2932 19576 2941
rect 20628 3000 20680 3052
rect 15660 2907 15712 2916
rect 11336 2796 11388 2848
rect 11704 2796 11756 2848
rect 12348 2796 12400 2848
rect 13176 2839 13228 2848
rect 13176 2805 13185 2839
rect 13185 2805 13219 2839
rect 13219 2805 13228 2839
rect 13176 2796 13228 2805
rect 13268 2796 13320 2848
rect 15660 2873 15669 2907
rect 15669 2873 15703 2907
rect 15703 2873 15712 2907
rect 15660 2864 15712 2873
rect 16028 2907 16080 2916
rect 16028 2873 16037 2907
rect 16037 2873 16071 2907
rect 16071 2873 16080 2907
rect 16028 2864 16080 2873
rect 16396 2864 16448 2916
rect 14004 2839 14056 2848
rect 14004 2805 14013 2839
rect 14013 2805 14047 2839
rect 14047 2805 14056 2839
rect 14004 2796 14056 2805
rect 14464 2839 14516 2848
rect 14464 2805 14473 2839
rect 14473 2805 14507 2839
rect 14507 2805 14516 2839
rect 14464 2796 14516 2805
rect 14740 2839 14792 2848
rect 14740 2805 14749 2839
rect 14749 2805 14783 2839
rect 14783 2805 14792 2839
rect 14740 2796 14792 2805
rect 15200 2796 15252 2848
rect 15476 2796 15528 2848
rect 16488 2796 16540 2848
rect 17684 2796 17736 2848
rect 17960 2796 18012 2848
rect 18144 2864 18196 2916
rect 19340 2864 19392 2916
rect 19800 2907 19852 2916
rect 19800 2873 19809 2907
rect 19809 2873 19843 2907
rect 19843 2873 19852 2907
rect 19800 2864 19852 2873
rect 19892 2864 19944 2916
rect 20260 2907 20312 2916
rect 20260 2873 20269 2907
rect 20269 2873 20303 2907
rect 20303 2873 20312 2907
rect 20260 2864 20312 2873
rect 20628 2907 20680 2916
rect 18236 2796 18288 2848
rect 18512 2796 18564 2848
rect 19708 2796 19760 2848
rect 20628 2873 20637 2907
rect 20637 2873 20671 2907
rect 20671 2873 20680 2907
rect 20628 2864 20680 2873
rect 22192 2932 22244 2984
rect 21456 2839 21508 2848
rect 21456 2805 21465 2839
rect 21465 2805 21499 2839
rect 21499 2805 21508 2839
rect 21456 2796 21508 2805
rect 22008 2839 22060 2848
rect 22008 2805 22017 2839
rect 22017 2805 22051 2839
rect 22051 2805 22060 2839
rect 22008 2796 22060 2805
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 1400 2592 1452 2644
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 3516 2592 3568 2644
rect 4804 2592 4856 2644
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 1492 2456 1544 2508
rect 1676 2499 1728 2508
rect 1676 2465 1685 2499
rect 1685 2465 1719 2499
rect 1719 2465 1728 2499
rect 1676 2456 1728 2465
rect 2596 2499 2648 2508
rect 572 2388 624 2440
rect 2596 2465 2605 2499
rect 2605 2465 2639 2499
rect 2639 2465 2648 2499
rect 2596 2456 2648 2465
rect 3884 2524 3936 2576
rect 4160 2524 4212 2576
rect 4712 2524 4764 2576
rect 6276 2592 6328 2644
rect 6736 2635 6788 2644
rect 6736 2601 6745 2635
rect 6745 2601 6779 2635
rect 6779 2601 6788 2635
rect 6736 2592 6788 2601
rect 7012 2635 7064 2644
rect 7012 2601 7021 2635
rect 7021 2601 7055 2635
rect 7055 2601 7064 2635
rect 7012 2592 7064 2601
rect 5816 2524 5868 2576
rect 7472 2592 7524 2644
rect 8668 2592 8720 2644
rect 9036 2592 9088 2644
rect 7564 2524 7616 2576
rect 9588 2567 9640 2576
rect 9588 2533 9597 2567
rect 9597 2533 9631 2567
rect 9631 2533 9640 2567
rect 9588 2524 9640 2533
rect 10048 2592 10100 2644
rect 10508 2635 10560 2644
rect 10508 2601 10517 2635
rect 10517 2601 10551 2635
rect 10551 2601 10560 2635
rect 10508 2592 10560 2601
rect 12164 2592 12216 2644
rect 12440 2592 12492 2644
rect 12808 2635 12860 2644
rect 12808 2601 12817 2635
rect 12817 2601 12851 2635
rect 12851 2601 12860 2635
rect 12808 2592 12860 2601
rect 13084 2592 13136 2644
rect 13176 2524 13228 2576
rect 13728 2524 13780 2576
rect 14004 2567 14056 2576
rect 14004 2533 14013 2567
rect 14013 2533 14047 2567
rect 14047 2533 14056 2567
rect 14004 2524 14056 2533
rect 4896 2499 4948 2508
rect 4896 2465 4905 2499
rect 4905 2465 4939 2499
rect 4939 2465 4948 2499
rect 4896 2456 4948 2465
rect 5448 2456 5500 2508
rect 6000 2499 6052 2508
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 6552 2456 6604 2508
rect 7196 2499 7248 2508
rect 7196 2465 7205 2499
rect 7205 2465 7239 2499
rect 7239 2465 7248 2499
rect 7196 2456 7248 2465
rect 1032 2320 1084 2372
rect 2504 2388 2556 2440
rect 3608 2388 3660 2440
rect 6092 2431 6144 2440
rect 3792 2320 3844 2372
rect 6092 2397 6101 2431
rect 6101 2397 6135 2431
rect 6135 2397 6144 2431
rect 6092 2388 6144 2397
rect 5264 2320 5316 2372
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 2044 2252 2096 2304
rect 2136 2295 2188 2304
rect 2136 2261 2145 2295
rect 2145 2261 2179 2295
rect 2179 2261 2188 2295
rect 2136 2252 2188 2261
rect 4804 2252 4856 2304
rect 8668 2456 8720 2508
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 7656 2320 7708 2372
rect 8576 2320 8628 2372
rect 9404 2320 9456 2372
rect 12716 2456 12768 2508
rect 12992 2456 13044 2508
rect 13268 2499 13320 2508
rect 13268 2465 13277 2499
rect 13277 2465 13311 2499
rect 13311 2465 13320 2499
rect 13268 2456 13320 2465
rect 11060 2431 11112 2440
rect 11060 2397 11069 2431
rect 11069 2397 11103 2431
rect 11103 2397 11112 2431
rect 11060 2388 11112 2397
rect 12348 2388 12400 2440
rect 13452 2456 13504 2508
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14188 2456 14240 2465
rect 14464 2524 14516 2576
rect 14832 2524 14884 2576
rect 17040 2592 17092 2644
rect 17960 2592 18012 2644
rect 15568 2524 15620 2576
rect 16580 2567 16632 2576
rect 16580 2533 16589 2567
rect 16589 2533 16623 2567
rect 16623 2533 16632 2567
rect 16580 2524 16632 2533
rect 16764 2524 16816 2576
rect 17408 2567 17460 2576
rect 17408 2533 17417 2567
rect 17417 2533 17451 2567
rect 17451 2533 17460 2567
rect 17408 2524 17460 2533
rect 17776 2524 17828 2576
rect 18604 2635 18656 2644
rect 18604 2601 18613 2635
rect 18613 2601 18647 2635
rect 18647 2601 18656 2635
rect 19064 2635 19116 2644
rect 18604 2592 18656 2601
rect 19064 2601 19073 2635
rect 19073 2601 19107 2635
rect 19107 2601 19116 2635
rect 19064 2592 19116 2601
rect 19340 2592 19392 2644
rect 20352 2592 20404 2644
rect 19432 2524 19484 2576
rect 20812 2567 20864 2576
rect 20812 2533 20821 2567
rect 20821 2533 20855 2567
rect 20855 2533 20864 2567
rect 20812 2524 20864 2533
rect 20996 2524 21048 2576
rect 15200 2456 15252 2508
rect 12072 2320 12124 2372
rect 8484 2252 8536 2304
rect 9036 2252 9088 2304
rect 11888 2252 11940 2304
rect 13544 2388 13596 2440
rect 15292 2388 15344 2440
rect 17316 2388 17368 2440
rect 18236 2456 18288 2508
rect 18052 2388 18104 2440
rect 19708 2456 19760 2508
rect 18880 2388 18932 2440
rect 19248 2388 19300 2440
rect 21088 2388 21140 2440
rect 12716 2320 12768 2372
rect 14832 2320 14884 2372
rect 16856 2320 16908 2372
rect 17684 2320 17736 2372
rect 14372 2252 14424 2304
rect 15384 2295 15436 2304
rect 15384 2261 15393 2295
rect 15393 2261 15427 2295
rect 15427 2261 15436 2295
rect 15384 2252 15436 2261
rect 15752 2295 15804 2304
rect 15752 2261 15761 2295
rect 15761 2261 15795 2295
rect 15795 2261 15804 2295
rect 15752 2252 15804 2261
rect 18604 2252 18656 2304
rect 19616 2252 19668 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 1584 2048 1636 2100
rect 6000 2048 6052 2100
rect 11796 2048 11848 2100
rect 6092 1980 6144 2032
rect 6460 1980 6512 2032
rect 10508 1980 10560 2032
rect 11428 1980 11480 2032
rect 13268 1980 13320 2032
rect 2044 1844 2096 1896
rect 3056 1776 3108 1828
rect 4896 1776 4948 1828
rect 6000 1776 6052 1828
rect 6552 1776 6604 1828
rect 8668 1912 8720 1964
rect 9864 1912 9916 1964
rect 8852 1844 8904 1896
rect 10140 1776 10192 1828
rect 2136 1708 2188 1760
rect 6460 1708 6512 1760
rect 7196 1708 7248 1760
rect 9680 1640 9732 1692
rect 9588 1572 9640 1624
rect 11244 1572 11296 1624
rect 14372 1436 14424 1488
rect 15752 1436 15804 1488
rect 14004 1368 14056 1420
rect 15384 1368 15436 1420
<< metal2 >>
rect 202 22200 258 23000
rect 570 22200 626 23000
rect 938 22200 994 23000
rect 1306 22200 1362 23000
rect 1398 22672 1454 22681
rect 1398 22607 1454 22616
rect 216 19854 244 22200
rect 584 20398 612 22200
rect 952 20466 980 22200
rect 940 20460 992 20466
rect 940 20402 992 20408
rect 572 20392 624 20398
rect 572 20334 624 20340
rect 204 19848 256 19854
rect 204 19790 256 19796
rect 1320 19242 1348 22200
rect 1412 20058 1440 22607
rect 1674 22200 1730 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2870 22200 2926 23000
rect 2962 22264 3018 22273
rect 1584 20324 1636 20330
rect 1584 20266 1636 20272
rect 1492 20256 1544 20262
rect 1490 20224 1492 20233
rect 1544 20224 1546 20233
rect 1490 20159 1546 20168
rect 1400 20052 1452 20058
rect 1400 19994 1452 20000
rect 1492 19712 1544 19718
rect 1490 19680 1492 19689
rect 1544 19680 1546 19689
rect 1490 19615 1546 19624
rect 1596 19514 1624 20266
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1400 19304 1452 19310
rect 1398 19272 1400 19281
rect 1452 19272 1454 19281
rect 1308 19236 1360 19242
rect 1398 19207 1454 19216
rect 1308 19178 1360 19184
rect 1320 18630 1348 19178
rect 1688 19174 1716 22200
rect 1858 20632 1914 20641
rect 1858 20567 1860 20576
rect 1912 20567 1914 20576
rect 1860 20538 1912 20544
rect 2056 20058 2084 22200
rect 2226 21040 2282 21049
rect 2226 20975 2282 20984
rect 2240 20602 2268 20975
rect 2228 20596 2280 20602
rect 2228 20538 2280 20544
rect 2412 20392 2464 20398
rect 2412 20334 2464 20340
rect 2136 20324 2188 20330
rect 2136 20266 2188 20272
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 1400 18896 1452 18902
rect 1398 18864 1400 18873
rect 1452 18864 1454 18873
rect 1780 18834 1808 19790
rect 1952 19304 2004 19310
rect 1950 19272 1952 19281
rect 2004 19272 2006 19281
rect 1860 19236 1912 19242
rect 1950 19207 2006 19216
rect 1860 19178 1912 19184
rect 1872 18970 1900 19178
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 1398 18799 1454 18808
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1308 18624 1360 18630
rect 1308 18566 1360 18572
rect 1858 18456 1914 18465
rect 1964 18426 1992 18770
rect 1858 18391 1860 18400
rect 1912 18391 1914 18400
rect 1952 18420 2004 18426
rect 1860 18362 1912 18368
rect 1952 18362 2004 18368
rect 2056 18329 2084 19858
rect 2148 18873 2176 20266
rect 2228 19984 2280 19990
rect 2228 19926 2280 19932
rect 2240 18970 2268 19926
rect 2332 19446 2360 20266
rect 2424 19922 2452 20334
rect 2516 20262 2544 22200
rect 2884 21962 2912 22200
rect 2962 22199 3018 22208
rect 3238 22200 3294 23000
rect 3606 22200 3662 23000
rect 3974 22200 4030 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5170 22200 5226 23000
rect 5538 22200 5594 23000
rect 5906 22200 5962 23000
rect 6274 22200 6330 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7470 22200 7526 23000
rect 7838 22200 7894 23000
rect 8206 22200 8262 23000
rect 8574 22200 8630 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9770 22200 9826 23000
rect 10138 22200 10194 23000
rect 10506 22200 10562 23000
rect 10874 22200 10930 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12070 22200 12126 23000
rect 12438 22200 12494 23000
rect 12806 22200 12862 23000
rect 13174 22200 13230 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14370 22200 14426 23000
rect 14738 22200 14794 23000
rect 15106 22200 15162 23000
rect 15474 22200 15530 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16670 22200 16726 23000
rect 17038 22200 17094 23000
rect 17406 22200 17462 23000
rect 17498 22264 17554 22273
rect 2872 21956 2924 21962
rect 2872 21898 2924 21904
rect 2870 21856 2926 21865
rect 2870 21791 2926 21800
rect 2778 21448 2834 21457
rect 2778 21383 2834 21392
rect 2792 20602 2820 21383
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2884 20534 2912 21791
rect 2872 20528 2924 20534
rect 2872 20470 2924 20476
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2596 20324 2648 20330
rect 2596 20266 2648 20272
rect 2504 20256 2556 20262
rect 2504 20198 2556 20204
rect 2412 19916 2464 19922
rect 2412 19858 2464 19864
rect 2424 19514 2452 19858
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 2320 19440 2372 19446
rect 2320 19382 2372 19388
rect 2504 19304 2556 19310
rect 2504 19246 2556 19252
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2134 18864 2190 18873
rect 2134 18799 2190 18808
rect 2042 18320 2098 18329
rect 2042 18255 2098 18264
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 1544 18048 1546 18057
rect 1490 17983 1546 17992
rect 2424 17921 2452 19110
rect 2516 18970 2544 19246
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 2516 18601 2544 18770
rect 2608 18737 2636 20266
rect 2700 19922 2728 20402
rect 2778 19952 2834 19961
rect 2688 19916 2740 19922
rect 2778 19887 2834 19896
rect 2688 19858 2740 19864
rect 2700 19378 2728 19858
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2792 19310 2820 19887
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2688 19236 2740 19242
rect 2688 19178 2740 19184
rect 2594 18728 2650 18737
rect 2594 18663 2650 18672
rect 2700 18630 2728 19178
rect 2688 18624 2740 18630
rect 2502 18592 2558 18601
rect 2688 18566 2740 18572
rect 2502 18527 2558 18536
rect 2884 18426 2912 19654
rect 2976 19174 3004 22199
rect 3148 21956 3200 21962
rect 3148 21898 3200 21904
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3068 19922 3096 19994
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 3068 18834 3096 19858
rect 3160 19242 3188 21898
rect 3252 20398 3280 22200
rect 3240 20392 3292 20398
rect 3620 20380 3648 22200
rect 3700 20392 3752 20398
rect 3620 20352 3700 20380
rect 3240 20334 3292 20340
rect 3700 20334 3752 20340
rect 3988 20262 4016 22200
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3240 20052 3292 20058
rect 3240 19994 3292 20000
rect 3252 19718 3280 19994
rect 3344 19922 3372 20198
rect 3884 19984 3936 19990
rect 3884 19926 3936 19932
rect 3976 19984 4028 19990
rect 3976 19926 4028 19932
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 3700 19916 3752 19922
rect 3700 19858 3752 19864
rect 3240 19712 3292 19718
rect 3240 19654 3292 19660
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 3160 18970 3188 19178
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 3252 18290 3280 19654
rect 3344 18902 3372 19858
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3332 18896 3384 18902
rect 3332 18838 3384 18844
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3436 18086 3464 19654
rect 3712 19514 3740 19858
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 3804 19417 3832 19654
rect 3790 19408 3846 19417
rect 3790 19343 3846 19352
rect 3792 19168 3844 19174
rect 3792 19110 3844 19116
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 2410 17912 2466 17921
rect 2410 17847 2466 17856
rect 1952 17740 2004 17746
rect 1952 17682 2004 17688
rect 1766 17640 1822 17649
rect 1766 17575 1768 17584
rect 1820 17575 1822 17584
rect 1768 17546 1820 17552
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17241 1532 17478
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1768 17060 1820 17066
rect 1768 17002 1820 17008
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1504 16833 1532 16934
rect 1490 16824 1546 16833
rect 1780 16794 1808 17002
rect 1964 16794 1992 17682
rect 2412 17672 2464 17678
rect 2976 17649 3004 18022
rect 3160 17882 3188 18022
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3240 17808 3292 17814
rect 3240 17750 3292 17756
rect 2412 17614 2464 17620
rect 2962 17640 3018 17649
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 2320 17536 2372 17542
rect 2320 17478 2372 17484
rect 2240 17134 2268 17478
rect 2332 17202 2360 17478
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 1490 16759 1546 16768
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1504 16289 1532 16390
rect 1490 16280 1546 16289
rect 1490 16215 1546 16224
rect 1780 16114 1808 16730
rect 2320 16652 2372 16658
rect 2424 16640 2452 17614
rect 2596 17604 2648 17610
rect 2962 17575 3018 17584
rect 2596 17546 2648 17552
rect 2608 17270 2636 17546
rect 3252 17490 3280 17750
rect 3252 17462 3464 17490
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 2372 16612 2452 16640
rect 2320 16594 2372 16600
rect 2332 16114 2360 16594
rect 3160 16590 3188 17002
rect 3240 16720 3292 16726
rect 3240 16662 3292 16668
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2424 16250 2452 16390
rect 3252 16250 3280 16662
rect 3344 16250 3372 17274
rect 3436 16810 3464 17462
rect 3528 16946 3556 18702
rect 3608 18148 3660 18154
rect 3608 18090 3660 18096
rect 3620 17678 3648 18090
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3712 17542 3740 18022
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3804 17202 3832 19110
rect 3896 18902 3924 19926
rect 3988 19514 4016 19926
rect 4068 19916 4120 19922
rect 4356 19904 4384 22200
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4436 20460 4488 20466
rect 4436 20402 4488 20408
rect 4120 19876 4384 19904
rect 4068 19858 4120 19864
rect 4448 19802 4476 20402
rect 4816 20398 4844 22200
rect 5080 20528 5132 20534
rect 5080 20470 5132 20476
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 4712 20256 4764 20262
rect 4710 20224 4712 20233
rect 4764 20224 4766 20233
rect 4710 20159 4766 20168
rect 4068 19780 4120 19786
rect 4068 19722 4120 19728
rect 4356 19774 4476 19802
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3974 19272 4030 19281
rect 3974 19207 4030 19216
rect 3884 18896 3936 18902
rect 3884 18838 3936 18844
rect 3988 18834 4016 19207
rect 4080 18970 4108 19722
rect 4160 19168 4212 19174
rect 4356 19145 4384 19774
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4816 19496 4844 20334
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4632 19468 4844 19496
rect 4632 19242 4660 19468
rect 4908 19394 4936 20198
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 4724 19366 4936 19394
rect 4724 19334 4752 19366
rect 4724 19306 4844 19334
rect 5000 19310 5028 19654
rect 4620 19236 4672 19242
rect 4620 19178 4672 19184
rect 4160 19110 4212 19116
rect 4342 19136 4398 19145
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 3884 18624 3936 18630
rect 3882 18592 3884 18601
rect 3936 18592 3938 18601
rect 3882 18527 3938 18536
rect 3988 18193 4016 18770
rect 3974 18184 4030 18193
rect 4080 18154 4108 18906
rect 4172 18358 4200 19110
rect 4342 19071 4398 19080
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 3974 18119 4030 18128
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 3988 17814 4016 18022
rect 4264 17882 4292 18702
rect 4436 18692 4488 18698
rect 4356 18652 4436 18680
rect 4356 18290 4384 18652
rect 4436 18634 4488 18640
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4526 17912 4582 17921
rect 4252 17876 4304 17882
rect 4526 17847 4528 17856
rect 4252 17818 4304 17824
rect 4580 17847 4582 17856
rect 4528 17818 4580 17824
rect 3976 17808 4028 17814
rect 3976 17750 4028 17756
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3528 16918 3648 16946
rect 3436 16782 3556 16810
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 1858 15872 1914 15881
rect 1858 15807 1914 15816
rect 1872 15706 1900 15807
rect 2332 15706 2360 16050
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 1398 15464 1454 15473
rect 1398 15399 1400 15408
rect 1452 15399 1454 15408
rect 1400 15370 1452 15376
rect 1596 15094 1624 15506
rect 1964 15162 1992 15506
rect 2044 15360 2096 15366
rect 2044 15302 2096 15308
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 1584 15088 1636 15094
rect 1398 15056 1454 15065
rect 1584 15030 1636 15036
rect 1398 14991 1400 15000
rect 1452 14991 1454 15000
rect 1400 14962 1452 14968
rect 2056 14958 2084 15302
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 1858 14648 1914 14657
rect 1858 14583 1860 14592
rect 1912 14583 1914 14592
rect 1860 14554 1912 14560
rect 2056 14550 2084 14894
rect 2044 14544 2096 14550
rect 2044 14486 2096 14492
rect 1492 14272 1544 14278
rect 1490 14240 1492 14249
rect 1544 14240 1546 14249
rect 1490 14175 1546 14184
rect 2240 14074 2268 14894
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2424 14006 2452 14350
rect 2516 14278 2544 14758
rect 2792 14618 2820 15846
rect 2884 15162 2912 15914
rect 3436 15706 3464 16594
rect 3528 16522 3556 16782
rect 3516 16516 3568 16522
rect 3516 16458 3568 16464
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3240 15632 3292 15638
rect 3240 15574 3292 15580
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 3252 15026 3280 15574
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2872 14544 2924 14550
rect 3148 14544 3200 14550
rect 2924 14492 3004 14498
rect 2872 14486 3004 14492
rect 3148 14486 3200 14492
rect 2884 14470 3004 14486
rect 2872 14340 2924 14346
rect 2872 14282 2924 14288
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 1400 13864 1452 13870
rect 1768 13864 1820 13870
rect 1400 13806 1452 13812
rect 1766 13832 1768 13841
rect 2320 13864 2372 13870
rect 1820 13832 1822 13841
rect 1412 13433 1440 13806
rect 2320 13806 2372 13812
rect 1766 13767 1822 13776
rect 2136 13796 2188 13802
rect 2136 13738 2188 13744
rect 2148 13530 2176 13738
rect 2332 13530 2360 13806
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 1398 13424 1454 13433
rect 2424 13394 2452 13670
rect 1398 13359 1454 13368
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 1768 13252 1820 13258
rect 1768 13194 1820 13200
rect 1400 13184 1452 13190
rect 1400 13126 1452 13132
rect 1412 12481 1440 13126
rect 1780 12782 1808 13194
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12889 1900 13126
rect 1964 12986 1992 13330
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 1858 12880 1914 12889
rect 1858 12815 1914 12824
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1952 12708 2004 12714
rect 1952 12650 2004 12656
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1398 12472 1454 12481
rect 1398 12407 1454 12416
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1412 10849 1440 12242
rect 1504 12073 1532 12582
rect 1964 12238 1992 12650
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1490 12064 1546 12073
rect 1490 11999 1546 12008
rect 1964 11898 1992 12174
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 1582 11792 1638 11801
rect 1582 11727 1638 11736
rect 1596 11354 1624 11727
rect 2044 11620 2096 11626
rect 2044 11562 2096 11568
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1398 10840 1454 10849
rect 1398 10775 1454 10784
rect 1504 10441 1532 11154
rect 1688 10674 1716 11290
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1768 10464 1820 10470
rect 1490 10432 1546 10441
rect 1768 10406 1820 10412
rect 1490 10367 1546 10376
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1688 9586 1716 9998
rect 1780 9722 1808 10406
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1950 9344 2006 9353
rect 1504 8362 1532 9318
rect 1950 9279 2006 9288
rect 1766 8664 1822 8673
rect 1766 8599 1768 8608
rect 1820 8599 1822 8608
rect 1768 8570 1820 8576
rect 1780 8430 1808 8570
rect 1964 8566 1992 9279
rect 1860 8560 1912 8566
rect 1858 8528 1860 8537
rect 1952 8560 2004 8566
rect 1912 8528 1914 8537
rect 1952 8502 2004 8508
rect 1858 8463 1914 8472
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 7857 1532 8298
rect 1674 8120 1730 8129
rect 1674 8055 1730 8064
rect 1490 7848 1546 7857
rect 1490 7783 1546 7792
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1504 7041 1532 7278
rect 1490 7032 1546 7041
rect 1490 6967 1546 6976
rect 1688 6934 1716 8055
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1964 7546 1992 7890
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1676 6928 1728 6934
rect 1490 6896 1546 6905
rect 2056 6914 2084 11562
rect 2240 10810 2268 12242
rect 2516 10826 2544 14214
rect 2884 13394 2912 14282
rect 2976 14074 3004 14470
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3160 13802 3188 14486
rect 3252 14414 3280 14962
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3528 14618 3556 14758
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 2608 12442 2636 13330
rect 2976 13274 3004 13330
rect 2884 13246 3004 13274
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 11694 2636 12038
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2608 11354 2636 11630
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2424 10798 2544 10826
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 8906 2176 9998
rect 2240 9994 2268 10406
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2332 9178 2360 9318
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2136 8900 2188 8906
rect 2136 8842 2188 8848
rect 2136 8288 2188 8294
rect 2136 8230 2188 8236
rect 2148 8022 2176 8230
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 2134 7168 2190 7177
rect 2134 7103 2190 7112
rect 1676 6870 1728 6876
rect 1964 6886 2084 6914
rect 1490 6831 1492 6840
rect 1544 6831 1546 6840
rect 1492 6802 1544 6808
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 1122 6216 1178 6225
rect 1122 6151 1178 6160
rect 1216 6180 1268 6186
rect 938 5808 994 5817
rect 938 5743 994 5752
rect 204 2916 256 2922
rect 204 2858 256 2864
rect 216 800 244 2858
rect 572 2440 624 2446
rect 572 2382 624 2388
rect 584 800 612 2382
rect 952 1873 980 5743
rect 1032 2372 1084 2378
rect 1032 2314 1084 2320
rect 938 1864 994 1873
rect 938 1799 994 1808
rect 1044 800 1072 2314
rect 1136 1057 1164 6151
rect 1216 6122 1268 6128
rect 1228 5681 1256 6122
rect 1308 5772 1360 5778
rect 1308 5714 1360 5720
rect 1214 5672 1270 5681
rect 1214 5607 1270 5616
rect 1320 5273 1348 5714
rect 1306 5264 1362 5273
rect 1306 5199 1362 5208
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1320 4457 1348 5102
rect 1306 4448 1362 4457
rect 1306 4383 1362 4392
rect 1308 4072 1360 4078
rect 1306 4040 1308 4049
rect 1360 4040 1362 4049
rect 1306 3975 1362 3984
rect 1412 3641 1440 6598
rect 1504 6089 1532 6802
rect 1964 6458 1992 6886
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1490 6080 1546 6089
rect 1490 6015 1546 6024
rect 1780 5370 1808 6190
rect 1952 5840 2004 5846
rect 1952 5782 2004 5788
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1964 5234 1992 5782
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1766 4992 1822 5001
rect 1766 4927 1822 4936
rect 1582 4040 1638 4049
rect 1582 3975 1638 3984
rect 1596 3942 1624 3975
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1398 3632 1454 3641
rect 1398 3567 1400 3576
rect 1452 3567 1454 3576
rect 1400 3538 1452 3544
rect 1412 3507 1440 3538
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 1122 1048 1178 1057
rect 1122 983 1178 992
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1320 241 1348 2926
rect 1492 2916 1544 2922
rect 1492 2858 1544 2864
rect 1400 2644 1452 2650
rect 1400 2586 1452 2592
rect 1412 800 1440 2586
rect 1504 2514 1532 2858
rect 1688 2514 1716 3334
rect 1780 3097 1808 4927
rect 1964 4826 1992 5170
rect 2042 5128 2098 5137
rect 2042 5063 2098 5072
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1766 3088 1822 3097
rect 1766 3023 1822 3032
rect 1872 2990 1900 3878
rect 2056 3738 2084 5063
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2056 3097 2084 3130
rect 2042 3088 2098 3097
rect 2148 3058 2176 7103
rect 2332 7041 2360 8978
rect 2424 7313 2452 10798
rect 2596 10532 2648 10538
rect 2596 10474 2648 10480
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2410 7304 2466 7313
rect 2410 7239 2466 7248
rect 2318 7032 2374 7041
rect 2318 6967 2320 6976
rect 2372 6967 2374 6976
rect 2320 6938 2372 6944
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2240 6322 2268 6598
rect 2424 6390 2452 7239
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2516 6118 2544 9998
rect 2608 9994 2636 10474
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2608 9586 2636 9930
rect 2792 9674 2820 12718
rect 2884 12714 2912 13246
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2884 11762 2912 12650
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2976 11898 3004 12582
rect 3068 11898 3096 13398
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2884 10470 2912 11154
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2884 10198 2912 10406
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2688 9648 2740 9654
rect 2792 9646 2912 9674
rect 2688 9590 2740 9596
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2608 8974 2636 9522
rect 2700 9364 2728 9590
rect 2884 9518 2912 9646
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2700 9336 2820 9364
rect 2792 9178 2820 9336
rect 2884 9217 2912 9454
rect 2870 9208 2926 9217
rect 2780 9172 2832 9178
rect 2870 9143 2926 9152
rect 2780 9114 2832 9120
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2700 8838 2728 8978
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2700 6322 2728 8774
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2792 7562 2820 8366
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2884 7818 2912 8298
rect 2976 8022 3004 11494
rect 3160 10266 3188 13738
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3252 13326 3280 13670
rect 3330 13560 3386 13569
rect 3330 13495 3332 13504
rect 3384 13495 3386 13504
rect 3332 13466 3384 13472
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3252 12714 3280 13262
rect 3620 12753 3648 16918
rect 3882 16552 3938 16561
rect 3700 16516 3752 16522
rect 3882 16487 3938 16496
rect 3700 16458 3752 16464
rect 3712 15502 3740 16458
rect 3792 15972 3844 15978
rect 3792 15914 3844 15920
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3804 15434 3832 15914
rect 3792 15428 3844 15434
rect 3792 15370 3844 15376
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3606 12744 3662 12753
rect 3240 12708 3292 12714
rect 3606 12679 3662 12688
rect 3240 12650 3292 12656
rect 3712 12356 3740 14486
rect 3804 12434 3832 14758
rect 3896 14006 3924 16487
rect 3976 15088 4028 15094
rect 3976 15030 4028 15036
rect 3988 14414 4016 15030
rect 4080 14822 4108 17614
rect 4172 17270 4200 17682
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 4356 16726 4384 17274
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 4344 16720 4396 16726
rect 4344 16662 4396 16668
rect 4448 16436 4476 17002
rect 4356 16408 4476 16436
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4172 14958 4200 15438
rect 4264 15162 4292 15846
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4172 14618 4200 14894
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 3976 14408 4028 14414
rect 3974 14376 3976 14385
rect 4028 14376 4030 14385
rect 3974 14311 4030 14320
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3896 12617 3924 13942
rect 4172 13705 4200 14554
rect 4356 14550 4384 16408
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4436 15972 4488 15978
rect 4436 15914 4488 15920
rect 4448 15706 4476 15914
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4816 15620 4844 19306
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 4908 17882 4936 19246
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 5000 17678 5028 18226
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 5000 17202 5028 17614
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 4816 15592 4936 15620
rect 4712 15564 4764 15570
rect 4764 15524 4844 15552
rect 4712 15506 4764 15512
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4344 14544 4396 14550
rect 4344 14486 4396 14492
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 3974 13696 4030 13705
rect 3974 13631 4030 13640
rect 4158 13696 4214 13705
rect 4158 13631 4214 13640
rect 3988 13394 4016 13631
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 3988 12782 4016 13330
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3976 12640 4028 12646
rect 3882 12608 3938 12617
rect 3976 12582 4028 12588
rect 3882 12543 3938 12552
rect 3988 12442 4016 12582
rect 3976 12436 4028 12442
rect 3804 12406 3924 12434
rect 3712 12328 3832 12356
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3252 11354 3280 12174
rect 3620 11898 3648 12242
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3330 11248 3386 11257
rect 3330 11183 3332 11192
rect 3384 11183 3386 11192
rect 3332 11154 3384 11160
rect 3344 10266 3372 11154
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 8480 3096 9318
rect 3160 9178 3188 10066
rect 3436 9926 3464 10066
rect 3424 9920 3476 9926
rect 3422 9888 3424 9897
rect 3476 9888 3478 9897
rect 3422 9823 3478 9832
rect 3620 9674 3648 11494
rect 3712 11082 3740 11698
rect 3700 11076 3752 11082
rect 3700 11018 3752 11024
rect 3712 10470 3740 11018
rect 3804 10538 3832 12328
rect 3896 11558 3924 12406
rect 3976 12378 4028 12384
rect 4080 12374 4108 12786
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4066 11656 4122 11665
rect 4172 11642 4200 12242
rect 4264 11898 4292 14418
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4356 13530 4384 14350
rect 4448 14346 4476 14758
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4710 13832 4766 13841
rect 4710 13767 4712 13776
rect 4764 13767 4766 13776
rect 4712 13738 4764 13744
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4436 13388 4488 13394
rect 4356 13348 4436 13376
rect 4356 12986 4384 13348
rect 4436 13330 4488 13336
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4250 11656 4306 11665
rect 4172 11614 4250 11642
rect 4066 11591 4122 11600
rect 4356 11626 4384 12582
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4250 11591 4306 11600
rect 4344 11620 4396 11626
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3896 10810 3924 11086
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3804 9722 3832 10134
rect 3528 9646 3648 9674
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3240 9512 3292 9518
rect 3238 9480 3240 9489
rect 3292 9480 3294 9489
rect 3528 9450 3556 9646
rect 3238 9415 3294 9424
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3146 9072 3202 9081
rect 3620 9042 3648 9318
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 3146 9007 3148 9016
rect 3200 9007 3202 9016
rect 3608 9036 3660 9042
rect 3148 8978 3200 8984
rect 3608 8978 3660 8984
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3330 8936 3386 8945
rect 3068 8452 3188 8480
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3068 8090 3096 8298
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2962 7848 3018 7857
rect 2872 7812 2924 7818
rect 2962 7783 3018 7792
rect 2872 7754 2924 7760
rect 2792 7546 2912 7562
rect 2792 7540 2924 7546
rect 2792 7534 2872 7540
rect 2872 7482 2924 7488
rect 2976 7290 3004 7783
rect 2884 7274 3004 7290
rect 2872 7268 3004 7274
rect 2924 7262 3004 7268
rect 2872 7210 2924 7216
rect 3160 7002 3188 8452
rect 3252 7954 3280 8910
rect 3712 8922 3740 9046
rect 3896 9042 3924 10746
rect 3988 9654 4016 11290
rect 4080 11286 4108 11591
rect 4344 11562 4396 11568
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 4172 10742 4200 11494
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4264 10810 4292 11154
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4250 10704 4306 10713
rect 4250 10639 4306 10648
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4080 10266 4108 10542
rect 4264 10470 4292 10639
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4080 9674 4108 10202
rect 4264 9994 4292 10406
rect 4356 10266 4384 11086
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4540 10062 4568 10474
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 3976 9648 4028 9654
rect 4080 9646 4292 9674
rect 3976 9590 4028 9596
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3330 8871 3332 8880
rect 3384 8871 3386 8880
rect 3620 8894 3740 8922
rect 3332 8842 3384 8848
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3252 7449 3280 7890
rect 3344 7750 3372 8298
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3514 8256 3570 8265
rect 3436 7750 3464 8230
rect 3514 8191 3570 8200
rect 3528 7954 3556 8191
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3238 7440 3294 7449
rect 3238 7375 3294 7384
rect 3344 7342 3372 7686
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3252 6882 3280 7142
rect 3344 6934 3372 7142
rect 3068 6854 3280 6882
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2884 6202 2912 6326
rect 2700 6174 2912 6202
rect 2976 6202 3004 6734
rect 3068 6662 3096 6854
rect 3240 6792 3292 6798
rect 3436 6746 3464 7482
rect 3528 6934 3556 7890
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3620 6769 3648 8894
rect 3792 8424 3844 8430
rect 3896 8412 3924 8978
rect 3844 8384 3924 8412
rect 3792 8366 3844 8372
rect 3988 8242 4016 9590
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3804 8214 4016 8242
rect 3804 7546 3832 8214
rect 4080 8106 4108 9386
rect 4172 9042 4200 9522
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4172 8634 4200 8978
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4264 8294 4292 9646
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4816 8634 4844 15524
rect 4908 14090 4936 15592
rect 5000 15502 5028 17138
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 5000 14958 5028 15438
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 4988 14272 5040 14278
rect 4986 14240 4988 14249
rect 5040 14240 5042 14249
rect 4986 14175 5042 14184
rect 4908 14062 5028 14090
rect 4896 14000 4948 14006
rect 4896 13942 4948 13948
rect 4908 13462 4936 13942
rect 5000 13462 5028 14062
rect 4896 13456 4948 13462
rect 4896 13398 4948 13404
rect 4988 13456 5040 13462
rect 4988 13398 5040 13404
rect 5092 12782 5120 20470
rect 5184 20398 5212 22200
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5172 20392 5224 20398
rect 5172 20334 5224 20340
rect 5184 19174 5212 20334
rect 5276 19922 5304 20470
rect 5448 20324 5500 20330
rect 5448 20266 5500 20272
rect 5460 20058 5488 20266
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5552 19990 5580 22200
rect 5632 20392 5684 20398
rect 5684 20352 5856 20380
rect 5632 20334 5684 20340
rect 5630 20224 5686 20233
rect 5630 20159 5686 20168
rect 5540 19984 5592 19990
rect 5540 19926 5592 19932
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5276 18970 5304 19858
rect 5644 19378 5672 20159
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5736 19310 5764 19790
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5460 18834 5488 19246
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5446 18592 5502 18601
rect 5446 18527 5502 18536
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5184 18086 5212 18362
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17066 5212 18022
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 5276 16454 5304 17818
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 15638 5212 15846
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 5184 15366 5212 15574
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5264 14816 5316 14822
rect 5184 14776 5264 14804
rect 5184 14278 5212 14776
rect 5264 14758 5316 14764
rect 5172 14272 5224 14278
rect 5170 14240 5172 14249
rect 5224 14240 5226 14249
rect 5170 14175 5226 14184
rect 5368 13954 5396 18158
rect 5460 17921 5488 18527
rect 5446 17912 5502 17921
rect 5446 17847 5502 17856
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5460 17338 5488 17614
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5552 16114 5580 17750
rect 5644 17134 5672 18838
rect 5736 18630 5764 19246
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5736 17270 5764 18566
rect 5828 17320 5856 20352
rect 5920 19310 5948 22200
rect 6288 20398 6316 22200
rect 6000 20392 6052 20398
rect 6000 20334 6052 20340
rect 6276 20392 6328 20398
rect 6368 20392 6420 20398
rect 6276 20334 6328 20340
rect 6366 20360 6368 20369
rect 6420 20360 6422 20369
rect 6012 19990 6040 20334
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6000 19984 6052 19990
rect 6000 19926 6052 19932
rect 6012 19446 6040 19926
rect 6000 19440 6052 19446
rect 6000 19382 6052 19388
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 17814 6040 19110
rect 6104 18952 6132 20198
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6196 19514 6224 19654
rect 6288 19514 6316 20334
rect 6366 20295 6422 20304
rect 6656 19990 6684 22200
rect 7116 20806 7144 22200
rect 7104 20800 7156 20806
rect 7104 20742 7156 20748
rect 7116 20398 7144 20742
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 6736 20324 6788 20330
rect 6736 20266 6788 20272
rect 7288 20324 7340 20330
rect 7288 20266 7340 20272
rect 6644 19984 6696 19990
rect 6644 19926 6696 19932
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 6276 19508 6328 19514
rect 6564 19496 6592 19858
rect 6564 19468 6684 19496
rect 6276 19450 6328 19456
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6460 18964 6512 18970
rect 6104 18924 6408 18952
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5828 17292 5948 17320
rect 5724 17264 5776 17270
rect 5724 17206 5776 17212
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5184 13926 5396 13954
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 4988 12708 5040 12714
rect 4988 12650 5040 12656
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 12374 4936 12582
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4908 11694 4936 12038
rect 5000 11762 5028 12650
rect 5080 12368 5132 12374
rect 5080 12310 5132 12316
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 4908 9674 4936 11222
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5000 10198 5028 11154
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 4908 9646 5028 9674
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4908 8906 4936 9386
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4894 8392 4950 8401
rect 4894 8327 4950 8336
rect 4908 8294 4936 8327
rect 5000 8294 5028 9646
rect 5092 9586 5120 12310
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4264 8266 4384 8294
rect 4080 8078 4200 8106
rect 4068 8016 4120 8022
rect 4172 7993 4200 8078
rect 4068 7958 4120 7964
rect 4158 7984 4214 7993
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3292 6740 3464 6746
rect 3240 6734 3464 6740
rect 3148 6724 3200 6730
rect 3252 6718 3464 6734
rect 3606 6760 3662 6769
rect 3606 6695 3662 6704
rect 3148 6666 3200 6672
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2976 6174 3096 6202
rect 2700 6118 2728 6174
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2688 6112 2740 6118
rect 2964 6112 3016 6118
rect 2688 6054 2740 6060
rect 2870 6080 2926 6089
rect 2964 6054 3016 6060
rect 2870 6015 2926 6024
rect 2884 5914 2912 6015
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2700 5234 2728 5510
rect 2688 5228 2740 5234
rect 2608 5188 2688 5216
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2320 5024 2372 5030
rect 2504 5024 2556 5030
rect 2320 4966 2372 4972
rect 2424 4984 2504 5012
rect 2240 3738 2268 4966
rect 2332 4826 2360 4966
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2042 3023 2098 3032
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2240 2990 2268 3334
rect 2424 3074 2452 4984
rect 2504 4966 2556 4972
rect 2608 4486 2636 5188
rect 2688 5170 2740 5176
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2778 4856 2834 4865
rect 2778 4791 2834 4800
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2700 4282 2728 4626
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2700 3534 2728 4218
rect 2792 3670 2820 4791
rect 2884 4214 2912 5034
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2976 4146 3004 6054
rect 3068 4758 3096 6174
rect 3160 5914 3188 6666
rect 3238 6488 3294 6497
rect 3238 6423 3294 6432
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3252 5778 3280 6423
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3238 5672 3294 5681
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 3068 4026 3096 4490
rect 2976 3998 3096 4026
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2596 3528 2648 3534
rect 2502 3496 2558 3505
rect 2596 3470 2648 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2502 3431 2504 3440
rect 2556 3431 2558 3440
rect 2504 3402 2556 3408
rect 2608 3194 2636 3470
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2424 3046 2636 3074
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 1492 2508 1544 2514
rect 1492 2450 1544 2456
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1596 2106 1624 2246
rect 1584 2100 1636 2106
rect 1584 2042 1636 2048
rect 1872 800 1900 2926
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2056 1902 2084 2246
rect 2044 1896 2096 1902
rect 2044 1838 2096 1844
rect 2148 1766 2176 2246
rect 2136 1760 2188 1766
rect 2136 1702 2188 1708
rect 2240 800 2268 2926
rect 2412 2848 2464 2854
rect 2410 2816 2412 2825
rect 2504 2848 2556 2854
rect 2464 2816 2466 2825
rect 2504 2790 2556 2796
rect 2410 2751 2466 2760
rect 2516 2446 2544 2790
rect 2608 2514 2636 3046
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 2700 800 2728 2926
rect 2884 2650 2912 3538
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 1306 232 1362 241
rect 1306 167 1362 176
rect 1398 0 1454 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 2976 649 3004 3998
rect 3160 2990 3188 5646
rect 3238 5607 3294 5616
rect 3252 3398 3280 5607
rect 3344 4010 3372 6054
rect 3528 5166 3556 6122
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3620 5012 3648 6695
rect 3712 6458 3740 7142
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6497 3832 6598
rect 3790 6488 3846 6497
rect 3700 6452 3752 6458
rect 3790 6423 3846 6432
rect 3700 6394 3752 6400
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3804 6118 3832 6326
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3792 6112 3844 6118
rect 3988 6100 4016 7686
rect 4080 7410 4108 7958
rect 4158 7919 4214 7928
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4172 7546 4200 7822
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4080 6905 4108 7210
rect 4172 6934 4200 7278
rect 4160 6928 4212 6934
rect 4066 6896 4122 6905
rect 4160 6870 4212 6876
rect 4066 6831 4122 6840
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6254 4108 6598
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 3988 6072 4108 6100
rect 3792 6054 3844 6060
rect 3712 5914 3740 6054
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3804 5574 3832 6054
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3988 5778 4016 5850
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3712 5273 3740 5510
rect 3790 5400 3846 5409
rect 4080 5370 4108 6072
rect 4172 6066 4200 6870
rect 4264 6458 4292 7890
rect 4356 7392 4384 8266
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5184 8090 5212 13926
rect 5356 13864 5408 13870
rect 5262 13832 5318 13841
rect 5356 13806 5408 13812
rect 5262 13767 5318 13776
rect 5276 13530 5304 13767
rect 5368 13705 5396 13806
rect 5354 13696 5410 13705
rect 5354 13631 5410 13640
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5276 12646 5304 13466
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5368 13025 5396 13398
rect 5354 13016 5410 13025
rect 5354 12951 5410 12960
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5368 12374 5396 12951
rect 5460 12424 5488 15302
rect 5552 14958 5580 15914
rect 5644 15502 5672 16594
rect 5736 15638 5764 16934
rect 5828 16046 5856 17138
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 5920 15688 5948 17292
rect 6012 16726 6040 17614
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6012 15706 6040 15846
rect 5828 15660 5948 15688
rect 6000 15700 6052 15706
rect 5724 15632 5776 15638
rect 5724 15574 5776 15580
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5644 15162 5672 15438
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5552 13569 5580 14282
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5538 13560 5594 13569
rect 5538 13495 5594 13504
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5552 12646 5580 13126
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5460 12396 5580 12424
rect 5356 12368 5408 12374
rect 5552 12345 5580 12396
rect 5356 12310 5408 12316
rect 5538 12336 5594 12345
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5448 12300 5500 12306
rect 5538 12271 5594 12280
rect 5448 12242 5500 12248
rect 5276 12050 5304 12242
rect 5354 12200 5410 12209
rect 5354 12135 5356 12144
rect 5408 12135 5410 12144
rect 5356 12106 5408 12112
rect 5276 12022 5396 12050
rect 5262 11928 5318 11937
rect 5262 11863 5318 11872
rect 5276 11014 5304 11863
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5276 10674 5304 10746
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5276 10062 5304 10610
rect 5368 10470 5396 12022
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5276 9450 5304 9998
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5368 9330 5396 10406
rect 5460 9518 5488 12242
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5552 11762 5580 12038
rect 5644 11898 5672 13874
rect 5736 13569 5764 14350
rect 5828 14226 5856 15660
rect 6000 15642 6052 15648
rect 5908 15564 5960 15570
rect 5960 15524 6040 15552
rect 5908 15506 5960 15512
rect 6012 14822 6040 15524
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 5828 14198 5948 14226
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5722 13560 5778 13569
rect 5722 13495 5778 13504
rect 5736 12986 5764 13495
rect 5828 13394 5856 14010
rect 5920 13870 5948 14198
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 5920 13530 5948 13670
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5906 13424 5962 13433
rect 5816 13388 5868 13394
rect 5906 13359 5962 13368
rect 5816 13330 5868 13336
rect 5920 13326 5948 13359
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5814 13152 5870 13161
rect 5814 13087 5870 13096
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5828 12850 5856 13087
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5736 12442 5764 12786
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11286 5580 11494
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5644 10810 5672 11562
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5630 10704 5686 10713
rect 5630 10639 5686 10648
rect 5644 10606 5672 10639
rect 5736 10606 5764 10950
rect 5632 10600 5684 10606
rect 5538 10568 5594 10577
rect 5632 10542 5684 10548
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5538 10503 5540 10512
rect 5592 10503 5594 10512
rect 5540 10474 5592 10480
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5276 9302 5396 9330
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4802 7576 4858 7585
rect 4724 7520 4802 7528
rect 4724 7511 4858 7520
rect 4724 7500 4844 7511
rect 4356 7364 4476 7392
rect 4448 7290 4476 7364
rect 4448 7262 4660 7290
rect 4632 7206 4660 7262
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4540 7002 4568 7142
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4528 6996 4580 7002
rect 4528 6938 4580 6944
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4252 6248 4304 6254
rect 4250 6216 4252 6225
rect 4304 6216 4306 6225
rect 4250 6151 4306 6160
rect 4172 6038 4292 6066
rect 4158 5944 4214 5953
rect 4158 5879 4214 5888
rect 3790 5335 3792 5344
rect 3844 5335 3846 5344
rect 4068 5364 4120 5370
rect 3792 5306 3844 5312
rect 4068 5306 4120 5312
rect 3698 5264 3754 5273
rect 3698 5199 3754 5208
rect 3976 5228 4028 5234
rect 4172 5216 4200 5879
rect 4264 5778 4292 6038
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4356 5624 4384 6938
rect 4632 6905 4660 7142
rect 4618 6896 4674 6905
rect 4724 6866 4752 7500
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4618 6831 4674 6840
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4816 6390 4844 7346
rect 4436 6384 4488 6390
rect 4804 6384 4856 6390
rect 4436 6326 4488 6332
rect 4802 6352 4804 6361
rect 4856 6352 4858 6361
rect 4028 5188 4200 5216
rect 4264 5596 4384 5624
rect 3976 5170 4028 5176
rect 4264 5166 4292 5596
rect 4448 5556 4476 6326
rect 4802 6287 4858 6296
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 4816 5778 4844 6122
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4356 5528 4476 5556
rect 4356 5352 4384 5528
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4356 5324 4660 5352
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 3528 4984 3648 5012
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3436 3738 3464 4558
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3528 3618 3556 4984
rect 3896 4865 3924 5034
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3882 4856 3938 4865
rect 3882 4791 3938 4800
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3344 3590 3556 3618
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 3238 2952 3294 2961
rect 3238 2887 3240 2896
rect 3292 2887 3294 2896
rect 3240 2858 3292 2864
rect 3344 2650 3372 3590
rect 3620 3534 3648 3946
rect 3804 3641 3832 4422
rect 3988 4078 4016 4966
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 3790 3632 3846 3641
rect 3790 3567 3846 3576
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3436 2854 3464 3334
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 3528 2650 3556 3062
rect 3620 3058 3648 3470
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3620 2446 3648 2994
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3056 1828 3108 1834
rect 3056 1770 3108 1776
rect 3068 800 3096 1770
rect 3712 1442 3740 3130
rect 3804 3058 3832 3567
rect 3988 3534 4016 3878
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3896 2582 3924 3470
rect 4172 2990 4200 3878
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4172 2582 4200 2790
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 3792 2372 3844 2378
rect 3844 2332 3924 2360
rect 3792 2314 3844 2320
rect 3528 1414 3740 1442
rect 3528 800 3556 1414
rect 3896 800 3924 2332
rect 4264 1465 4292 4422
rect 4356 3942 4384 4558
rect 4632 4468 4660 5324
rect 4816 5234 4844 5714
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4690 4752 4966
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4632 4440 4844 4468
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4712 4208 4764 4214
rect 4618 4176 4674 4185
rect 4712 4150 4764 4156
rect 4618 4111 4674 4120
rect 4632 4078 4660 4111
rect 4436 4072 4488 4078
rect 4620 4072 4672 4078
rect 4488 4032 4568 4060
rect 4436 4014 4488 4020
rect 4344 3936 4396 3942
rect 4436 3936 4488 3942
rect 4344 3878 4396 3884
rect 4434 3904 4436 3913
rect 4488 3904 4490 3913
rect 4356 3738 4384 3878
rect 4434 3839 4490 3848
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4540 3602 4568 4032
rect 4620 4014 4672 4020
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4632 3380 4660 4014
rect 4724 3670 4752 4150
rect 4712 3664 4764 3670
rect 4710 3632 4712 3641
rect 4764 3632 4766 3641
rect 4710 3567 4766 3576
rect 4356 3352 4660 3380
rect 4250 1456 4306 1465
rect 4250 1391 4306 1400
rect 4356 800 4384 3352
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4724 2582 4752 2926
rect 4816 2650 4844 4440
rect 4908 3602 4936 7890
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5000 6322 5028 7482
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5092 6186 5120 7482
rect 5184 6458 5212 7822
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5184 6066 5212 6122
rect 5000 6038 5212 6066
rect 5000 5234 5028 6038
rect 5172 5568 5224 5574
rect 5092 5528 5172 5556
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5000 4554 5028 5170
rect 5092 5166 5120 5528
rect 5172 5510 5224 5516
rect 5276 5386 5304 9302
rect 5552 8430 5580 10066
rect 5828 10062 5856 12786
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 5920 12345 5948 12718
rect 5906 12336 5962 12345
rect 5906 12271 5962 12280
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 10810 5948 11494
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 6012 10470 6040 14758
rect 6104 11257 6132 18022
rect 6196 17678 6224 18770
rect 6274 18456 6330 18465
rect 6274 18391 6330 18400
rect 6288 18222 6316 18391
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6288 17746 6316 18022
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6196 16658 6224 17138
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6196 15502 6224 16390
rect 6288 16046 6316 16594
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6196 14657 6224 15438
rect 6288 15434 6316 15846
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6182 14648 6238 14657
rect 6182 14583 6238 14592
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 13938 6224 14350
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6196 13841 6224 13874
rect 6182 13832 6238 13841
rect 6182 13767 6238 13776
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6196 12782 6224 13330
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6090 11248 6146 11257
rect 6090 11183 6146 11192
rect 6104 11082 6132 11183
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 10198 6040 10406
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5644 8634 5672 9318
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5354 7576 5410 7585
rect 5354 7511 5410 7520
rect 5368 7410 5396 7511
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5460 7290 5488 8230
rect 5644 8022 5672 8570
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5736 7868 5764 9114
rect 5920 9042 5948 9318
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5828 8430 5856 8910
rect 6012 8634 6040 9998
rect 6104 9518 6132 9998
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6092 9376 6144 9382
rect 6196 9364 6224 12582
rect 6288 10282 6316 14486
rect 6380 10418 6408 18924
rect 6460 18906 6512 18912
rect 6472 18834 6500 18906
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6472 18222 6500 18362
rect 6460 18216 6512 18222
rect 6460 18158 6512 18164
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6472 17882 6500 18022
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6564 17762 6592 19314
rect 6656 18834 6684 19468
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6656 18290 6684 18770
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6748 17882 6776 20266
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6840 19174 6868 19858
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6932 18970 6960 19654
rect 7024 19514 7052 19994
rect 7104 19984 7156 19990
rect 7104 19926 7156 19932
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 7010 19408 7066 19417
rect 7010 19343 7066 19352
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 6932 18630 6960 18906
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6840 18465 6868 18566
rect 6826 18456 6882 18465
rect 6826 18391 6882 18400
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6932 17882 6960 18022
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6564 17734 6868 17762
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6472 15706 6500 16050
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6564 15638 6592 17070
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6552 15088 6604 15094
rect 6552 15030 6604 15036
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6472 12986 6500 14418
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6564 12481 6592 15030
rect 6656 14822 6684 15914
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6748 15162 6776 15438
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6748 14346 6776 15098
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6656 13258 6684 13874
rect 6840 13852 6868 17734
rect 6920 17060 6972 17066
rect 6920 17002 6972 17008
rect 6932 16454 6960 17002
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6932 16114 6960 16390
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6932 14618 6960 15846
rect 7024 15042 7052 19343
rect 7116 18970 7144 19926
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7208 18698 7236 20198
rect 7300 20058 7328 20266
rect 7288 20052 7340 20058
rect 7288 19994 7340 20000
rect 7300 19825 7328 19994
rect 7484 19990 7512 22200
rect 7852 20398 7880 22200
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 8116 20392 8168 20398
rect 8220 20380 8248 22200
rect 8300 20392 8352 20398
rect 8220 20352 8300 20380
rect 8116 20334 8168 20340
rect 8588 20380 8616 22200
rect 8852 20800 8904 20806
rect 8852 20742 8904 20748
rect 8760 20392 8812 20398
rect 8588 20352 8760 20380
rect 8300 20334 8352 20340
rect 8760 20334 8812 20340
rect 7748 20256 7800 20262
rect 8128 20244 8156 20334
rect 8128 20216 8248 20244
rect 7748 20198 7800 20204
rect 7472 19984 7524 19990
rect 7472 19926 7524 19932
rect 7380 19848 7432 19854
rect 7286 19816 7342 19825
rect 7380 19790 7432 19796
rect 7286 19751 7342 19760
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7208 17542 7236 17818
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7300 16969 7328 19654
rect 7392 17542 7420 19790
rect 7760 19718 7788 20198
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7472 19236 7524 19242
rect 7472 19178 7524 19184
rect 7484 17660 7512 19178
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7576 18766 7604 19110
rect 7668 18970 7696 19654
rect 8128 19242 8156 19790
rect 8220 19689 8248 20216
rect 8312 19990 8340 20334
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 8300 19712 8352 19718
rect 8206 19680 8262 19689
rect 8300 19654 8352 19660
rect 8206 19615 8262 19624
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 8220 18426 8248 18770
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7576 17785 7604 17818
rect 7562 17776 7618 17785
rect 7562 17711 7618 17720
rect 7564 17672 7616 17678
rect 7484 17632 7564 17660
rect 7564 17614 7616 17620
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 17338 7420 17478
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7576 17202 7604 17614
rect 7668 17338 7696 18022
rect 7760 17882 7788 18158
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 7748 17672 7800 17678
rect 7746 17640 7748 17649
rect 7800 17640 7802 17649
rect 7746 17575 7802 17584
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 8220 17241 8248 17818
rect 8206 17232 8262 17241
rect 7564 17196 7616 17202
rect 8206 17167 8262 17176
rect 7564 17138 7616 17144
rect 7286 16960 7342 16969
rect 7286 16895 7342 16904
rect 7576 16794 7604 17138
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7300 16572 7328 16730
rect 7300 16544 7420 16572
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7208 15162 7236 15438
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7024 15014 7144 15042
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 7024 14482 7052 14894
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 6748 13824 6868 13852
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6656 12850 6684 13194
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6642 12744 6698 12753
rect 6642 12679 6698 12688
rect 6656 12646 6684 12679
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6550 12472 6606 12481
rect 6748 12434 6776 13824
rect 6826 13696 6882 13705
rect 6826 13631 6882 13640
rect 6840 13394 6868 13631
rect 6918 13560 6974 13569
rect 6918 13495 6974 13504
rect 6932 13462 6960 13495
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6550 12407 6606 12416
rect 6656 12406 6776 12434
rect 6460 12368 6512 12374
rect 6460 12310 6512 12316
rect 6472 11898 6500 12310
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6472 10538 6500 11834
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6564 11286 6592 11698
rect 6656 11558 6684 12406
rect 6734 12336 6790 12345
rect 6840 12306 6868 13330
rect 7024 12986 7052 14418
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7116 12866 7144 15014
rect 7392 14822 7420 16544
rect 8312 15994 8340 19654
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 8404 16726 8432 17206
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8404 16114 8432 16662
rect 8496 16153 8524 20198
rect 8574 19816 8630 19825
rect 8574 19751 8630 19760
rect 8588 18222 8616 19751
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8576 17536 8628 17542
rect 8574 17504 8576 17513
rect 8628 17504 8630 17513
rect 8574 17439 8630 17448
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8588 16794 8616 17070
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8588 16561 8616 16730
rect 8574 16552 8630 16561
rect 8574 16487 8630 16496
rect 8482 16144 8538 16153
rect 8392 16108 8444 16114
rect 8482 16079 8538 16088
rect 8392 16050 8444 16056
rect 7656 15972 7708 15978
rect 8312 15966 8524 15994
rect 7656 15914 7708 15920
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7300 14618 7328 14758
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7208 13530 7236 14350
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 6932 12838 7144 12866
rect 6734 12271 6790 12280
rect 6828 12300 6880 12306
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6564 10674 6592 10950
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6460 10532 6512 10538
rect 6460 10474 6512 10480
rect 6380 10390 6592 10418
rect 6458 10296 6514 10305
rect 6288 10254 6408 10282
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6144 9336 6224 9364
rect 6092 9318 6144 9324
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6104 8514 6132 9318
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6012 8486 6132 8514
rect 6196 8498 6224 8978
rect 6288 8566 6316 10066
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6184 8492 6236 8498
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5368 7262 5488 7290
rect 5552 7840 5764 7868
rect 5368 6905 5396 7262
rect 5552 7206 5580 7840
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5644 7018 5672 7142
rect 5460 6990 5672 7018
rect 5354 6896 5410 6905
rect 5354 6831 5410 6840
rect 5368 6730 5396 6831
rect 5365 6724 5417 6730
rect 5365 6666 5417 6672
rect 5460 5914 5488 6990
rect 5540 6860 5592 6866
rect 5592 6820 5672 6848
rect 5540 6802 5592 6808
rect 5538 6760 5594 6769
rect 5538 6695 5594 6704
rect 5552 6662 5580 6695
rect 5540 6656 5592 6662
rect 5644 6633 5672 6820
rect 5828 6662 5856 8230
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5920 7177 5948 7210
rect 5906 7168 5962 7177
rect 5906 7103 5962 7112
rect 5816 6656 5868 6662
rect 5540 6598 5592 6604
rect 5630 6624 5686 6633
rect 5816 6598 5868 6604
rect 5630 6559 5686 6568
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5552 5953 5580 6258
rect 5538 5944 5594 5953
rect 5448 5908 5500 5914
rect 5538 5879 5540 5888
rect 5448 5850 5500 5856
rect 5592 5879 5594 5888
rect 5540 5850 5592 5856
rect 5644 5794 5672 6559
rect 6012 6497 6040 8486
rect 6184 8434 6236 8440
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6104 7002 6132 7278
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 7041 6316 7142
rect 6274 7032 6330 7041
rect 6092 6996 6144 7002
rect 6274 6967 6330 6976
rect 6092 6938 6144 6944
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 5998 6488 6054 6497
rect 5724 6452 5776 6458
rect 5998 6423 6054 6432
rect 5724 6394 5776 6400
rect 5184 5358 5304 5386
rect 5552 5766 5672 5794
rect 5736 5778 5764 6394
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5828 5914 5856 6054
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 6012 5828 6040 6423
rect 5920 5800 6040 5828
rect 5724 5772 5776 5778
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 5092 4146 5120 4966
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4988 3936 5040 3942
rect 4986 3904 4988 3913
rect 5040 3904 5042 3913
rect 4986 3839 5042 3848
rect 4986 3768 5042 3777
rect 4986 3703 5042 3712
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4908 2514 4936 2858
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 4804 2304 4856 2310
rect 4802 2272 4804 2281
rect 4856 2272 4858 2281
rect 4421 2204 4717 2224
rect 4802 2207 4858 2216
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4908 1834 4936 2450
rect 4896 1828 4948 1834
rect 4896 1770 4948 1776
rect 5000 1714 5028 3703
rect 5092 3194 5120 4082
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5184 2990 5212 5358
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5276 4622 5304 5170
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5276 4146 5304 4558
rect 5354 4312 5410 4321
rect 5354 4247 5410 4256
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5276 3670 5304 4082
rect 5368 3942 5396 4247
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5460 3738 5488 4966
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5276 2378 5304 3606
rect 5354 3360 5410 3369
rect 5354 3295 5410 3304
rect 5368 2825 5396 3295
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5354 2816 5410 2825
rect 5354 2751 5410 2760
rect 5460 2514 5488 3062
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 5460 1850 5488 2450
rect 5552 2417 5580 5766
rect 5724 5714 5776 5720
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5644 2650 5672 4694
rect 5736 4486 5764 5714
rect 5814 5672 5870 5681
rect 5814 5607 5870 5616
rect 5828 5574 5856 5607
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5920 5386 5948 5800
rect 5998 5672 6054 5681
rect 5998 5607 6054 5616
rect 5828 5358 5948 5386
rect 5828 5166 5856 5358
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5828 4593 5856 4626
rect 5814 4584 5870 4593
rect 5814 4519 5870 4528
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5814 4448 5870 4457
rect 5814 4383 5870 4392
rect 5828 4298 5856 4383
rect 5736 4270 5856 4298
rect 5736 4010 5764 4270
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5736 3777 5764 3946
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5722 3768 5778 3777
rect 5722 3703 5778 3712
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 5736 3194 5764 3606
rect 5828 3194 5856 3878
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5828 2582 5856 2790
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 5920 2428 5948 5102
rect 6012 4842 6040 5607
rect 6104 4978 6132 6802
rect 6182 6760 6238 6769
rect 6182 6695 6238 6704
rect 6196 6225 6224 6695
rect 6182 6216 6238 6225
rect 6182 6151 6238 6160
rect 6182 5808 6238 5817
rect 6182 5743 6184 5752
rect 6236 5743 6238 5752
rect 6184 5714 6236 5720
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6274 5536 6330 5545
rect 6196 5098 6224 5510
rect 6274 5471 6330 5480
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 6104 4950 6224 4978
rect 6012 4814 6132 4842
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6012 3534 6040 4082
rect 6104 3670 6132 4814
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6104 3126 6132 3470
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 6196 2825 6224 4950
rect 6288 4826 6316 5471
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6274 4584 6330 4593
rect 6274 4519 6330 4528
rect 6182 2816 6238 2825
rect 6182 2751 6238 2760
rect 6288 2650 6316 4519
rect 6380 3126 6408 10254
rect 6458 10231 6460 10240
rect 6512 10231 6514 10240
rect 6460 10202 6512 10208
rect 6472 6338 6500 10202
rect 6564 9722 6592 10390
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6564 6798 6592 9658
rect 6656 9654 6684 11086
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6656 8888 6684 9454
rect 6748 9353 6776 12271
rect 6828 12242 6880 12248
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 10169 6868 11494
rect 6932 10198 6960 12838
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7010 12608 7066 12617
rect 7010 12543 7066 12552
rect 6920 10192 6972 10198
rect 6826 10160 6882 10169
rect 6920 10134 6972 10140
rect 6826 10095 6882 10104
rect 6840 9625 6868 10095
rect 7024 10010 7052 12543
rect 7116 12170 7144 12650
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7208 11694 7236 12038
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 7116 10742 7144 11222
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 6932 9982 7052 10010
rect 6826 9616 6882 9625
rect 6826 9551 6882 9560
rect 6734 9344 6790 9353
rect 6734 9279 6790 9288
rect 6932 9110 6960 9982
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7024 9625 7052 9862
rect 7010 9616 7066 9625
rect 7010 9551 7066 9560
rect 7012 9512 7064 9518
rect 7010 9480 7012 9489
rect 7064 9480 7066 9489
rect 7010 9415 7066 9424
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6656 8860 6776 8888
rect 6748 8072 6776 8860
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6840 8430 6868 8774
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6932 8129 6960 8774
rect 7024 8430 7052 9318
rect 7116 9178 7144 10066
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 9382 7236 9998
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7208 9058 7236 9318
rect 7116 9030 7236 9058
rect 7116 8498 7144 9030
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 6918 8120 6974 8129
rect 6828 8084 6880 8090
rect 6748 8044 6828 8072
rect 7116 8090 7144 8298
rect 6918 8055 6974 8064
rect 7104 8084 7156 8090
rect 6828 8026 6880 8032
rect 7104 8026 7156 8032
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6748 7002 6776 7482
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 6642 6896 6698 6905
rect 6642 6831 6698 6840
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6472 6310 6592 6338
rect 6656 6322 6684 6831
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6748 6458 6776 6666
rect 6840 6458 6868 7686
rect 6918 7576 6974 7585
rect 6918 7511 6974 7520
rect 6932 7410 6960 7511
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6918 7304 6974 7313
rect 6918 7239 6974 7248
rect 7012 7268 7064 7274
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6458 6216 6514 6225
rect 6564 6202 6592 6310
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6734 6216 6790 6225
rect 6564 6174 6684 6202
rect 6458 6151 6514 6160
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 5538 2408 5594 2417
rect 5538 2343 5594 2352
rect 5644 2400 5948 2428
rect 4816 1686 5028 1714
rect 5184 1822 5488 1850
rect 4816 800 4844 1686
rect 5184 800 5212 1822
rect 5644 800 5672 2400
rect 6012 2106 6040 2450
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 6000 2100 6052 2106
rect 6000 2042 6052 2048
rect 6104 2038 6132 2382
rect 6472 2038 6500 6151
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6564 2514 6592 6054
rect 6656 3942 6684 6174
rect 6734 6151 6790 6160
rect 6748 5914 6776 6151
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6840 5710 6868 6394
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6932 5574 6960 7239
rect 7012 7210 7064 7216
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6734 5400 6790 5409
rect 6734 5335 6790 5344
rect 6920 5364 6972 5370
rect 6748 5030 6776 5335
rect 6920 5306 6972 5312
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6748 4214 6776 4422
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3398 6776 3878
rect 6840 3466 6868 4966
rect 6932 3534 6960 5306
rect 7024 5234 7052 7210
rect 7116 6798 7144 7346
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7010 4720 7066 4729
rect 7116 4690 7144 6598
rect 7208 6322 7236 8434
rect 7300 8378 7328 13806
rect 7392 12434 7420 14758
rect 7562 14648 7618 14657
rect 7562 14583 7618 14592
rect 7576 14550 7604 14583
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7484 13938 7512 14282
rect 7668 14074 7696 15914
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 7760 15706 7788 15846
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8220 15094 8248 15302
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7760 13954 7788 14962
rect 7838 14920 7894 14929
rect 7838 14855 7840 14864
rect 7892 14855 7894 14864
rect 7840 14826 7892 14832
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7668 13926 7788 13954
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7576 13433 7604 13670
rect 7668 13462 7696 13926
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7656 13456 7708 13462
rect 7562 13424 7618 13433
rect 7656 13398 7708 13404
rect 7562 13359 7618 13368
rect 7562 12880 7618 12889
rect 7562 12815 7564 12824
rect 7616 12815 7618 12824
rect 7564 12786 7616 12792
rect 7392 12406 7512 12434
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7392 12073 7420 12242
rect 7378 12064 7434 12073
rect 7378 11999 7434 12008
rect 7484 11914 7512 12406
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7392 11886 7512 11914
rect 7392 11529 7420 11886
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7378 11520 7434 11529
rect 7378 11455 7434 11464
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7392 11121 7420 11290
rect 7484 11218 7512 11562
rect 7576 11354 7604 12242
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7378 11112 7434 11121
rect 7378 11047 7434 11056
rect 7392 10810 7420 11047
rect 7668 10826 7696 13398
rect 7760 12714 7788 13806
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7840 12776 7892 12782
rect 8220 12753 8248 13670
rect 8404 13394 8432 15846
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 12782 8340 13126
rect 8300 12776 8352 12782
rect 7840 12718 7892 12724
rect 8206 12744 8262 12753
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7852 12628 7880 12718
rect 8300 12718 8352 12724
rect 8206 12679 8262 12688
rect 7821 12600 7880 12628
rect 8208 12640 8260 12646
rect 7821 12434 7849 12600
rect 8208 12582 8260 12588
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 7821 12406 7880 12434
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 10849 7788 12038
rect 7852 11830 7880 12406
rect 8024 12368 8076 12374
rect 7944 12328 8024 12356
rect 7944 11898 7972 12328
rect 8024 12310 8076 12316
rect 8114 12336 8170 12345
rect 8114 12271 8170 12280
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 8036 11626 8064 12174
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 8128 11540 8156 12271
rect 8220 12238 8248 12582
rect 8312 12306 8340 12718
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8312 11762 8340 12242
rect 8404 12073 8432 13330
rect 8496 12424 8524 15966
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8588 14822 8616 15506
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8588 14278 8616 14758
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8588 13258 8616 13466
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8574 13016 8630 13025
rect 8680 12986 8708 20198
rect 8772 20058 8800 20334
rect 8864 20330 8892 20742
rect 8956 20516 8984 22200
rect 9036 20528 9088 20534
rect 8956 20488 9036 20516
rect 9036 20470 9088 20476
rect 9416 20398 9444 22200
rect 9784 20398 9812 22200
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 8852 20324 8904 20330
rect 8852 20266 8904 20272
rect 9416 20058 9444 20334
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 9496 20256 9548 20262
rect 9496 20198 9548 20204
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9404 19712 9456 19718
rect 9126 19680 9182 19689
rect 9404 19654 9456 19660
rect 9126 19615 9182 19624
rect 8852 19236 8904 19242
rect 8852 19178 8904 19184
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 8864 18601 8892 19178
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8850 18592 8906 18601
rect 8850 18527 8906 18536
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8574 12951 8630 12960
rect 8668 12980 8720 12986
rect 8588 12646 8616 12951
rect 8668 12922 8720 12928
rect 8680 12753 8708 12922
rect 8666 12744 8722 12753
rect 8666 12679 8722 12688
rect 8576 12640 8628 12646
rect 8772 12617 8800 17750
rect 8864 17134 8892 18226
rect 8956 18154 8984 19110
rect 9048 18698 9076 19178
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 9048 18222 9076 18634
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 9048 17338 9076 18158
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 8956 16522 8984 16934
rect 9048 16590 9076 17274
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 8956 15881 8984 16458
rect 9048 15978 9076 16526
rect 9036 15972 9088 15978
rect 9036 15914 9088 15920
rect 8942 15872 8998 15881
rect 8942 15807 8998 15816
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 8852 14544 8904 14550
rect 8852 14486 8904 14492
rect 8864 14346 8892 14486
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8850 13968 8906 13977
rect 8850 13903 8906 13912
rect 8864 13462 8892 13903
rect 8852 13456 8904 13462
rect 8852 13398 8904 13404
rect 8576 12582 8628 12588
rect 8758 12608 8814 12617
rect 8758 12543 8814 12552
rect 8864 12481 8892 13398
rect 8850 12472 8906 12481
rect 8496 12396 8708 12424
rect 8850 12407 8906 12416
rect 8482 12336 8538 12345
rect 8482 12271 8538 12280
rect 8390 12064 8446 12073
rect 8390 11999 8446 12008
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8300 11552 8352 11558
rect 8128 11512 8248 11540
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7484 10798 7696 10826
rect 7746 10840 7802 10849
rect 7484 9704 7512 10798
rect 7746 10775 7802 10784
rect 7564 10736 7616 10742
rect 7562 10704 7564 10713
rect 7616 10704 7618 10713
rect 8036 10674 8064 10950
rect 7562 10639 7618 10648
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7564 10464 7616 10470
rect 7562 10432 7564 10441
rect 7616 10432 7618 10441
rect 7562 10367 7618 10376
rect 7668 10062 7696 10610
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7392 9676 7512 9704
rect 7392 8498 7420 9676
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7484 8906 7512 9522
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7300 8350 7420 8378
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 8090 7328 8230
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7392 6458 7420 8350
rect 7484 7886 7512 8842
rect 7576 8090 7604 9862
rect 7760 9432 7788 10474
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 8220 10266 8248 11512
rect 8300 11494 8352 11500
rect 8312 11082 8340 11494
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8298 10976 8354 10985
rect 8298 10911 8354 10920
rect 8312 10266 8340 10911
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8298 10024 8354 10033
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7930 9752 7986 9761
rect 7930 9687 7986 9696
rect 7668 9404 7788 9432
rect 7668 9092 7696 9404
rect 7944 9364 7972 9687
rect 8036 9489 8064 9862
rect 8022 9480 8078 9489
rect 8220 9450 8248 9998
rect 8298 9959 8354 9968
rect 8312 9926 8340 9959
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8298 9480 8354 9489
rect 8022 9415 8078 9424
rect 8208 9444 8260 9450
rect 8298 9415 8354 9424
rect 8208 9386 8260 9392
rect 7821 9336 7972 9364
rect 7821 9160 7849 9336
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 7821 9132 7972 9160
rect 7668 9064 7788 9092
rect 7760 8498 7788 9064
rect 7944 9042 7972 9132
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 8128 8276 8156 8978
rect 8220 8974 8248 9386
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 8378 8248 8774
rect 8312 8498 8340 9415
rect 8404 8673 8432 11999
rect 8496 9994 8524 12271
rect 8574 12064 8630 12073
rect 8574 11999 8630 12008
rect 8588 11694 8616 11999
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8588 11354 8616 11494
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8390 8664 8446 8673
rect 8390 8599 8446 8608
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8220 8350 8340 8378
rect 8128 8248 8248 8276
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7760 7750 7788 7958
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7656 7404 7708 7410
rect 7760 7392 7788 7686
rect 7708 7364 7788 7392
rect 7656 7346 7708 7352
rect 7472 7200 7524 7206
rect 7524 7160 7604 7188
rect 7472 7142 7524 7148
rect 7576 6769 7604 7160
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8220 7002 8248 8248
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8312 6882 8340 8350
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8404 8090 8432 8230
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8496 7970 8524 9930
rect 8588 8974 8616 11018
rect 8680 10985 8708 12396
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8772 11665 8800 12038
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8758 11656 8814 11665
rect 8758 11591 8814 11600
rect 8864 11558 8892 11766
rect 8760 11552 8812 11558
rect 8758 11520 8760 11529
rect 8852 11552 8904 11558
rect 8812 11520 8814 11529
rect 8852 11494 8904 11500
rect 8758 11455 8814 11464
rect 8666 10976 8722 10985
rect 8666 10911 8722 10920
rect 8850 10840 8906 10849
rect 8850 10775 8906 10784
rect 8760 10736 8812 10742
rect 8680 10684 8760 10690
rect 8680 10678 8812 10684
rect 8680 10662 8800 10678
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8404 7942 8524 7970
rect 8576 7948 8628 7954
rect 8404 7546 8432 7942
rect 8576 7890 8628 7896
rect 8588 7546 8616 7890
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8036 6854 8340 6882
rect 8576 6928 8628 6934
rect 8680 6916 8708 10662
rect 8864 10606 8892 10775
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8852 10464 8904 10470
rect 8758 10432 8814 10441
rect 8852 10406 8904 10412
rect 8758 10367 8814 10376
rect 8772 9110 8800 10367
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8772 7449 8800 8910
rect 8758 7440 8814 7449
rect 8758 7375 8814 7384
rect 8628 6888 8708 6916
rect 8576 6870 8628 6876
rect 7656 6792 7708 6798
rect 7562 6760 7618 6769
rect 7656 6734 7708 6740
rect 7562 6695 7618 6704
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 7378 6352 7434 6361
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 5681 7236 6258
rect 7300 6254 7328 6326
rect 7562 6352 7618 6361
rect 7472 6316 7524 6322
rect 7434 6296 7472 6304
rect 7378 6287 7472 6296
rect 7392 6276 7472 6287
rect 7562 6287 7618 6296
rect 7472 6258 7524 6264
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7576 6168 7604 6287
rect 7392 6140 7604 6168
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7194 5672 7250 5681
rect 7194 5607 7250 5616
rect 7196 5024 7248 5030
rect 7300 5001 7328 5714
rect 7392 5137 7420 6140
rect 7562 5808 7618 5817
rect 7668 5794 7696 6734
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7852 6390 7880 6598
rect 7840 6384 7892 6390
rect 7746 6352 7802 6361
rect 7840 6326 7892 6332
rect 7746 6287 7802 6296
rect 7760 6254 7788 6287
rect 7748 6248 7800 6254
rect 8036 6225 8064 6854
rect 8392 6792 8444 6798
rect 8312 6752 8392 6780
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 7748 6190 7800 6196
rect 8022 6216 8078 6225
rect 8022 6151 8078 6160
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7618 5766 7696 5794
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7562 5743 7618 5752
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7470 5400 7526 5409
rect 7470 5335 7526 5344
rect 7378 5128 7434 5137
rect 7484 5098 7512 5335
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7378 5063 7434 5072
rect 7472 5092 7524 5098
rect 7196 4966 7248 4972
rect 7286 4992 7342 5001
rect 7010 4655 7066 4664
rect 7104 4684 7156 4690
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6656 2922 6684 3130
rect 6644 2916 6696 2922
rect 6696 2876 6868 2904
rect 6644 2858 6696 2864
rect 6734 2816 6790 2825
rect 6734 2751 6790 2760
rect 6748 2650 6776 2751
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6092 2032 6144 2038
rect 6092 1974 6144 1980
rect 6460 2032 6512 2038
rect 6460 1974 6512 1980
rect 6564 1834 6592 2450
rect 6000 1828 6052 1834
rect 6000 1770 6052 1776
rect 6552 1828 6604 1834
rect 6552 1770 6604 1776
rect 6012 800 6040 1770
rect 6460 1760 6512 1766
rect 6460 1702 6512 1708
rect 6472 800 6500 1702
rect 6840 800 6868 2876
rect 7024 2650 7052 4655
rect 7104 4626 7156 4632
rect 7208 4282 7236 4966
rect 7286 4927 7342 4936
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7300 4729 7328 4762
rect 7286 4720 7342 4729
rect 7286 4655 7342 4664
rect 7392 4622 7420 5063
rect 7472 5034 7524 5040
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7116 3126 7144 3538
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7194 2544 7250 2553
rect 7194 2479 7196 2488
rect 7248 2479 7250 2488
rect 7196 2450 7248 2456
rect 7208 1766 7236 2450
rect 7196 1760 7248 1766
rect 7196 1702 7248 1708
rect 7300 800 7328 4558
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7392 4078 7420 4422
rect 7576 4282 7604 5170
rect 7668 4758 7696 5510
rect 7944 5273 7972 5782
rect 8024 5772 8076 5778
rect 8220 5760 8248 6598
rect 8076 5732 8248 5760
rect 8024 5714 8076 5720
rect 8208 5568 8260 5574
rect 8022 5536 8078 5545
rect 8208 5510 8260 5516
rect 8022 5471 8078 5480
rect 7930 5264 7986 5273
rect 7930 5199 7986 5208
rect 8036 5166 8064 5471
rect 8220 5234 8248 5510
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4826 7788 4966
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 8220 4706 8248 5170
rect 8312 5030 8340 6752
rect 8392 6734 8444 6740
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8496 6633 8524 6666
rect 8482 6624 8538 6633
rect 8482 6559 8538 6568
rect 8680 6390 8708 6888
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8220 4678 8340 4706
rect 8312 4622 8340 4678
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7484 3670 7512 4014
rect 8220 4010 8248 4558
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 8220 3602 8248 3946
rect 8312 3738 8340 4558
rect 8404 4078 8432 6054
rect 8588 5710 8616 6258
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8496 3618 8524 5510
rect 8680 5273 8708 5578
rect 8666 5264 8722 5273
rect 8666 5199 8722 5208
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8588 4457 8616 4966
rect 8574 4448 8630 4457
rect 8574 4383 8630 4392
rect 8680 4185 8708 5102
rect 8772 4729 8800 7375
rect 8758 4720 8814 4729
rect 8758 4655 8814 4664
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8666 4176 8722 4185
rect 8772 4146 8800 4422
rect 8864 4282 8892 10406
rect 8956 9654 8984 15642
rect 9048 15570 9076 15914
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9048 12986 9076 13466
rect 9140 13025 9168 19615
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9218 18592 9274 18601
rect 9218 18527 9274 18536
rect 9232 17542 9260 18527
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9232 14113 9260 16934
rect 9324 16250 9352 19246
rect 9416 16998 9444 19654
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9508 15910 9536 20198
rect 9588 18216 9640 18222
rect 9586 18184 9588 18193
rect 9640 18184 9642 18193
rect 9586 18119 9642 18128
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9600 16726 9628 17070
rect 9588 16720 9640 16726
rect 9588 16662 9640 16668
rect 9600 16250 9628 16662
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9496 15632 9548 15638
rect 9496 15574 9548 15580
rect 9508 15026 9536 15574
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9218 14104 9274 14113
rect 9218 14039 9274 14048
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9126 13016 9182 13025
rect 9036 12980 9088 12986
rect 9126 12951 9182 12960
rect 9036 12922 9088 12928
rect 9232 12832 9260 13942
rect 9416 13394 9444 14282
rect 9508 14278 9536 14962
rect 9586 14920 9642 14929
rect 9586 14855 9588 14864
rect 9640 14855 9642 14864
rect 9588 14826 9640 14832
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9324 13025 9352 13330
rect 9416 13138 9444 13330
rect 9508 13326 9536 14214
rect 9600 13938 9628 14486
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9416 13110 9536 13138
rect 9310 13016 9366 13025
rect 9310 12951 9366 12960
rect 9232 12804 9444 12832
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9218 12608 9274 12617
rect 9218 12543 9274 12552
rect 9126 12472 9182 12481
rect 9232 12442 9260 12543
rect 9126 12407 9182 12416
rect 9220 12436 9272 12442
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9048 11937 9076 12242
rect 9034 11928 9090 11937
rect 9034 11863 9090 11872
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9048 11354 9076 11698
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8956 9178 8984 9590
rect 9048 9518 9076 11290
rect 9140 10538 9168 12407
rect 9220 12378 9272 12384
rect 9324 12356 9352 12650
rect 9416 12481 9444 12804
rect 9508 12782 9536 13110
rect 9600 12918 9628 13738
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9402 12472 9458 12481
rect 9402 12407 9458 12416
rect 9324 12328 9444 12356
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9232 11082 9260 11834
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9232 10418 9260 11018
rect 9140 10390 9260 10418
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9140 9364 9168 10390
rect 9218 10296 9274 10305
rect 9218 10231 9274 10240
rect 9232 10062 9260 10231
rect 9324 10169 9352 10406
rect 9310 10160 9366 10169
rect 9310 10095 9366 10104
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9232 9489 9260 9862
rect 9218 9480 9274 9489
rect 9218 9415 9220 9424
rect 9272 9415 9274 9424
rect 9220 9386 9272 9392
rect 9048 9336 9168 9364
rect 9232 9355 9260 9386
rect 9324 9353 9352 9930
rect 9310 9344 9366 9353
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8956 8634 8984 8910
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8956 8090 8984 8230
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8942 6352 8998 6361
rect 8942 6287 8998 6296
rect 8956 6186 8984 6287
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8956 5545 8984 5782
rect 8942 5536 8998 5545
rect 8942 5471 8998 5480
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8956 4162 8984 5102
rect 8666 4111 8722 4120
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8864 4134 8984 4162
rect 8864 4026 8892 4134
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8404 3590 8524 3618
rect 8680 3998 8892 4026
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8576 3596 8628 3602
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 7748 3392 7800 3398
rect 7470 3360 7526 3369
rect 7748 3334 7800 3340
rect 7470 3295 7526 3304
rect 7484 2650 7512 3295
rect 7562 3088 7618 3097
rect 7562 3023 7618 3032
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7576 2582 7604 3023
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7668 2378 7696 2926
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 7760 1442 7788 3334
rect 8128 2922 8156 3470
rect 8220 3466 8248 3538
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8300 3188 8352 3194
rect 8404 3176 8432 3590
rect 8576 3538 8628 3544
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8496 3194 8524 3470
rect 8352 3148 8432 3176
rect 8484 3188 8536 3194
rect 8300 3130 8352 3136
rect 8484 3130 8536 3136
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8116 2916 8168 2922
rect 8116 2858 8168 2864
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8220 1442 8248 3062
rect 8588 2378 8616 3538
rect 8680 2961 8708 3998
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8772 3058 8800 3674
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8666 2952 8722 2961
rect 8666 2887 8722 2896
rect 8680 2650 8708 2887
rect 8772 2854 8800 2994
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8668 2508 8720 2514
rect 8668 2450 8720 2456
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 7668 1414 7788 1442
rect 8128 1414 8248 1442
rect 7668 800 7696 1414
rect 8128 800 8156 1414
rect 8496 800 8524 2246
rect 8680 1970 8708 2450
rect 8772 2446 8800 2790
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8668 1964 8720 1970
rect 8668 1906 8720 1912
rect 8864 1902 8892 2926
rect 8852 1896 8904 1902
rect 8852 1838 8904 1844
rect 8956 800 8984 4014
rect 9048 3738 9076 9336
rect 9310 9279 9366 9288
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9140 8430 9168 8774
rect 9218 8664 9274 8673
rect 9218 8599 9274 8608
rect 9232 8430 9260 8599
rect 9310 8528 9366 8537
rect 9416 8514 9444 12328
rect 9508 12073 9536 12718
rect 9600 12442 9628 12718
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9494 12064 9550 12073
rect 9494 11999 9550 12008
rect 9496 11552 9548 11558
rect 9494 11520 9496 11529
rect 9692 11529 9720 20266
rect 9784 19922 9812 20334
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9876 19310 9904 20538
rect 10152 20398 10180 22200
rect 10140 20392 10192 20398
rect 10046 20360 10102 20369
rect 10140 20334 10192 20340
rect 10046 20295 10102 20304
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 9784 17882 9812 18566
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9784 17241 9812 17614
rect 9876 17513 9904 17682
rect 9862 17504 9918 17513
rect 9862 17439 9918 17448
rect 9770 17232 9826 17241
rect 9770 17167 9826 17176
rect 9784 12481 9812 17167
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9876 16561 9904 16594
rect 9862 16552 9918 16561
rect 9862 16487 9918 16496
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9968 16130 9996 20198
rect 10060 19334 10088 20295
rect 10152 19786 10180 20334
rect 10520 19922 10548 22200
rect 10888 20534 10916 22200
rect 11256 20534 11284 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11716 20534 11744 22200
rect 12084 20534 12112 22200
rect 12452 20534 12480 22200
rect 12820 20534 12848 22200
rect 13188 20534 13216 22200
rect 13556 20534 13584 22200
rect 14016 20534 14044 22200
rect 10692 20528 10744 20534
rect 10692 20470 10744 20476
rect 10876 20528 10928 20534
rect 10876 20470 10928 20476
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 11704 20528 11756 20534
rect 11704 20470 11756 20476
rect 12072 20528 12124 20534
rect 12072 20470 12124 20476
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 13176 20528 13228 20534
rect 13176 20470 13228 20476
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 10704 20398 10732 20470
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10508 19916 10560 19922
rect 10508 19858 10560 19864
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10060 19306 10180 19334
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10060 17882 10088 18702
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 10060 16590 10088 17138
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9876 15910 9904 16118
rect 9968 16102 10088 16130
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9876 14074 9904 14758
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9864 13728 9916 13734
rect 9862 13696 9864 13705
rect 9916 13696 9918 13705
rect 9862 13631 9918 13640
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9770 12472 9826 12481
rect 9770 12407 9826 12416
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9784 11762 9812 12174
rect 9876 12170 9904 12922
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9548 11520 9550 11529
rect 9494 11455 9550 11464
rect 9678 11520 9734 11529
rect 9968 11506 9996 15982
rect 10060 12442 10088 16102
rect 10152 13841 10180 19306
rect 10244 16046 10272 19654
rect 10336 19514 10364 19858
rect 10704 19718 10732 20334
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11428 20324 11480 20330
rect 11428 20266 11480 20272
rect 12072 20324 12124 20330
rect 12072 20266 12124 20272
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 12808 20324 12860 20330
rect 12808 20266 12860 20272
rect 13176 20324 13228 20330
rect 13176 20266 13228 20272
rect 13544 20324 13596 20330
rect 13544 20266 13596 20272
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 14280 20324 14332 20330
rect 14280 20266 14332 20272
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10692 19712 10744 19718
rect 10692 19654 10744 19660
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10416 19168 10468 19174
rect 10416 19110 10468 19116
rect 10428 18970 10456 19110
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10612 18154 10640 19314
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10428 17882 10456 18022
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10336 16658 10364 17682
rect 10612 17678 10640 18090
rect 10796 17762 10824 20198
rect 11072 19310 11100 20266
rect 11440 20058 11468 20266
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11256 19514 11284 19858
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 10888 17882 10916 19110
rect 11072 18970 11100 19110
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10968 18896 11020 18902
rect 11020 18844 11100 18850
rect 10968 18838 11100 18844
rect 10980 18822 11100 18838
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 11072 18034 11100 18822
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11164 18358 11192 18770
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10796 17734 10916 17762
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10612 17202 10640 17614
rect 10784 17604 10836 17610
rect 10784 17546 10836 17552
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10416 16720 10468 16726
rect 10414 16688 10416 16697
rect 10468 16688 10470 16697
rect 10324 16652 10376 16658
rect 10414 16623 10470 16632
rect 10324 16594 10376 16600
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10138 13832 10194 13841
rect 10138 13767 10194 13776
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10152 13530 10180 13670
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10244 13258 10272 15506
rect 10336 14890 10364 16186
rect 10324 14884 10376 14890
rect 10324 14826 10376 14832
rect 10336 14793 10364 14826
rect 10322 14784 10378 14793
rect 10322 14719 10378 14728
rect 10428 14113 10456 16526
rect 10414 14104 10470 14113
rect 10414 14039 10470 14048
rect 10520 13841 10548 16730
rect 10612 14890 10640 16934
rect 10796 16794 10824 17546
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10888 16504 10916 17734
rect 10980 17134 11008 18022
rect 11072 18006 11192 18034
rect 11164 17678 11192 18006
rect 11152 17672 11204 17678
rect 11058 17640 11114 17649
rect 11152 17614 11204 17620
rect 11058 17575 11114 17584
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10980 16794 11008 16934
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10704 16476 10916 16504
rect 10704 14906 10732 16476
rect 10980 16436 11008 16730
rect 11072 16697 11100 17575
rect 11164 17270 11192 17614
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11058 16688 11114 16697
rect 11058 16623 11114 16632
rect 11152 16652 11204 16658
rect 11072 16590 11100 16623
rect 11152 16594 11204 16600
rect 11060 16584 11112 16590
rect 11164 16561 11192 16594
rect 11060 16526 11112 16532
rect 11150 16552 11206 16561
rect 11150 16487 11206 16496
rect 10888 16408 11008 16436
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10796 15502 10824 15914
rect 10888 15586 10916 16408
rect 11256 15706 11284 19246
rect 11808 19242 11836 19654
rect 12084 19446 12112 20266
rect 12452 19514 12480 20266
rect 12820 20058 12848 20266
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11796 19236 11848 19242
rect 11796 19178 11848 19184
rect 11808 18766 11836 19178
rect 11900 18970 11928 19314
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11336 17672 11388 17678
rect 11334 17640 11336 17649
rect 11388 17640 11390 17649
rect 11334 17575 11390 17584
rect 11624 17524 11652 18158
rect 11716 17678 11744 18294
rect 11900 18154 11928 18906
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 11992 17882 12020 18770
rect 12084 17882 12112 19110
rect 12268 18834 12296 19246
rect 12544 19174 12572 19858
rect 13188 19514 13216 20266
rect 13556 19514 13584 20266
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13648 19310 13676 19654
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12820 18970 12848 19246
rect 12900 19236 12952 19242
rect 12900 19178 12952 19184
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11624 17496 11744 17524
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11716 17134 11744 17496
rect 11992 17338 12020 17682
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11612 17060 11664 17066
rect 11612 17002 11664 17008
rect 11624 16794 11652 17002
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11716 15910 11744 16662
rect 11808 16114 11836 17138
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 10888 15558 11008 15586
rect 11164 15570 11192 15642
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10888 15162 10916 15438
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10600 14884 10652 14890
rect 10704 14878 10916 14906
rect 10600 14826 10652 14832
rect 10506 13832 10562 13841
rect 10324 13796 10376 13802
rect 10506 13767 10562 13776
rect 10324 13738 10376 13744
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10230 12880 10286 12889
rect 10140 12844 10192 12850
rect 10230 12815 10286 12824
rect 10140 12786 10192 12792
rect 10152 12617 10180 12786
rect 10138 12608 10194 12617
rect 10138 12543 10194 12552
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10060 12238 10088 12378
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10152 11762 10180 12378
rect 10244 12238 10272 12815
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9678 11455 9734 11464
rect 9784 11478 9996 11506
rect 10046 11520 10102 11529
rect 9784 11336 9812 11478
rect 10046 11455 10102 11464
rect 9692 11308 9812 11336
rect 9862 11384 9918 11393
rect 10060 11370 10088 11455
rect 9862 11319 9918 11328
rect 9968 11342 10088 11370
rect 9692 10742 9720 11308
rect 9876 11150 9904 11319
rect 9968 11286 9996 11342
rect 9956 11280 10008 11286
rect 10152 11234 10180 11698
rect 9956 11222 10008 11228
rect 10060 11206 10180 11234
rect 10060 11150 10088 11206
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9770 10976 9826 10985
rect 9770 10911 9826 10920
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9784 10674 9812 10911
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9508 10441 9536 10610
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9494 10432 9550 10441
rect 9494 10367 9550 10376
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9494 9208 9550 9217
rect 9494 9143 9550 9152
rect 9508 9042 9536 9143
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9600 8922 9628 10202
rect 9692 9217 9720 10542
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9678 9208 9734 9217
rect 9678 9143 9734 9152
rect 9784 8974 9812 10066
rect 9366 8486 9444 8514
rect 9508 8894 9628 8922
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9310 8463 9366 8472
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9324 8294 9352 8463
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9402 8256 9458 8265
rect 9402 8191 9458 8200
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 9310 7984 9366 7993
rect 9232 7478 9260 7958
rect 9310 7919 9366 7928
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 9324 7410 9352 7919
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9126 7168 9182 7177
rect 9126 7103 9182 7112
rect 9140 6497 9168 7103
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9126 6488 9182 6497
rect 9126 6423 9182 6432
rect 9126 6352 9182 6361
rect 9126 6287 9182 6296
rect 9140 6118 9168 6287
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9232 5166 9260 6938
rect 9312 6792 9364 6798
rect 9416 6780 9444 8191
rect 9364 6752 9444 6780
rect 9312 6734 9364 6740
rect 9404 6656 9456 6662
rect 9402 6624 9404 6633
rect 9456 6624 9458 6633
rect 9402 6559 9458 6568
rect 9508 6458 9536 8894
rect 9784 8838 9812 8910
rect 9772 8832 9824 8838
rect 9586 8800 9642 8809
rect 9642 8758 9720 8786
rect 9772 8774 9824 8780
rect 9586 8735 9642 8744
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9600 8022 9628 8366
rect 9588 8016 9640 8022
rect 9692 7993 9720 8758
rect 9588 7958 9640 7964
rect 9678 7984 9734 7993
rect 9678 7919 9734 7928
rect 9692 7188 9720 7919
rect 9784 7750 9812 8774
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9692 7160 9812 7188
rect 9784 6914 9812 7160
rect 9692 6886 9812 6914
rect 9692 6798 9720 6886
rect 9876 6866 9904 11086
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 9518 9996 10542
rect 10152 10520 10180 11086
rect 10060 10492 10180 10520
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9968 8090 9996 9454
rect 10060 8673 10088 10492
rect 10138 10432 10194 10441
rect 10138 10367 10194 10376
rect 10152 9178 10180 10367
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10140 8832 10192 8838
rect 10138 8800 10140 8809
rect 10192 8800 10194 8809
rect 10138 8735 10194 8744
rect 10046 8664 10102 8673
rect 10046 8599 10102 8608
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10152 8401 10180 8570
rect 10138 8392 10194 8401
rect 10048 8356 10100 8362
rect 10138 8327 10194 8336
rect 10048 8298 10100 8304
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9968 7313 9996 7414
rect 9954 7304 10010 7313
rect 9954 7239 10010 7248
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9680 6792 9732 6798
rect 9876 6769 9904 6802
rect 9680 6734 9732 6740
rect 9862 6760 9918 6769
rect 9862 6695 9918 6704
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9692 6497 9720 6598
rect 9678 6488 9734 6497
rect 9496 6452 9548 6458
rect 9678 6423 9734 6432
rect 9496 6394 9548 6400
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 9140 4690 9168 5034
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9232 4758 9260 4966
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9324 4570 9352 6122
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9232 4542 9352 4570
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9232 3670 9260 4542
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 4282 9352 4422
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9416 4010 9444 6054
rect 9508 5574 9536 6394
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9692 6089 9720 6326
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9678 6080 9734 6089
rect 9678 6015 9734 6024
rect 9784 5642 9812 6258
rect 9968 6254 9996 6598
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9678 5536 9734 5545
rect 9678 5471 9734 5480
rect 9692 4826 9720 5471
rect 9784 5166 9812 5578
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9876 4826 9904 6054
rect 9954 5944 10010 5953
rect 9954 5879 10010 5888
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9772 4616 9824 4622
rect 9824 4576 9904 4604
rect 9968 4593 9996 5879
rect 9772 4558 9824 4564
rect 9508 4214 9536 4558
rect 9876 4214 9904 4576
rect 9954 4584 10010 4593
rect 9954 4519 10010 4528
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9232 3398 9260 3606
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9416 3126 9444 3946
rect 9692 3398 9720 4082
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9784 3738 9812 3878
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9692 2990 9720 3334
rect 9770 3224 9826 3233
rect 9770 3159 9772 3168
rect 9824 3159 9826 3168
rect 9772 3130 9824 3136
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9772 2848 9824 2854
rect 9678 2816 9734 2825
rect 9772 2790 9824 2796
rect 9678 2751 9734 2760
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9048 2310 9076 2586
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9416 800 9444 2314
rect 9600 2281 9628 2518
rect 9692 2446 9720 2751
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9586 2272 9642 2281
rect 9586 2207 9642 2216
rect 9600 1630 9628 2207
rect 9692 1698 9720 2382
rect 9680 1692 9732 1698
rect 9680 1634 9732 1640
rect 9588 1624 9640 1630
rect 9588 1566 9640 1572
rect 9784 800 9812 2790
rect 9876 1970 9904 4150
rect 10060 3942 10088 8298
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3670 10088 3878
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 10046 3496 10102 3505
rect 10046 3431 10102 3440
rect 10060 2650 10088 3431
rect 10152 2922 10180 8230
rect 10244 7546 10272 12174
rect 10336 9178 10364 13738
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10428 12238 10456 13670
rect 10520 12889 10548 13767
rect 10612 13682 10640 14826
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14532 10824 14758
rect 10796 14504 10833 14532
rect 10692 14408 10744 14414
rect 10805 14362 10833 14504
rect 10692 14350 10744 14356
rect 10704 14278 10732 14350
rect 10796 14346 10833 14362
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10704 14006 10732 14214
rect 10782 14104 10838 14113
rect 10782 14039 10838 14048
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10612 13654 10732 13682
rect 10598 13560 10654 13569
rect 10598 13495 10654 13504
rect 10506 12880 10562 12889
rect 10506 12815 10562 12824
rect 10508 12776 10560 12782
rect 10612 12764 10640 13495
rect 10704 12986 10732 13654
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10560 12736 10640 12764
rect 10508 12718 10560 12724
rect 10520 12374 10548 12718
rect 10508 12368 10560 12374
rect 10508 12310 10560 12316
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10414 12064 10470 12073
rect 10414 11999 10470 12008
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10428 9110 10456 11999
rect 10520 11694 10548 12310
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10508 11688 10560 11694
rect 10612 11665 10640 11834
rect 10508 11630 10560 11636
rect 10598 11656 10654 11665
rect 10598 11591 10654 11600
rect 10692 11552 10744 11558
rect 10598 11520 10654 11529
rect 10692 11494 10744 11500
rect 10598 11455 10654 11464
rect 10506 11384 10562 11393
rect 10612 11354 10640 11455
rect 10506 11319 10562 11328
rect 10600 11348 10652 11354
rect 10520 11218 10548 11319
rect 10600 11290 10652 11296
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10704 11150 10732 11494
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10690 10976 10746 10985
rect 10690 10911 10746 10920
rect 10598 10840 10654 10849
rect 10598 10775 10654 10784
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10520 9722 10548 10474
rect 10612 10441 10640 10775
rect 10598 10432 10654 10441
rect 10598 10367 10654 10376
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10416 9104 10468 9110
rect 10336 9052 10416 9058
rect 10336 9046 10468 9052
rect 10336 9030 10456 9046
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10336 7426 10364 9030
rect 10520 8974 10548 9658
rect 10612 9518 10640 9998
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10428 8650 10456 8910
rect 10428 8622 10548 8650
rect 10612 8634 10640 8978
rect 10520 8566 10548 8622
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10428 8022 10456 8434
rect 10704 8344 10732 10911
rect 10612 8316 10732 8344
rect 10612 8022 10640 8316
rect 10796 8242 10824 14039
rect 10888 13569 10916 14878
rect 10980 14385 11008 15558
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11072 14550 11100 14962
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 11164 14618 11192 14826
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 10966 14376 11022 14385
rect 10966 14311 11022 14320
rect 10874 13560 10930 13569
rect 10874 13495 10930 13504
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10888 12850 10916 13330
rect 10980 12889 11008 14311
rect 11060 14272 11112 14278
rect 11348 14260 11376 14894
rect 11426 14512 11482 14521
rect 11426 14447 11428 14456
rect 11480 14447 11482 14456
rect 11428 14418 11480 14424
rect 11060 14214 11112 14220
rect 11256 14232 11376 14260
rect 11072 13462 11100 14214
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11058 13016 11114 13025
rect 11058 12951 11114 12960
rect 10966 12880 11022 12889
rect 10876 12844 10928 12850
rect 10966 12815 11022 12824
rect 10876 12786 10928 12792
rect 10888 12442 10916 12786
rect 10968 12640 11020 12646
rect 10966 12608 10968 12617
rect 11020 12608 11022 12617
rect 10966 12543 11022 12552
rect 10966 12472 11022 12481
rect 10876 12436 10928 12442
rect 10966 12407 11022 12416
rect 10876 12378 10928 12384
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10888 11354 10916 12242
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10980 10588 11008 12407
rect 11072 11626 11100 12951
rect 11256 12850 11284 14232
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11348 13705 11376 13806
rect 11334 13696 11390 13705
rect 11334 13631 11390 13640
rect 11426 13560 11482 13569
rect 11426 13495 11482 13504
rect 11440 13297 11468 13495
rect 11426 13288 11482 13297
rect 11426 13223 11482 13232
rect 11716 13190 11744 15846
rect 11808 14958 11836 16050
rect 11900 15706 11928 17002
rect 12268 16250 12296 18770
rect 12820 18698 12848 18906
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12912 18630 12940 19178
rect 13728 19168 13780 19174
rect 13832 19156 13860 20266
rect 14292 19514 14320 20266
rect 14384 19990 14412 22200
rect 14752 20534 14780 22200
rect 15120 20534 15148 22200
rect 15488 20534 15516 22200
rect 15856 20534 15884 22200
rect 16316 20534 16344 22200
rect 16684 20534 16712 22200
rect 17052 20534 17080 22200
rect 17420 20534 17448 22200
rect 17498 22199 17554 22208
rect 17774 22200 17830 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 18970 22200 19026 23000
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 19890 22672 19946 22681
rect 19890 22607 19946 22616
rect 14740 20528 14792 20534
rect 14740 20470 14792 20476
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 15476 20528 15528 20534
rect 15476 20470 15528 20476
rect 15844 20528 15896 20534
rect 15844 20470 15896 20476
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16672 20528 16724 20534
rect 16672 20470 16724 20476
rect 17040 20528 17092 20534
rect 17040 20470 17092 20476
rect 17408 20528 17460 20534
rect 17408 20470 17460 20476
rect 14648 20324 14700 20330
rect 14648 20266 14700 20272
rect 15200 20324 15252 20330
rect 15200 20266 15252 20272
rect 15660 20324 15712 20330
rect 15660 20266 15712 20272
rect 16028 20324 16080 20330
rect 16028 20266 16080 20272
rect 16488 20324 16540 20330
rect 16488 20266 16540 20272
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 17408 20324 17460 20330
rect 17408 20266 17460 20272
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14004 19304 14056 19310
rect 14464 19304 14516 19310
rect 14004 19246 14056 19252
rect 14384 19252 14464 19258
rect 14384 19246 14516 19252
rect 13780 19128 13860 19156
rect 13728 19110 13780 19116
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12360 17270 12388 17546
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12360 16130 12388 17206
rect 12452 17202 12480 18158
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12544 16658 12572 18022
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12268 16102 12388 16130
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11900 15366 11928 15642
rect 11980 15496 12032 15502
rect 11978 15464 11980 15473
rect 12032 15464 12034 15473
rect 11978 15399 12034 15408
rect 11888 15360 11940 15366
rect 11886 15328 11888 15337
rect 11980 15360 12032 15366
rect 11940 15328 11942 15337
rect 11980 15302 12032 15308
rect 11886 15263 11942 15272
rect 11992 15201 12020 15302
rect 11978 15192 12034 15201
rect 11978 15127 12034 15136
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11808 14498 11836 14894
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 12176 14793 12204 14826
rect 12162 14784 12218 14793
rect 12162 14719 12218 14728
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 11808 14470 11928 14498
rect 11900 14278 11928 14470
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11808 13530 11836 14214
rect 11992 14006 12020 14418
rect 12176 14414 12204 14554
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 11980 14000 12032 14006
rect 12032 13960 12112 13988
rect 11980 13942 12032 13948
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11900 13530 11928 13874
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11610 12472 11666 12481
rect 11610 12407 11666 12416
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11348 12084 11376 12310
rect 11150 12064 11206 12073
rect 11150 11999 11206 12008
rect 11256 12056 11376 12084
rect 11624 12084 11652 12407
rect 11716 12306 11744 12786
rect 11900 12714 11928 13466
rect 11992 12986 12020 13670
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11900 12594 11928 12650
rect 11900 12566 12020 12594
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11624 12056 11744 12084
rect 11164 11762 11192 11999
rect 11256 11762 11284 12056
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11716 11812 11744 12056
rect 11624 11784 11744 11812
rect 11808 11801 11836 12378
rect 11992 12238 12020 12566
rect 12084 12442 12112 13960
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12176 13530 12204 13670
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 12268 13410 12296 16102
rect 12452 16046 12480 16526
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12440 15496 12492 15502
rect 12544 15484 12572 16594
rect 12728 15706 12756 16594
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12912 15502 12940 18566
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13096 16658 13124 17614
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13464 17338 13492 17546
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13464 17202 13492 17274
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13268 17060 13320 17066
rect 13268 17002 13320 17008
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 13280 16590 13308 17002
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13280 16250 13308 16526
rect 13556 16250 13584 17682
rect 13832 17066 13860 18362
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13832 16833 13860 17002
rect 13818 16824 13874 16833
rect 13818 16759 13874 16768
rect 13924 16658 13952 17070
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13740 16046 13768 16390
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13188 15502 13216 15982
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 12492 15456 12572 15484
rect 12900 15496 12952 15502
rect 12440 15438 12492 15444
rect 12900 15438 12952 15444
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 12346 15192 12402 15201
rect 12346 15127 12348 15136
rect 12400 15127 12402 15136
rect 12348 15098 12400 15104
rect 12452 14958 12480 15438
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12360 14385 12388 14758
rect 12452 14414 12480 14894
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12440 14408 12492 14414
rect 12346 14376 12402 14385
rect 12440 14350 12492 14356
rect 12346 14311 12402 14320
rect 12360 13530 12388 14311
rect 12544 14074 12572 14554
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12636 13716 12664 14486
rect 13004 14414 13032 14894
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12820 14113 12848 14350
rect 12806 14104 12862 14113
rect 12806 14039 12862 14048
rect 13096 13802 13124 15030
rect 13188 15026 13216 15438
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13188 14822 13216 14962
rect 13280 14822 13308 15506
rect 13464 15473 13492 15506
rect 13450 15464 13506 15473
rect 13450 15399 13506 15408
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13372 14074 13400 14214
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13464 13938 13492 14214
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13556 13870 13584 14962
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13648 14006 13676 14486
rect 13740 14249 13768 15982
rect 13832 15162 13860 16594
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15706 13952 15846
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13726 14240 13782 14249
rect 13726 14175 13782 14184
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13084 13796 13136 13802
rect 13084 13738 13136 13744
rect 12544 13688 12664 13716
rect 12808 13728 12860 13734
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12268 13382 12480 13410
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11794 11792 11850 11801
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11072 10742 11100 11562
rect 11164 11558 11192 11698
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 10980 10560 11100 10588
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 11072 10418 11100 10560
rect 11164 10538 11192 11494
rect 11256 11150 11284 11698
rect 11624 11150 11652 11784
rect 11794 11727 11850 11736
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11256 10810 11284 11086
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 10980 10266 11008 10406
rect 11072 10390 11192 10418
rect 11058 10296 11114 10305
rect 10968 10260 11020 10266
rect 11058 10231 11114 10240
rect 10968 10202 11020 10208
rect 10968 10056 11020 10062
rect 10888 10016 10968 10044
rect 10888 8634 10916 10016
rect 10968 9998 11020 10004
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 9518 11008 9862
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10980 9178 11008 9318
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 11072 8809 11100 10231
rect 11164 9466 11192 10390
rect 11624 10282 11652 10610
rect 11624 10254 11744 10282
rect 11808 10266 11836 11727
rect 11992 11626 12020 12038
rect 12084 11898 12112 12174
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 11980 11620 12032 11626
rect 11980 11562 12032 11568
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11256 9654 11284 9930
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11716 9704 11744 10254
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11532 9676 11744 9704
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11164 9438 11284 9466
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11164 9178 11192 9318
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11058 8800 11114 8809
rect 11058 8735 11114 8744
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10888 8265 10916 8298
rect 10704 8214 10824 8242
rect 10874 8256 10930 8265
rect 10416 8016 10468 8022
rect 10600 8016 10652 8022
rect 10416 7958 10468 7964
rect 10520 7976 10600 8004
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10428 7721 10456 7822
rect 10414 7712 10470 7721
rect 10414 7647 10470 7656
rect 10244 7398 10364 7426
rect 10244 5012 10272 7398
rect 10416 7268 10468 7274
rect 10416 7210 10468 7216
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10336 7002 10364 7142
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10322 6896 10378 6905
rect 10322 6831 10324 6840
rect 10376 6831 10378 6840
rect 10324 6802 10376 6808
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10336 5846 10364 6598
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10428 5522 10456 7210
rect 10520 6905 10548 7976
rect 10600 7958 10652 7964
rect 10600 7744 10652 7750
rect 10598 7712 10600 7721
rect 10652 7712 10654 7721
rect 10598 7647 10654 7656
rect 10598 7576 10654 7585
rect 10598 7511 10654 7520
rect 10612 7313 10640 7511
rect 10598 7304 10654 7313
rect 10598 7239 10654 7248
rect 10600 7200 10652 7206
rect 10598 7168 10600 7177
rect 10652 7168 10654 7177
rect 10598 7103 10654 7112
rect 10506 6896 10562 6905
rect 10506 6831 10562 6840
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10520 5778 10548 6734
rect 10704 6662 10732 8214
rect 10874 8191 10930 8200
rect 10980 8090 11008 8434
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10612 5953 10640 6054
rect 10598 5944 10654 5953
rect 10598 5879 10654 5888
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10336 5494 10456 5522
rect 10336 5137 10364 5494
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10322 5128 10378 5137
rect 10322 5063 10378 5072
rect 10244 4984 10364 5012
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10244 3040 10272 3946
rect 10336 3738 10364 4984
rect 10428 3942 10456 5306
rect 10520 4758 10548 5714
rect 10796 5710 10824 8026
rect 10980 7274 11008 8026
rect 11072 7324 11100 8570
rect 11164 7721 11192 8978
rect 11256 8634 11284 9438
rect 11532 9178 11560 9676
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11702 9480 11758 9489
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11532 9042 11560 9114
rect 11624 9110 11652 9454
rect 11702 9415 11758 9424
rect 11716 9382 11744 9415
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11900 9042 11928 11086
rect 11992 10849 12020 11154
rect 12176 11082 12204 12242
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12162 10976 12218 10985
rect 12162 10911 12218 10920
rect 11978 10840 12034 10849
rect 11978 10775 11980 10784
rect 12032 10775 12034 10784
rect 11980 10746 12032 10752
rect 11992 10715 12020 10746
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11992 9110 12020 9522
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11150 7712 11206 7721
rect 11150 7647 11206 7656
rect 11256 7478 11284 8434
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11072 7296 11192 7324
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 11164 7206 11192 7296
rect 11426 7304 11482 7313
rect 11426 7239 11482 7248
rect 11440 7206 11468 7239
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 10874 7032 10930 7041
rect 10874 6967 10930 6976
rect 10784 5704 10836 5710
rect 10704 5652 10784 5658
rect 10704 5646 10836 5652
rect 10704 5630 10824 5646
rect 10704 5166 10732 5630
rect 10782 5536 10838 5545
rect 10782 5471 10838 5480
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10244 3012 10364 3040
rect 10336 2961 10364 3012
rect 10322 2952 10378 2961
rect 10140 2916 10192 2922
rect 10140 2858 10192 2864
rect 10232 2916 10284 2922
rect 10322 2887 10378 2896
rect 10232 2858 10284 2864
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9864 1964 9916 1970
rect 9864 1906 9916 1912
rect 10152 1834 10180 2858
rect 10140 1828 10192 1834
rect 10140 1770 10192 1776
rect 10244 800 10272 2858
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10520 2553 10548 2586
rect 10506 2544 10562 2553
rect 10506 2479 10562 2488
rect 10520 2038 10548 2479
rect 10508 2032 10560 2038
rect 10508 1974 10560 1980
rect 10612 800 10640 4014
rect 10704 3398 10732 5102
rect 10796 4622 10824 5471
rect 10888 5012 10916 6967
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 6769 11008 6802
rect 10966 6760 11022 6769
rect 10966 6695 11022 6704
rect 11072 6474 11100 7142
rect 11164 7041 11192 7142
rect 11440 7041 11468 7142
rect 11150 7032 11206 7041
rect 11150 6967 11206 6976
rect 11426 7032 11482 7041
rect 11426 6967 11482 6976
rect 11152 6928 11204 6934
rect 11532 6916 11560 7142
rect 11204 6888 11560 6916
rect 11152 6870 11204 6876
rect 11152 6792 11204 6798
rect 11204 6752 11836 6780
rect 11152 6734 11204 6740
rect 11808 6662 11836 6752
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 10980 6458 11100 6474
rect 10968 6452 11100 6458
rect 11020 6446 11100 6452
rect 11150 6488 11206 6497
rect 11352 6480 11648 6500
rect 11206 6458 11284 6474
rect 11206 6452 11296 6458
rect 11206 6446 11244 6452
rect 11150 6423 11206 6432
rect 10968 6394 11020 6400
rect 11244 6394 11296 6400
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11426 6352 11482 6361
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10980 5914 11008 6054
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 11072 5166 11100 6326
rect 11336 6316 11388 6322
rect 11426 6287 11482 6296
rect 11336 6258 11388 6264
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11164 5234 11192 6054
rect 11256 5846 11284 6122
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11244 5636 11296 5642
rect 11348 5624 11376 6258
rect 11440 6118 11468 6287
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11610 6216 11666 6225
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11532 5953 11560 6190
rect 11610 6151 11666 6160
rect 11624 6118 11652 6151
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11518 5944 11574 5953
rect 11518 5879 11574 5888
rect 11624 5778 11652 6054
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11296 5596 11376 5624
rect 11244 5578 11296 5584
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11612 5024 11664 5030
rect 10888 4984 11192 5012
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10704 2990 10732 3334
rect 10796 3126 10824 3606
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 10692 2984 10744 2990
rect 10692 2926 10744 2932
rect 10888 2854 10916 4082
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10980 2990 11008 3946
rect 11072 3505 11100 4558
rect 11164 3641 11192 4984
rect 11612 4966 11664 4972
rect 11624 4758 11652 4966
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11150 3632 11206 3641
rect 11150 3567 11206 3576
rect 11058 3496 11114 3505
rect 11058 3431 11114 3440
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 11072 2446 11100 3334
rect 11164 3194 11192 3567
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11164 1442 11192 2858
rect 11256 1630 11284 4558
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11716 4078 11744 6598
rect 11808 5846 11836 6598
rect 11900 6202 11928 8842
rect 11900 6174 12020 6202
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11900 5953 11928 6054
rect 11886 5944 11942 5953
rect 11886 5879 11942 5888
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11808 4570 11836 5578
rect 11900 5166 11928 5714
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4690 11928 4966
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11808 4542 11928 4570
rect 11794 4448 11850 4457
rect 11794 4383 11850 4392
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11716 3194 11744 3538
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11334 3088 11390 3097
rect 11334 3023 11390 3032
rect 11348 2854 11376 3023
rect 11716 2854 11744 3130
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11808 2106 11836 4383
rect 11900 3097 11928 4542
rect 11992 3738 12020 6174
rect 12084 5642 12112 10610
rect 12176 10198 12204 10911
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12162 9888 12218 9897
rect 12162 9823 12218 9832
rect 12176 9722 12204 9823
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12176 8809 12204 8978
rect 12162 8800 12218 8809
rect 12162 8735 12218 8744
rect 12268 8616 12296 13126
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11801 12388 12038
rect 12346 11792 12402 11801
rect 12346 11727 12402 11736
rect 12452 11218 12480 13382
rect 12544 12322 12572 13688
rect 12808 13670 12860 13676
rect 12992 13728 13044 13734
rect 13648 13682 13676 13942
rect 12992 13670 13044 13676
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12636 12442 12664 13126
rect 12728 12850 12756 13330
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12716 12368 12768 12374
rect 12544 12294 12664 12322
rect 12716 12310 12768 12316
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 11830 12572 12038
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12636 10985 12664 12294
rect 12728 11762 12756 12310
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12820 11558 12848 13670
rect 13004 13530 13032 13670
rect 13556 13654 13676 13682
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 13556 13462 13584 13654
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13280 12646 13308 13194
rect 13358 12880 13414 12889
rect 13648 12850 13676 13466
rect 13358 12815 13414 12824
rect 13636 12844 13688 12850
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12912 11218 12940 12378
rect 13096 12374 13124 12582
rect 13372 12442 13400 12815
rect 13636 12786 13688 12792
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13450 12472 13506 12481
rect 13360 12436 13412 12442
rect 13450 12407 13452 12416
rect 13360 12378 13412 12384
rect 13504 12407 13506 12416
rect 13452 12378 13504 12384
rect 13648 12374 13676 12582
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13174 11656 13230 11665
rect 13174 11591 13230 11600
rect 13188 11286 13216 11591
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12622 10976 12678 10985
rect 12622 10911 12678 10920
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12176 8588 12296 8616
rect 12176 8430 12204 8588
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 8090 12204 8230
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12268 7954 12296 8434
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 12268 7721 12296 7890
rect 12254 7712 12310 7721
rect 12254 7647 12310 7656
rect 12360 7041 12388 10474
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12544 9897 12572 10134
rect 12728 9926 12756 10542
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12716 9920 12768 9926
rect 12530 9888 12586 9897
rect 12716 9862 12768 9868
rect 12530 9823 12586 9832
rect 12438 9752 12494 9761
rect 12438 9687 12440 9696
rect 12492 9687 12494 9696
rect 12440 9658 12492 9664
rect 12622 9616 12678 9625
rect 12622 9551 12678 9560
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12544 9178 12572 9386
rect 12636 9217 12664 9551
rect 12714 9480 12770 9489
rect 12820 9450 12848 10406
rect 12714 9415 12770 9424
rect 12808 9444 12860 9450
rect 12622 9208 12678 9217
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12532 9172 12584 9178
rect 12622 9143 12678 9152
rect 12532 9114 12584 9120
rect 12452 8922 12480 9114
rect 12530 8936 12586 8945
rect 12452 8894 12530 8922
rect 12530 8871 12586 8880
rect 12728 8838 12756 9415
rect 12808 9386 12860 9392
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12452 7818 12480 8298
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12346 7032 12402 7041
rect 12256 6996 12308 7002
rect 12452 7002 12480 7278
rect 12544 7188 12572 8570
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12636 7857 12664 7958
rect 12622 7848 12678 7857
rect 12622 7783 12678 7792
rect 12544 7160 12664 7188
rect 12346 6967 12402 6976
rect 12440 6996 12492 7002
rect 12256 6938 12308 6944
rect 12440 6938 12492 6944
rect 12162 6760 12218 6769
rect 12162 6695 12218 6704
rect 12176 5681 12204 6695
rect 12268 6458 12296 6938
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 12438 6896 12494 6905
rect 12360 6458 12388 6870
rect 12438 6831 12494 6840
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12162 5672 12218 5681
rect 12072 5636 12124 5642
rect 12162 5607 12218 5616
rect 12072 5578 12124 5584
rect 12268 5574 12296 6258
rect 12346 5944 12402 5953
rect 12452 5914 12480 6831
rect 12530 6624 12586 6633
rect 12530 6559 12586 6568
rect 12346 5879 12348 5888
rect 12400 5879 12402 5888
rect 12440 5908 12492 5914
rect 12348 5850 12400 5856
rect 12440 5850 12492 5856
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 12256 5228 12308 5234
rect 12176 5188 12256 5216
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11886 3088 11942 3097
rect 11886 3023 11942 3032
rect 12084 2378 12112 4626
rect 12176 4622 12204 5188
rect 12256 5170 12308 5176
rect 12360 5030 12388 5714
rect 12544 5642 12572 6559
rect 12636 6186 12664 7160
rect 12728 6322 12756 8502
rect 12820 8362 12848 8978
rect 12912 8362 12940 11154
rect 13280 11098 13308 12310
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13556 11354 13584 11494
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13544 11144 13596 11150
rect 13358 11112 13414 11121
rect 13280 11070 13358 11098
rect 13648 11132 13676 11494
rect 13740 11286 13768 14175
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13596 11104 13676 11132
rect 13544 11086 13596 11092
rect 13358 11047 13414 11056
rect 13452 11076 13504 11082
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13280 10606 13308 10746
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13174 10432 13230 10441
rect 13372 10418 13400 11047
rect 13452 11018 13504 11024
rect 13464 10606 13492 11018
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13372 10390 13492 10418
rect 13174 10367 13230 10376
rect 13188 9722 13216 10367
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 12990 9616 13046 9625
rect 12990 9551 13046 9560
rect 13176 9580 13228 9586
rect 13004 9518 13032 9551
rect 13176 9522 13228 9528
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13084 9376 13136 9382
rect 12990 9344 13046 9353
rect 13084 9318 13136 9324
rect 12990 9279 13046 9288
rect 13004 9178 13032 9279
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12820 7886 12848 8298
rect 13004 8242 13032 9114
rect 13096 8906 13124 9318
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 12912 8214 13032 8242
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 6662 12848 7822
rect 12912 7410 12940 8214
rect 12990 8120 13046 8129
rect 12990 8055 13046 8064
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6866 12940 7142
rect 13004 6934 13032 8055
rect 13096 7886 13124 8842
rect 13188 7954 13216 9522
rect 13280 9178 13308 10066
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13372 9042 13400 9318
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13266 8800 13322 8809
rect 13266 8735 13322 8744
rect 13280 8634 13308 8735
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13372 8090 13400 8230
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13084 7744 13136 7750
rect 13082 7712 13084 7721
rect 13136 7712 13138 7721
rect 13082 7647 13138 7656
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12912 6390 12940 6802
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12820 5817 12848 6122
rect 12900 5840 12952 5846
rect 12806 5808 12862 5817
rect 12900 5782 12952 5788
rect 12806 5743 12862 5752
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12820 5234 12848 5510
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12176 4146 12204 4558
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12164 3936 12216 3942
rect 12162 3904 12164 3913
rect 12216 3904 12218 3913
rect 12162 3839 12218 3848
rect 12268 3618 12296 4626
rect 12348 4480 12400 4486
rect 12346 4448 12348 4457
rect 12400 4448 12402 4457
rect 12346 4383 12402 4392
rect 12452 4162 12480 4626
rect 12544 4214 12572 5034
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12176 3590 12296 3618
rect 12360 4134 12480 4162
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12636 4146 12664 4490
rect 12624 4140 12676 4146
rect 12176 2650 12204 3590
rect 12360 2972 12388 4134
rect 12624 4082 12676 4088
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12438 3768 12494 3777
rect 12544 3738 12572 3946
rect 12438 3703 12494 3712
rect 12532 3732 12584 3738
rect 12452 3670 12480 3703
rect 12532 3674 12584 3680
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12636 3534 12664 4082
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12728 3738 12756 3878
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12820 3346 12848 3878
rect 12912 3670 12940 5782
rect 13096 5234 13124 7346
rect 13188 7002 13216 7890
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13188 6798 13216 6938
rect 13176 6792 13228 6798
rect 13280 6769 13308 7890
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13372 7585 13400 7686
rect 13358 7576 13414 7585
rect 13358 7511 13414 7520
rect 13372 7478 13400 7511
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 7002 13400 7142
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13176 6734 13228 6740
rect 13266 6760 13322 6769
rect 13188 6610 13216 6734
rect 13266 6695 13322 6704
rect 13188 6582 13308 6610
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13188 6225 13216 6394
rect 13174 6216 13230 6225
rect 13174 6151 13230 6160
rect 13280 5778 13308 6582
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13464 6202 13492 10390
rect 13556 10130 13584 11086
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13544 10124 13596 10130
rect 13648 10112 13676 10678
rect 13740 10470 13768 11222
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13728 10124 13780 10130
rect 13648 10084 13728 10112
rect 13544 10066 13596 10072
rect 13728 10066 13780 10072
rect 13556 8974 13584 10066
rect 13740 9586 13768 10066
rect 13832 10010 13860 13806
rect 13924 13734 13952 14758
rect 14016 14618 14044 19246
rect 14384 19230 14504 19246
rect 14384 17762 14412 19230
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18850 14504 19110
rect 14568 18970 14596 19858
rect 14660 19514 14688 20266
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 15212 19174 15240 20266
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14476 18822 14596 18850
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14476 17882 14504 18158
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14384 17734 14504 17762
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 15994 14320 16526
rect 14200 15966 14320 15994
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14108 15162 14136 15506
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14200 14906 14228 15966
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14292 15434 14320 15846
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 14096 14884 14148 14890
rect 14200 14878 14320 14906
rect 14096 14826 14148 14832
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 14016 12986 14044 14554
rect 14108 13161 14136 14826
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14094 13152 14150 13161
rect 14094 13087 14150 13096
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14016 12646 14044 12922
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13924 11014 13952 12582
rect 14200 12434 14228 14758
rect 14108 12406 14228 12434
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13924 10130 13952 10542
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 14016 10062 14044 12310
rect 14108 10606 14136 12406
rect 14292 12186 14320 14878
rect 14384 14822 14412 15642
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14384 13870 14412 14758
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14200 12158 14320 12186
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14108 10266 14136 10406
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14004 10056 14056 10062
rect 13832 9982 13952 10010
rect 14004 9998 14056 10004
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 9178 13768 9318
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13556 7478 13584 8434
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13556 7342 13584 7414
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13556 6934 13584 7278
rect 13648 7274 13676 8978
rect 13740 8430 13768 8978
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13740 8090 13768 8230
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13818 7984 13874 7993
rect 13818 7919 13820 7928
rect 13872 7919 13874 7928
rect 13820 7890 13872 7896
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13556 6322 13584 6598
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13372 5817 13400 6190
rect 13464 6174 13676 6202
rect 13358 5808 13414 5817
rect 13268 5772 13320 5778
rect 13358 5743 13414 5752
rect 13268 5714 13320 5720
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13188 5001 13216 5238
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13556 5030 13584 5170
rect 13268 5024 13320 5030
rect 13174 4992 13230 5001
rect 13268 4966 13320 4972
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13174 4927 13230 4936
rect 13188 4826 13216 4927
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13096 4706 13124 4762
rect 13096 4678 13216 4706
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12268 2944 12388 2972
rect 12452 3318 12848 3346
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 11428 2032 11480 2038
rect 11428 1974 11480 1980
rect 11244 1624 11296 1630
rect 11244 1566 11296 1572
rect 11072 1414 11192 1442
rect 11072 800 11100 1414
rect 11440 800 11468 1974
rect 11900 800 11928 2246
rect 12268 800 12296 2944
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12360 2446 12388 2790
rect 12452 2650 12480 3318
rect 12912 2922 12940 3470
rect 12992 3460 13044 3466
rect 12992 3402 13044 3408
rect 13004 2990 13032 3402
rect 13096 3126 13124 4014
rect 13188 3890 13216 4678
rect 13280 4078 13308 4966
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13372 3942 13400 4966
rect 13542 4720 13598 4729
rect 13542 4655 13598 4664
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13360 3936 13412 3942
rect 13188 3862 13308 3890
rect 13360 3878 13412 3884
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 13188 3058 13216 3334
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12728 2514 12756 2858
rect 13280 2854 13308 3862
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13372 2990 13400 3538
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13176 2848 13228 2854
rect 12990 2816 13046 2825
rect 13176 2790 13228 2796
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 12990 2751 13046 2760
rect 12806 2680 12862 2689
rect 12806 2615 12808 2624
rect 12860 2615 12862 2624
rect 12808 2586 12860 2592
rect 13004 2514 13032 2751
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12716 2372 12768 2378
rect 12716 2314 12768 2320
rect 12728 800 12756 2314
rect 13096 800 13124 2586
rect 13188 2582 13216 2790
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13464 2514 13492 4082
rect 13556 3602 13584 4655
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13556 2990 13584 3334
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13648 2825 13676 6174
rect 13740 5012 13768 7822
rect 13924 7750 13952 9982
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 14016 8974 14044 9590
rect 14094 9072 14150 9081
rect 14094 9007 14150 9016
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14016 7886 14044 8230
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13818 7576 13874 7585
rect 13818 7511 13874 7520
rect 13832 5846 13860 7511
rect 13924 7342 13952 7686
rect 14016 7410 14044 7822
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 14108 7342 14136 9007
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14200 7290 14228 12158
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14292 11694 14320 12038
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14292 9994 14320 11630
rect 14384 10810 14412 13330
rect 14476 12050 14504 17734
rect 14568 14770 14596 18822
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 14660 14958 14688 18634
rect 14752 15586 14780 19110
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 15304 16998 15332 17682
rect 15488 17241 15516 19246
rect 15672 18426 15700 20266
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15948 19174 15976 20198
rect 16040 19446 16068 20266
rect 16500 19514 16528 20266
rect 16868 19514 16896 20266
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 16946 20088 17002 20097
rect 17236 20058 17264 20198
rect 16946 20023 16948 20032
rect 17000 20023 17002 20032
rect 17224 20052 17276 20058
rect 16948 19994 17000 20000
rect 17224 19994 17276 20000
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 17052 19825 17080 19858
rect 17038 19816 17094 19825
rect 17038 19751 17094 19760
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 17328 19446 17356 19858
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 17316 19440 17368 19446
rect 17316 19382 17368 19388
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 16132 18834 16160 19246
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 15660 18420 15712 18426
rect 15660 18362 15712 18368
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15474 17232 15530 17241
rect 15474 17167 15530 17176
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 15304 16726 15332 16934
rect 15292 16720 15344 16726
rect 15292 16662 15344 16668
rect 15304 16114 15332 16662
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15304 15638 15332 16050
rect 15292 15632 15344 15638
rect 14752 15558 14872 15586
rect 15292 15574 15344 15580
rect 15396 15570 15424 16390
rect 15580 16250 15608 17682
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15764 17066 15792 17614
rect 15856 17610 15884 18158
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 15844 17604 15896 17610
rect 15844 17546 15896 17552
rect 15752 17060 15804 17066
rect 15752 17002 15804 17008
rect 15764 16794 15792 17002
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 14844 15502 14872 15558
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14844 14890 14872 15438
rect 15200 15360 15252 15366
rect 15396 15348 15424 15506
rect 15252 15320 15424 15348
rect 15200 15302 15252 15308
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14646 14784 14702 14793
rect 14568 14742 14646 14770
rect 14646 14719 14702 14728
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14568 13977 14596 14418
rect 14554 13968 14610 13977
rect 14554 13903 14610 13912
rect 14568 13530 14596 13903
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14568 12374 14596 13330
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14476 12022 14596 12050
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14292 9654 14320 9930
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14292 8129 14320 9454
rect 14384 9042 14412 10746
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14278 8120 14334 8129
rect 14278 8055 14334 8064
rect 14108 7002 14136 7278
rect 14200 7262 14320 7290
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14002 6760 14058 6769
rect 13912 6724 13964 6730
rect 14002 6695 14058 6704
rect 13912 6666 13964 6672
rect 13924 6390 13952 6666
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 14016 6118 14044 6695
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13832 5166 13860 5782
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13924 5234 13952 5510
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13924 5098 13952 5170
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13820 5024 13872 5030
rect 13740 4984 13820 5012
rect 13820 4966 13872 4972
rect 13820 4684 13872 4690
rect 13924 4672 13952 5034
rect 14016 4690 14044 5646
rect 14108 5642 14136 6326
rect 14200 6254 14228 7142
rect 14292 6322 14320 7262
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14292 5846 14320 6258
rect 14384 6225 14412 7142
rect 14370 6216 14426 6225
rect 14370 6151 14426 6160
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14280 5840 14332 5846
rect 14280 5782 14332 5788
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14292 5234 14320 5782
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14384 5114 14412 6054
rect 14292 5086 14412 5114
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 13872 4644 13952 4672
rect 14004 4684 14056 4690
rect 13820 4626 13872 4632
rect 14004 4626 14056 4632
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13634 2816 13690 2825
rect 13634 2751 13690 2760
rect 13740 2582 13768 3946
rect 14108 3670 14136 4966
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14200 3738 14228 4422
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 14016 2582 14044 2790
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 14004 2576 14056 2582
rect 14004 2518 14056 2524
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 14188 2508 14240 2514
rect 14292 2496 14320 5086
rect 14372 5024 14424 5030
rect 14370 4992 14372 5001
rect 14424 4992 14426 5001
rect 14370 4927 14426 4936
rect 14370 4720 14426 4729
rect 14370 4655 14426 4664
rect 14384 4622 14412 4655
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14384 2990 14412 4218
rect 14476 4078 14504 11834
rect 14568 11234 14596 12022
rect 14660 11370 14688 14719
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 12374 14780 14214
rect 15120 13892 15332 13920
rect 15120 13802 15148 13892
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 15016 13456 15068 13462
rect 15014 13424 15016 13433
rect 15068 13424 15070 13433
rect 15014 13359 15070 13368
rect 15212 13326 15240 13738
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 14844 13161 14872 13262
rect 14830 13152 14886 13161
rect 14830 13087 14886 13096
rect 14830 13016 14886 13025
rect 14830 12951 14886 12960
rect 14844 12850 14872 12951
rect 15212 12918 15240 13262
rect 15304 13025 15332 13892
rect 15290 13016 15346 13025
rect 15290 12951 15346 12960
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14752 11898 14780 12174
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 14660 11342 14780 11370
rect 14568 11206 14688 11234
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14568 10674 14596 11086
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14568 10266 14596 10406
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14568 9450 14596 9590
rect 14660 9518 14688 11206
rect 14752 10810 14780 11342
rect 15212 11286 15240 12378
rect 15200 11280 15252 11286
rect 14830 11248 14886 11257
rect 15200 11222 15252 11228
rect 14830 11183 14886 11192
rect 14924 11212 14976 11218
rect 14844 11150 14872 11183
rect 14924 11154 14976 11160
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14936 10742 14964 11154
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14752 10146 14780 10542
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 14752 10118 15148 10146
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14568 8838 14596 8978
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14568 6866 14596 8774
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14556 6656 14608 6662
rect 14554 6624 14556 6633
rect 14608 6624 14610 6633
rect 14554 6559 14610 6568
rect 14554 6352 14610 6361
rect 14554 6287 14610 6296
rect 14568 6254 14596 6287
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14568 5273 14596 6190
rect 14554 5264 14610 5273
rect 14554 5199 14610 5208
rect 14568 4690 14596 5199
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14660 4078 14688 9318
rect 14752 9058 14780 9998
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14844 9450 14872 9862
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 15120 9364 15148 10118
rect 15212 9518 15240 10950
rect 15304 10849 15332 10950
rect 15290 10840 15346 10849
rect 15290 10775 15346 10784
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15304 10266 15332 10474
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15120 9336 15332 9364
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14752 9030 14872 9058
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 7954 14780 8774
rect 14844 8362 14872 9030
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 15120 7478 15148 7958
rect 15212 7750 15240 8774
rect 15304 8022 15332 9336
rect 15292 8016 15344 8022
rect 15292 7958 15344 7964
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15304 7206 15332 7958
rect 15396 7857 15424 15320
rect 15764 15026 15792 16730
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15488 14550 15516 14962
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15658 13832 15714 13841
rect 15658 13767 15714 13776
rect 15672 13734 15700 13767
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15580 12628 15608 13670
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 15764 12986 15792 13194
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15580 12600 15700 12628
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15474 11112 15530 11121
rect 15474 11047 15530 11056
rect 15488 10130 15516 11047
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15580 9654 15608 11834
rect 15672 10266 15700 12600
rect 15856 12434 15884 15846
rect 16132 15706 16160 15846
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16212 15360 16264 15366
rect 16212 15302 16264 15308
rect 15948 15026 15976 15302
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 16132 14958 16160 15302
rect 16224 15162 16252 15302
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15948 13530 15976 14758
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16026 13968 16082 13977
rect 16026 13903 16082 13912
rect 16040 13682 16068 13903
rect 16132 13802 16160 14214
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 16040 13654 16160 13682
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 16132 13462 16160 13654
rect 16224 13530 16252 15098
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 16120 13456 16172 13462
rect 16120 13398 16172 13404
rect 16040 12850 16068 13398
rect 16118 13288 16174 13297
rect 16118 13223 16174 13232
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 16040 12434 16068 12650
rect 15764 12406 15884 12434
rect 15948 12406 16068 12434
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15672 9926 15700 10202
rect 15764 10130 15792 12406
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15568 9648 15620 9654
rect 15474 9616 15530 9625
rect 15568 9590 15620 9596
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15474 9551 15530 9560
rect 15488 9382 15516 9551
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15488 8430 15516 8842
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15474 8256 15530 8265
rect 15474 8191 15530 8200
rect 15382 7848 15438 7857
rect 15382 7783 15438 7792
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 15488 6934 15516 8191
rect 15580 8090 15608 9114
rect 15672 9110 15700 9590
rect 15856 9586 15884 12038
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15672 8634 15700 8774
rect 15764 8634 15792 8978
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15856 8362 15884 9522
rect 15948 8480 15976 12406
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 16040 11626 16068 12106
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 16040 10674 16068 11018
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16132 9518 16160 13223
rect 16224 13190 16252 13466
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16316 12220 16344 15846
rect 16408 15162 16436 17682
rect 16592 15201 16620 18566
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16776 17338 16804 17614
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16776 16726 16804 17274
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16578 15192 16634 15201
rect 16396 15156 16448 15162
rect 16578 15127 16634 15136
rect 16396 15098 16448 15104
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16500 13326 16528 14010
rect 16488 13320 16540 13326
rect 16408 13280 16488 13308
rect 16408 13025 16436 13280
rect 16488 13262 16540 13268
rect 16394 13016 16450 13025
rect 16394 12951 16450 12960
rect 16408 12850 16436 12951
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16408 12442 16436 12650
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16500 12374 16528 12854
rect 16592 12434 16620 15127
rect 16948 14884 17000 14890
rect 16948 14826 17000 14832
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16670 14104 16726 14113
rect 16670 14039 16726 14048
rect 16684 14006 16712 14039
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16868 13870 16896 14418
rect 16960 14074 16988 14826
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16868 13530 16896 13806
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16868 12714 16896 13466
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16856 12436 16908 12442
rect 16592 12406 16712 12434
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 16580 12232 16632 12238
rect 16316 12192 16528 12220
rect 16304 11688 16356 11694
rect 16224 11648 16304 11676
rect 16224 10112 16252 11648
rect 16304 11630 16356 11636
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16316 10810 16344 11494
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16408 10742 16436 11494
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16500 10588 16528 12192
rect 16580 12174 16632 12180
rect 16592 11121 16620 12174
rect 16684 12073 16712 12406
rect 16856 12378 16908 12384
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16776 12238 16804 12310
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16670 12064 16726 12073
rect 16670 11999 16726 12008
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 16578 11112 16634 11121
rect 16578 11047 16634 11056
rect 16408 10560 16528 10588
rect 16304 10124 16356 10130
rect 16224 10084 16304 10112
rect 16304 10066 16356 10072
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16316 8537 16344 10066
rect 16302 8528 16358 8537
rect 15948 8452 16252 8480
rect 16302 8463 16358 8472
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 14752 5370 14780 6666
rect 15580 6662 15608 8026
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15672 7206 15700 7822
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 14844 6322 14872 6598
rect 15672 6361 15700 7142
rect 15764 6882 15792 7890
rect 15856 7818 15884 8298
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15764 6854 15884 6882
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15658 6352 15714 6361
rect 14832 6316 14884 6322
rect 15764 6322 15792 6734
rect 15658 6287 15714 6296
rect 15752 6316 15804 6322
rect 14832 6258 14884 6264
rect 15752 6258 15804 6264
rect 14844 6186 14872 6258
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14752 4185 14780 5034
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15304 4282 15332 4422
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 14738 4176 14794 4185
rect 14738 4111 14794 4120
rect 15292 4140 15344 4146
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14568 3670 14596 3878
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 14660 2990 14688 3878
rect 14752 3738 14780 4111
rect 15292 4082 15344 4088
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15120 2990 15148 3538
rect 15212 3194 15240 3878
rect 15304 3466 15332 4082
rect 15396 4010 15424 6054
rect 15488 5914 15516 6190
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15764 5642 15792 6258
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15672 4690 15700 5306
rect 15764 5166 15792 5578
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15856 4457 15884 6854
rect 15842 4448 15898 4457
rect 15842 4383 15898 4392
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15396 3641 15424 3946
rect 15764 3913 15792 4218
rect 15948 4078 15976 8230
rect 16040 7886 16068 8298
rect 16028 7880 16080 7886
rect 16026 7848 16028 7857
rect 16080 7848 16082 7857
rect 16026 7783 16082 7792
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16040 6780 16068 7686
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16132 7002 16160 7142
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 16120 6792 16172 6798
rect 16040 6752 16120 6780
rect 16120 6734 16172 6740
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16040 6254 16068 6598
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 16132 4593 16160 6734
rect 16224 6662 16252 8452
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16224 5710 16252 6598
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16316 5556 16344 8463
rect 16408 7750 16436 10560
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16500 10266 16528 10406
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16684 10146 16712 11562
rect 16762 10976 16818 10985
rect 16762 10911 16818 10920
rect 16776 10810 16804 10911
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16500 10118 16712 10146
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16224 5528 16344 5556
rect 16118 4584 16174 4593
rect 16118 4519 16174 4528
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15750 3904 15806 3913
rect 15750 3839 15806 3848
rect 15382 3632 15438 3641
rect 15382 3567 15438 3576
rect 16224 3534 16252 5528
rect 16408 5370 16436 7346
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16408 5234 16436 5306
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 16408 4758 16436 5170
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16396 4072 16448 4078
rect 16500 4060 16528 10118
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16592 7954 16620 9590
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16684 7834 16712 9522
rect 16764 9512 16816 9518
rect 16762 9480 16764 9489
rect 16816 9480 16818 9489
rect 16762 9415 16818 9424
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16776 8566 16804 8978
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16776 7886 16804 8502
rect 16592 7806 16712 7834
rect 16764 7880 16816 7886
rect 16868 7857 16896 12378
rect 16960 12170 16988 12718
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16960 11286 16988 11630
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16960 9654 16988 10542
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 17052 8945 17080 19110
rect 17236 18630 17264 19246
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17420 18426 17448 20266
rect 17512 19786 17540 22199
rect 17788 20516 17816 22200
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 17960 20528 18012 20534
rect 17788 20488 17960 20516
rect 17960 20470 18012 20476
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17776 20324 17828 20330
rect 17776 20266 17828 20272
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17512 18766 17540 19246
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17604 18698 17632 19110
rect 17696 18986 17724 19858
rect 17788 19514 17816 20266
rect 17880 19922 17908 20334
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 17880 19394 17908 19654
rect 17788 19378 17908 19394
rect 17776 19372 17908 19378
rect 17828 19366 17908 19372
rect 17776 19314 17828 19320
rect 17972 19174 18000 20266
rect 18064 19922 18092 20742
rect 18156 20602 18184 22200
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18616 20534 18644 22200
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 18064 19417 18092 19858
rect 18050 19408 18106 19417
rect 18050 19343 18106 19352
rect 18052 19236 18104 19242
rect 18052 19178 18104 19184
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17696 18958 18000 18986
rect 17592 18692 17644 18698
rect 17592 18634 17644 18640
rect 17972 18630 18000 18958
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 18064 18329 18092 19178
rect 18156 18970 18184 20402
rect 18984 20398 19012 22200
rect 19352 20806 19380 22200
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19720 20466 19748 22200
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 18880 20324 18932 20330
rect 18880 20266 18932 20272
rect 18512 20256 18564 20262
rect 18510 20224 18512 20233
rect 18564 20224 18566 20233
rect 18510 20159 18566 20168
rect 18786 20224 18842 20233
rect 18786 20159 18842 20168
rect 18694 19952 18750 19961
rect 18694 19887 18750 19896
rect 18708 19854 18736 19887
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18418 19408 18474 19417
rect 18418 19343 18474 19352
rect 18432 18970 18460 19343
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18616 18902 18644 19654
rect 18800 19310 18828 20159
rect 18892 19334 18920 20266
rect 18984 19446 19012 20334
rect 19062 20088 19118 20097
rect 19062 20023 19118 20032
rect 19076 19990 19104 20023
rect 19064 19984 19116 19990
rect 19064 19926 19116 19932
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 19076 19446 19104 19790
rect 19168 19514 19196 20334
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19260 19961 19288 19994
rect 19246 19952 19302 19961
rect 19246 19887 19302 19896
rect 19352 19718 19380 20334
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 19430 20224 19486 20233
rect 19430 20159 19486 20168
rect 19444 19922 19472 20159
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 18972 19440 19024 19446
rect 18972 19382 19024 19388
rect 19064 19440 19116 19446
rect 19064 19382 19116 19388
rect 18788 19304 18840 19310
rect 18892 19306 19104 19334
rect 18788 19246 18840 19252
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18604 18896 18656 18902
rect 18708 18873 18736 19110
rect 18604 18838 18656 18844
rect 18694 18864 18750 18873
rect 18694 18799 18750 18808
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18694 18728 18750 18737
rect 18616 18578 18644 18702
rect 18694 18663 18696 18672
rect 18748 18663 18750 18672
rect 18972 18692 19024 18698
rect 18696 18634 18748 18640
rect 18972 18634 19024 18640
rect 18616 18550 18736 18578
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18050 18320 18106 18329
rect 18050 18255 18106 18264
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17420 16658 17448 17070
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17420 15026 17448 16594
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17236 14278 17264 14826
rect 17420 14482 17448 14962
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17406 14240 17462 14249
rect 17236 13326 17264 14214
rect 17512 14226 17540 15574
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17972 14822 18000 15438
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17972 14550 18000 14758
rect 17960 14544 18012 14550
rect 17960 14486 18012 14492
rect 17462 14198 17540 14226
rect 17406 14175 17462 14184
rect 17420 13870 17448 14175
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17420 12782 17448 13194
rect 17788 12986 17816 13262
rect 17880 12986 17908 13330
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17972 12889 18000 13806
rect 18064 13190 18092 15438
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18156 13938 18184 14418
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 18708 13870 18736 18550
rect 18984 18290 19012 18634
rect 19076 18306 19104 19306
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19168 18630 19196 19246
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19260 18970 19288 19178
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 19352 18426 19380 18702
rect 19536 18698 19564 20266
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19720 18970 19748 19858
rect 19904 19854 19932 22607
rect 20074 22200 20130 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21270 22200 21326 23000
rect 21638 22200 21694 23000
rect 22006 22200 22062 23000
rect 22374 22200 22430 23000
rect 22742 22200 22798 23000
rect 20088 20346 20116 22200
rect 20456 21162 20484 22200
rect 20626 21448 20682 21457
rect 20626 21383 20682 21392
rect 20364 21134 20484 21162
rect 20260 20392 20312 20398
rect 19996 20318 20116 20346
rect 20258 20360 20260 20369
rect 20312 20360 20314 20369
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19800 19712 19852 19718
rect 19800 19654 19852 19660
rect 19708 18964 19760 18970
rect 19708 18906 19760 18912
rect 19616 18896 19668 18902
rect 19616 18838 19668 18844
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19628 18426 19656 18838
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19812 18358 19840 19654
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19904 18834 19932 19110
rect 19996 18970 20024 20318
rect 20258 20295 20314 20304
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20088 19990 20116 20198
rect 20076 19984 20128 19990
rect 20076 19926 20128 19932
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19892 18828 19944 18834
rect 19892 18770 19944 18776
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19800 18352 19852 18358
rect 18972 18284 19024 18290
rect 19076 18278 19472 18306
rect 19800 18294 19852 18300
rect 18972 18226 19024 18232
rect 18972 18148 19024 18154
rect 18972 18090 19024 18096
rect 18984 14618 19012 18090
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 18786 14376 18842 14385
rect 18786 14311 18842 14320
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 18340 13530 18368 13738
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18708 13394 18736 13806
rect 18800 13734 18828 14311
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18788 13728 18840 13734
rect 18788 13670 18840 13676
rect 18800 13462 18828 13670
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17958 12880 18014 12889
rect 17958 12815 18014 12824
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17500 12708 17552 12714
rect 17500 12650 17552 12656
rect 17512 12306 17540 12650
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17038 8936 17094 8945
rect 17038 8871 17094 8880
rect 17144 8673 17172 12038
rect 17512 11694 17540 12242
rect 17604 11937 17632 12378
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17774 12064 17830 12073
rect 17590 11928 17646 11937
rect 17590 11863 17646 11872
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17420 11082 17448 11562
rect 17696 11354 17724 12038
rect 17774 11999 17830 12008
rect 17788 11354 17816 11999
rect 18064 11830 18092 12242
rect 18156 11898 18184 13330
rect 18892 13326 18920 13874
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18892 12918 18920 13262
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18788 12368 18840 12374
rect 18510 12336 18566 12345
rect 18788 12310 18840 12316
rect 18510 12271 18566 12280
rect 18524 12170 18552 12271
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18512 12164 18564 12170
rect 18512 12106 18564 12112
rect 18616 12102 18644 12174
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18052 11824 18104 11830
rect 18052 11766 18104 11772
rect 18064 11694 18092 11766
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17314 10704 17370 10713
rect 17314 10639 17370 10648
rect 17592 10668 17644 10674
rect 17328 10606 17356 10639
rect 17592 10610 17644 10616
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17130 8664 17186 8673
rect 17052 8622 17130 8650
rect 16764 7822 16816 7828
rect 16854 7848 16910 7857
rect 16592 6633 16620 7806
rect 16854 7783 16910 7792
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16672 7336 16724 7342
rect 16670 7304 16672 7313
rect 16724 7304 16726 7313
rect 16670 7239 16726 7248
rect 16776 7177 16804 7686
rect 16762 7168 16818 7177
rect 16762 7103 16818 7112
rect 16672 6792 16724 6798
rect 16776 6769 16804 7103
rect 16672 6734 16724 6740
rect 16762 6760 16818 6769
rect 16578 6624 16634 6633
rect 16578 6559 16634 6568
rect 16592 4078 16620 6559
rect 16684 5778 16712 6734
rect 16762 6695 16818 6704
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16776 5098 16804 6054
rect 16868 5778 16896 7783
rect 16948 7268 17000 7274
rect 16948 7210 17000 7216
rect 16960 7002 16988 7210
rect 17052 7041 17080 8622
rect 17130 8599 17186 8608
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17144 7410 17172 8298
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17038 7032 17094 7041
rect 16948 6996 17000 7002
rect 17038 6967 17094 6976
rect 16948 6938 17000 6944
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16960 5166 16988 6054
rect 17052 5914 17080 6054
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17236 5778 17264 10406
rect 17328 10266 17356 10542
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17604 10198 17632 10610
rect 17696 10606 17724 11290
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17788 10538 17816 11290
rect 18064 11150 18092 11290
rect 18708 11234 18736 12038
rect 18800 11665 18828 12310
rect 18892 12102 18920 12718
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18878 11792 18934 11801
rect 18878 11727 18880 11736
rect 18932 11727 18934 11736
rect 18880 11698 18932 11704
rect 18786 11656 18842 11665
rect 18786 11591 18842 11600
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18432 11206 18736 11234
rect 18432 11150 18460 11206
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 17972 10266 18000 10610
rect 18064 10577 18092 11086
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18892 10606 18920 11290
rect 18880 10600 18932 10606
rect 18050 10568 18106 10577
rect 18880 10542 18932 10548
rect 18050 10503 18106 10512
rect 18984 10470 19012 14554
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 19076 13870 19104 14350
rect 19168 14074 19196 14350
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19076 11762 19104 12718
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19260 12442 19288 12582
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19168 11801 19196 12038
rect 19154 11792 19210 11801
rect 19064 11756 19116 11762
rect 19154 11727 19210 11736
rect 19064 11698 19116 11704
rect 19168 11558 19196 11727
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19168 11014 19196 11290
rect 19352 11234 19380 16594
rect 19444 13530 19472 18278
rect 19904 18222 19932 18770
rect 19996 18630 20024 18770
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19720 17882 19748 18158
rect 19708 17876 19760 17882
rect 19708 17818 19760 17824
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19536 14958 19564 15302
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19628 14618 19656 15506
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19536 14074 19564 14418
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 19720 13870 19748 17818
rect 19904 17134 19932 18158
rect 19996 18154 20024 18566
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 20088 17626 20116 19110
rect 20180 18426 20208 20198
rect 20258 20088 20314 20097
rect 20258 20023 20314 20032
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 20168 17740 20220 17746
rect 20168 17682 20220 17688
rect 19996 17598 20116 17626
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 19904 15706 19932 16662
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19444 11354 19472 12650
rect 19996 12442 20024 17598
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19524 11824 19576 11830
rect 19524 11766 19576 11772
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19352 11206 19472 11234
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 19352 10826 19380 11086
rect 19260 10810 19380 10826
rect 19248 10804 19380 10810
rect 19300 10798 19380 10804
rect 19248 10746 19300 10752
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18984 10266 19012 10406
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 17592 10192 17644 10198
rect 19076 10146 19104 10202
rect 17592 10134 17644 10140
rect 17604 10062 17632 10134
rect 18984 10118 19104 10146
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17604 9586 17632 9998
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18984 9722 19012 10118
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17972 9450 18000 9658
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 17328 7002 17356 9318
rect 18524 9178 18552 9318
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17682 8936 17738 8945
rect 17420 7818 17448 8910
rect 17682 8871 17738 8880
rect 17696 8430 17724 8871
rect 17788 8634 17816 9114
rect 18050 9072 18106 9081
rect 18050 9007 18052 9016
rect 18104 9007 18106 9016
rect 18052 8978 18104 8984
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 18234 8936 18290 8945
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17604 8022 17632 8298
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17972 7886 18000 8910
rect 18234 8871 18236 8880
rect 18288 8871 18290 8880
rect 18236 8842 18288 8848
rect 18144 8832 18196 8838
rect 18142 8800 18144 8809
rect 18196 8800 18198 8809
rect 18142 8735 18198 8744
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17776 7472 17828 7478
rect 17590 7440 17646 7449
rect 17776 7414 17828 7420
rect 17590 7375 17646 7384
rect 17604 7342 17632 7375
rect 17788 7342 17816 7414
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17328 6322 17356 6802
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17512 6322 17540 6734
rect 17604 6633 17632 6734
rect 17696 6662 17724 7142
rect 17684 6656 17736 6662
rect 17590 6624 17646 6633
rect 17684 6598 17736 6604
rect 17590 6559 17646 6568
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17420 5914 17448 6054
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17696 5370 17724 6054
rect 17776 5636 17828 5642
rect 17776 5578 17828 5584
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16764 5092 16816 5098
rect 16764 5034 16816 5040
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 16960 4078 16988 4150
rect 16448 4032 16528 4060
rect 16580 4072 16632 4078
rect 16396 4014 16448 4020
rect 16580 4014 16632 4020
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 15292 3460 15344 3466
rect 15292 3402 15344 3408
rect 16316 3398 16344 3878
rect 16396 3460 16448 3466
rect 16396 3402 16448 3408
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15856 2990 15884 3334
rect 15948 2990 15976 3334
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 15108 2984 15160 2990
rect 15384 2984 15436 2990
rect 15108 2926 15160 2932
rect 15382 2952 15384 2961
rect 15844 2984 15896 2990
rect 15436 2952 15438 2961
rect 15844 2926 15896 2932
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 16408 2922 16436 3402
rect 16500 2990 16528 3878
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 15382 2887 15438 2896
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 14464 2848 14516 2854
rect 14370 2816 14426 2825
rect 14464 2790 14516 2796
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 14370 2751 14426 2760
rect 14240 2468 14320 2496
rect 14188 2450 14240 2456
rect 13280 2038 13308 2450
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 13268 2032 13320 2038
rect 13268 1974 13320 1980
rect 13556 800 13584 2382
rect 14384 2310 14412 2751
rect 14476 2582 14504 2790
rect 14464 2576 14516 2582
rect 14752 2564 14780 2790
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 14832 2576 14884 2582
rect 14752 2536 14832 2564
rect 14464 2518 14516 2524
rect 14832 2518 14884 2524
rect 15212 2514 15240 2790
rect 15488 2564 15516 2790
rect 15568 2576 15620 2582
rect 15488 2536 15568 2564
rect 15568 2518 15620 2524
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 14832 2372 14884 2378
rect 14832 2314 14884 2320
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 14372 1488 14424 1494
rect 14372 1430 14424 1436
rect 14004 1420 14056 1426
rect 14004 1362 14056 1368
rect 14016 800 14044 1362
rect 14384 800 14412 1430
rect 14844 800 14872 2314
rect 15304 1170 15332 2382
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 15396 1426 15424 2246
rect 15384 1420 15436 1426
rect 15384 1362 15436 1368
rect 15212 1142 15332 1170
rect 15212 800 15240 1142
rect 15672 800 15700 2858
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 15764 1494 15792 2246
rect 15752 1488 15804 1494
rect 15752 1430 15804 1436
rect 16040 800 16068 2858
rect 16488 2848 16540 2854
rect 16488 2790 16540 2796
rect 16500 800 16528 2790
rect 16592 2582 16620 3062
rect 16776 2582 16804 3878
rect 17052 2650 17080 4966
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17144 3670 17172 3878
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17236 3602 17264 4762
rect 17328 4690 17356 4966
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17684 4684 17736 4690
rect 17684 4626 17736 4632
rect 17696 4282 17724 4626
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17604 3602 17632 4082
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17592 3460 17644 3466
rect 17592 3402 17644 3408
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17328 2774 17356 3334
rect 17604 3194 17632 3402
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17696 2854 17724 3334
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 17328 2746 17448 2774
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 16764 2576 16816 2582
rect 17052 2553 17080 2586
rect 17420 2582 17448 2746
rect 17788 2582 17816 5578
rect 17880 4826 17908 6258
rect 17972 6186 18000 7210
rect 18064 6866 18092 8502
rect 18156 8480 18184 8735
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18156 8452 18368 8480
rect 18340 8362 18368 8452
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18432 7732 18460 8230
rect 18156 7704 18460 7732
rect 18156 7585 18184 7704
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18142 7576 18198 7585
rect 18282 7568 18578 7588
rect 18142 7511 18198 7520
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18340 7002 18368 7142
rect 18418 7032 18474 7041
rect 18328 6996 18380 7002
rect 18418 6967 18474 6976
rect 18328 6938 18380 6944
rect 18432 6866 18460 6967
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 18064 5234 18092 6258
rect 18156 6254 18184 6734
rect 18524 6730 18552 7414
rect 18616 7206 18644 9658
rect 18788 9648 18840 9654
rect 18788 9590 18840 9596
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18616 6361 18644 7142
rect 18602 6352 18658 6361
rect 18602 6287 18658 6296
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18156 5914 18184 6190
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18144 5636 18196 5642
rect 18144 5578 18196 5584
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 18064 4706 18092 5170
rect 18156 5030 18184 5578
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18236 5092 18288 5098
rect 18236 5034 18288 5040
rect 18420 5092 18472 5098
rect 18420 5034 18472 5040
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18156 4865 18184 4966
rect 18142 4856 18198 4865
rect 18142 4791 18198 4800
rect 18064 4678 18184 4706
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 18064 4282 18092 4558
rect 18052 4276 18104 4282
rect 18156 4264 18184 4678
rect 18248 4622 18276 5034
rect 18432 4826 18460 5034
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18708 4264 18736 9454
rect 18800 9178 18828 9590
rect 19076 9518 19104 9998
rect 19064 9512 19116 9518
rect 18984 9472 19064 9500
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18800 7206 18828 8978
rect 18984 8906 19012 9472
rect 19064 9454 19116 9460
rect 19064 9036 19116 9042
rect 19064 8978 19116 8984
rect 18972 8900 19024 8906
rect 18892 8860 18972 8888
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18800 6225 18828 7142
rect 18892 6322 18920 8860
rect 18972 8842 19024 8848
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18984 7886 19012 8434
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18984 7410 19012 7822
rect 19076 7546 19104 8978
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 18970 6896 19026 6905
rect 18970 6831 19026 6840
rect 18984 6798 19012 6831
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 19076 6497 19104 7210
rect 19062 6488 19118 6497
rect 19062 6423 19118 6432
rect 19168 6390 19196 10542
rect 19338 10296 19394 10305
rect 19338 10231 19394 10240
rect 19352 10130 19380 10231
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19444 10010 19472 11206
rect 19352 9982 19472 10010
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 7546 19288 9862
rect 19352 8838 19380 9982
rect 19432 9920 19484 9926
rect 19430 9888 19432 9897
rect 19484 9888 19486 9897
rect 19430 9823 19486 9832
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19340 8424 19392 8430
rect 19338 8392 19340 8401
rect 19392 8392 19394 8401
rect 19338 8327 19394 8336
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19246 7440 19302 7449
rect 19246 7375 19302 7384
rect 19260 7342 19288 7375
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19352 7154 19380 8026
rect 19444 7546 19472 8978
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19536 7342 19564 11766
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19628 8838 19656 11154
rect 19720 11014 19748 12242
rect 19996 11898 20024 12242
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19812 11354 19840 11630
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19708 11008 19760 11014
rect 19708 10950 19760 10956
rect 19996 10810 20024 11154
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19800 10464 19852 10470
rect 19800 10406 19852 10412
rect 19720 9722 19748 10406
rect 19708 9716 19760 9722
rect 19708 9658 19760 9664
rect 19812 9382 19840 10406
rect 19904 10130 19932 10610
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 20088 9194 20116 17478
rect 20180 16998 20208 17682
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20272 15706 20300 20023
rect 20364 18766 20392 21134
rect 20442 21040 20498 21049
rect 20442 20975 20498 20984
rect 20456 20534 20484 20975
rect 20640 20618 20668 21383
rect 20810 20632 20866 20641
rect 20640 20590 20760 20618
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 20536 20528 20588 20534
rect 20536 20470 20588 20476
rect 20444 19984 20496 19990
rect 20444 19926 20496 19932
rect 20456 18970 20484 19926
rect 20548 19786 20576 20470
rect 20732 19990 20760 20590
rect 20810 20567 20866 20576
rect 20824 20534 20852 20567
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20720 19984 20772 19990
rect 20720 19926 20772 19932
rect 20916 19904 20944 22200
rect 21284 21978 21312 22200
rect 21100 21950 21312 21978
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 21008 20097 21036 20334
rect 20994 20088 21050 20097
rect 20994 20023 21050 20032
rect 20996 19916 21048 19922
rect 20916 19876 20996 19904
rect 20536 19780 20588 19786
rect 20536 19722 20588 19728
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20548 18902 20576 19382
rect 20916 19310 20944 19876
rect 20996 19858 21048 19864
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20732 19174 20760 19246
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20548 18442 20576 18838
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20364 18414 20576 18442
rect 20640 18426 20668 18770
rect 20628 18420 20680 18426
rect 20364 17678 20392 18414
rect 20628 18362 20680 18368
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20456 17882 20484 18226
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20640 17882 20668 18022
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 20916 17746 20944 19246
rect 21100 19174 21128 21950
rect 21270 21856 21326 21865
rect 21270 21791 21326 21800
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21192 20233 21220 20402
rect 21178 20224 21234 20233
rect 21178 20159 21234 20168
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21284 18902 21312 21791
rect 21652 20602 21680 22200
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 21362 20360 21418 20369
rect 21362 20295 21418 20304
rect 21548 20324 21600 20330
rect 21376 19514 21404 20295
rect 21548 20266 21600 20272
rect 21456 19712 21508 19718
rect 21560 19689 21588 20266
rect 22020 19990 22048 22200
rect 22388 20398 22416 22200
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22008 19984 22060 19990
rect 22008 19926 22060 19932
rect 21456 19654 21508 19660
rect 21546 19680 21602 19689
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21468 19281 21496 19654
rect 21546 19615 21602 19624
rect 21454 19272 21510 19281
rect 21454 19207 21510 19216
rect 22756 18970 22784 22200
rect 22744 18964 22796 18970
rect 22744 18906 22796 18912
rect 21272 18896 21324 18902
rect 21272 18838 21324 18844
rect 21546 18864 21602 18873
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 21364 18828 21416 18834
rect 21546 18799 21548 18808
rect 21364 18770 21416 18776
rect 21600 18799 21602 18808
rect 21548 18770 21600 18776
rect 21008 18358 21036 18770
rect 21178 18456 21234 18465
rect 21178 18391 21234 18400
rect 21192 18358 21220 18391
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 21180 18352 21232 18358
rect 21180 18294 21232 18300
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20548 16998 20576 17682
rect 20916 17202 20944 17682
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20180 15162 20208 15438
rect 20456 15366 20484 15506
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20456 13462 20484 15302
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 20180 12442 20208 12718
rect 20168 12436 20220 12442
rect 20272 12434 20300 13330
rect 20272 12406 20392 12434
rect 20168 12378 20220 12384
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 19812 9166 20116 9194
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19524 7336 19576 7342
rect 19524 7278 19576 7284
rect 19524 7200 19576 7206
rect 19352 7148 19524 7154
rect 19352 7142 19576 7148
rect 19352 7126 19564 7142
rect 19246 7032 19302 7041
rect 19246 6967 19302 6976
rect 19260 6866 19288 6967
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19156 6384 19208 6390
rect 19156 6326 19208 6332
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 18786 6216 18842 6225
rect 18786 6151 18842 6160
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18800 5166 18828 6054
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18800 4826 18828 4966
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18156 4236 18276 4264
rect 18052 4218 18104 4224
rect 18248 4185 18276 4236
rect 18524 4236 18736 4264
rect 18234 4176 18290 4185
rect 18234 4111 18290 4120
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17972 3482 18000 4014
rect 18248 3602 18276 4111
rect 18524 3602 18552 4236
rect 18800 4162 18828 4626
rect 18892 4554 18920 4762
rect 18880 4548 18932 4554
rect 18880 4490 18932 4496
rect 18708 4134 18828 4162
rect 18708 4026 18736 4134
rect 18616 3998 18736 4026
rect 18786 4040 18842 4049
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 17880 3454 18000 3482
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 17880 3074 17908 3454
rect 18156 3074 18184 3470
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 17880 3058 18092 3074
rect 18156 3058 18276 3074
rect 17880 3052 18104 3058
rect 17880 3046 18052 3052
rect 18156 3052 18288 3058
rect 18156 3046 18236 3052
rect 18052 2994 18104 3000
rect 18236 2994 18288 3000
rect 17866 2952 17922 2961
rect 17866 2887 17922 2896
rect 18144 2916 18196 2922
rect 17880 2666 17908 2887
rect 18144 2858 18196 2864
rect 17960 2848 18012 2854
rect 18012 2808 18092 2836
rect 17960 2790 18012 2796
rect 17880 2650 18000 2666
rect 17880 2644 18012 2650
rect 17880 2638 17960 2644
rect 17960 2586 18012 2592
rect 17408 2576 17460 2582
rect 16764 2518 16816 2524
rect 17038 2544 17094 2553
rect 17408 2518 17460 2524
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17038 2479 17094 2488
rect 18064 2446 18092 2808
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 16868 800 16896 2314
rect 17328 800 17356 2382
rect 17684 2372 17736 2378
rect 17684 2314 17736 2320
rect 17696 800 17724 2314
rect 18156 800 18184 2858
rect 18248 2854 18276 2994
rect 18420 2984 18472 2990
rect 18472 2944 18552 2972
rect 18420 2926 18472 2932
rect 18524 2854 18552 2944
rect 18236 2848 18288 2854
rect 18512 2848 18564 2854
rect 18236 2790 18288 2796
rect 18510 2816 18512 2825
rect 18564 2816 18566 2825
rect 18248 2514 18276 2790
rect 18510 2751 18566 2760
rect 18616 2650 18644 3998
rect 18786 3975 18842 3984
rect 18880 4004 18932 4010
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18708 2553 18736 3878
rect 18800 3738 18828 3975
rect 18880 3946 18932 3952
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18694 2544 18750 2553
rect 18236 2508 18288 2514
rect 18694 2479 18750 2488
rect 18236 2450 18288 2456
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18616 800 18644 2246
rect 18800 1329 18828 3334
rect 18892 3194 18920 3946
rect 18880 3188 18932 3194
rect 18880 3130 18932 3136
rect 18892 2446 18920 3130
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18984 2281 19012 6054
rect 19260 5896 19288 6258
rect 19260 5868 19472 5896
rect 19064 5840 19116 5846
rect 19062 5808 19064 5817
rect 19116 5808 19118 5817
rect 19062 5743 19118 5752
rect 19156 5772 19208 5778
rect 19208 5732 19380 5760
rect 19156 5714 19208 5720
rect 19352 5370 19380 5732
rect 19444 5710 19472 5868
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19064 4820 19116 4826
rect 19064 4762 19116 4768
rect 19076 3618 19104 4762
rect 19260 4690 19288 5306
rect 19536 5302 19564 7126
rect 19628 5370 19656 8774
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19720 7954 19748 8366
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 19524 5296 19576 5302
rect 19444 5256 19524 5284
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19168 4593 19196 4626
rect 19154 4584 19210 4593
rect 19154 4519 19210 4528
rect 19156 4480 19208 4486
rect 19340 4480 19392 4486
rect 19208 4440 19288 4468
rect 19156 4422 19208 4428
rect 19154 4176 19210 4185
rect 19154 4111 19156 4120
rect 19208 4111 19210 4120
rect 19156 4082 19208 4088
rect 19260 4060 19288 4440
rect 19340 4422 19392 4428
rect 19352 4282 19380 4422
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19340 4072 19392 4078
rect 19260 4032 19340 4060
rect 19340 4014 19392 4020
rect 19076 3590 19196 3618
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 19076 2650 19104 3334
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 19168 2530 19196 3590
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19248 3120 19300 3126
rect 19248 3062 19300 3068
rect 19260 2689 19288 3062
rect 19352 3058 19380 3334
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19444 2961 19472 5256
rect 19524 5238 19576 5244
rect 19628 4740 19656 5306
rect 19536 4712 19656 4740
rect 19536 4049 19564 4712
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19522 4040 19578 4049
rect 19522 3975 19578 3984
rect 19524 3936 19576 3942
rect 19522 3904 19524 3913
rect 19576 3904 19578 3913
rect 19522 3839 19578 3848
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19536 2990 19564 3470
rect 19628 3466 19656 4558
rect 19720 3942 19748 7278
rect 19812 4842 19840 9166
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 19904 8498 19932 8978
rect 20180 8634 20208 12038
rect 20272 11898 20300 12106
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 20272 9625 20300 11018
rect 20258 9616 20314 9625
rect 20258 9551 20314 9560
rect 20260 9444 20312 9450
rect 20260 9386 20312 9392
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 19892 8492 19944 8498
rect 19892 8434 19944 8440
rect 19904 7750 19932 8434
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19996 8090 20024 8230
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19904 6798 19932 7686
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 19996 6866 20024 7414
rect 20180 7290 20208 7890
rect 20088 7262 20208 7290
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19890 6352 19946 6361
rect 19890 6287 19946 6296
rect 19904 4978 19932 6287
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 19996 5914 20024 6054
rect 20088 5914 20116 7262
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20180 7002 20208 7142
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 20272 6662 20300 9386
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20180 6186 20208 6598
rect 20258 6488 20314 6497
rect 20258 6423 20314 6432
rect 20168 6180 20220 6186
rect 20168 6122 20220 6128
rect 20166 6080 20222 6089
rect 20166 6015 20222 6024
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19996 5273 20024 5646
rect 20180 5642 20208 6015
rect 20168 5636 20220 5642
rect 20168 5578 20220 5584
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 19982 5264 20038 5273
rect 19982 5199 20038 5208
rect 20088 5098 20116 5510
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 20180 5030 20208 5306
rect 20168 5024 20220 5030
rect 19904 4950 20116 4978
rect 20168 4966 20220 4972
rect 19982 4856 20038 4865
rect 19812 4814 19932 4842
rect 19800 4548 19852 4554
rect 19800 4490 19852 4496
rect 19812 4146 19840 4490
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19616 3460 19668 3466
rect 19616 3402 19668 3408
rect 19616 3120 19668 3126
rect 19616 3062 19668 3068
rect 19524 2984 19576 2990
rect 19430 2952 19486 2961
rect 19340 2916 19392 2922
rect 19524 2926 19576 2932
rect 19430 2887 19486 2896
rect 19340 2858 19392 2864
rect 19246 2680 19302 2689
rect 19352 2650 19380 2858
rect 19628 2774 19656 3062
rect 19720 2854 19748 3878
rect 19812 3534 19840 4082
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19904 2922 19932 4814
rect 19982 4791 19984 4800
rect 20036 4791 20038 4800
rect 19984 4762 20036 4768
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19996 4146 20024 4626
rect 20088 4570 20116 4950
rect 20272 4826 20300 6423
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20088 4542 20300 4570
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20088 4146 20116 4422
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19996 3194 20024 3538
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19800 2916 19852 2922
rect 19800 2858 19852 2864
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19444 2746 19656 2774
rect 19246 2615 19302 2624
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19444 2582 19472 2746
rect 19432 2576 19484 2582
rect 19168 2502 19380 2530
rect 19432 2518 19484 2524
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 19352 2394 19380 2502
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 19720 2394 19748 2450
rect 18970 2272 19026 2281
rect 18970 2207 19026 2216
rect 18786 1320 18842 1329
rect 18786 1255 18842 1264
rect 19260 1170 19288 2382
rect 19352 2366 19748 2394
rect 19616 2304 19668 2310
rect 19616 2246 19668 2252
rect 19628 1170 19656 2246
rect 18984 1142 19288 1170
rect 19444 1142 19656 1170
rect 18984 800 19012 1142
rect 19444 800 19472 1142
rect 19812 800 19840 2858
rect 20180 2825 20208 4422
rect 20272 3466 20300 4542
rect 20260 3460 20312 3466
rect 20260 3402 20312 3408
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 20166 2816 20222 2825
rect 20166 2751 20222 2760
rect 20272 800 20300 2858
rect 20364 2650 20392 12406
rect 20444 11688 20496 11694
rect 20442 11656 20444 11665
rect 20496 11656 20498 11665
rect 20442 11591 20498 11600
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20456 10810 20484 11154
rect 20444 10804 20496 10810
rect 20444 10746 20496 10752
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 20456 9654 20484 10066
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 20548 9330 20576 16934
rect 20824 16794 20852 17070
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20640 15162 20668 15982
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 21180 15972 21232 15978
rect 21180 15914 21232 15920
rect 20732 15706 20760 15914
rect 20904 15904 20956 15910
rect 21192 15881 21220 15914
rect 20904 15846 20956 15852
rect 21178 15872 21234 15881
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20916 15638 20944 15846
rect 21178 15807 21234 15816
rect 20904 15632 20956 15638
rect 20904 15574 20956 15580
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20640 14278 20668 14418
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20640 12102 20668 14214
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20732 11898 20760 12650
rect 20824 12238 20852 14758
rect 21178 14648 21234 14657
rect 21178 14583 21234 14592
rect 21192 14550 21220 14583
rect 21180 14544 21232 14550
rect 21180 14486 21232 14492
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20456 9302 20576 9330
rect 20456 7886 20484 9302
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20548 8430 20576 8774
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20456 7002 20484 7686
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 20456 6497 20484 6666
rect 20442 6488 20498 6497
rect 20442 6423 20498 6432
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20456 5370 20484 5578
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 20548 4214 20576 7890
rect 20640 5914 20668 11562
rect 20732 10810 20760 11630
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20824 11014 20852 11494
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20916 9466 20944 13126
rect 21178 12472 21234 12481
rect 21178 12407 21234 12416
rect 21192 12374 21220 12407
rect 21180 12368 21232 12374
rect 21180 12310 21232 12316
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 21008 11898 21036 12242
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 21100 10538 21128 11086
rect 21088 10532 21140 10538
rect 21088 10474 21140 10480
rect 21180 10532 21232 10538
rect 21180 10474 21232 10480
rect 21100 10441 21128 10474
rect 21086 10432 21142 10441
rect 21086 10367 21142 10376
rect 21192 10169 21220 10474
rect 21178 10160 21234 10169
rect 21178 10095 21234 10104
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 20732 9438 20944 9466
rect 20732 8673 20760 9438
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20718 8664 20774 8673
rect 20718 8599 20774 8608
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20732 7818 20760 8434
rect 20824 7993 20852 8774
rect 20916 8634 20944 9318
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20810 7984 20866 7993
rect 20810 7919 20866 7928
rect 20812 7880 20864 7886
rect 20810 7848 20812 7857
rect 20864 7848 20866 7857
rect 20720 7812 20772 7818
rect 20810 7783 20866 7792
rect 20720 7754 20772 7760
rect 20732 7410 20760 7754
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20732 6390 20760 7346
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20812 6928 20864 6934
rect 20916 6914 20944 7142
rect 20864 6886 20944 6914
rect 20812 6870 20864 6876
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20626 5808 20682 5817
rect 20626 5743 20682 5752
rect 20536 4208 20588 4214
rect 20536 4150 20588 4156
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 20456 2553 20484 4014
rect 20548 3670 20576 4150
rect 20536 3664 20588 3670
rect 20536 3606 20588 3612
rect 20640 3602 20668 5743
rect 20732 4826 20760 6054
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20824 5166 20852 5306
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 20916 4978 20944 6886
rect 21008 6730 21036 9318
rect 21100 9178 21128 9522
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21088 8356 21140 8362
rect 21088 8298 21140 8304
rect 21100 6866 21128 8298
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 21088 6180 21140 6186
rect 21088 6122 21140 6128
rect 21100 6089 21128 6122
rect 21192 6118 21220 8366
rect 21284 8004 21312 18022
rect 21376 17338 21404 18770
rect 21548 18148 21600 18154
rect 21548 18090 21600 18096
rect 21560 18057 21588 18090
rect 21546 18048 21602 18057
rect 21546 17983 21602 17992
rect 21546 17640 21602 17649
rect 21546 17575 21548 17584
rect 21600 17575 21602 17584
rect 22008 17604 22060 17610
rect 21548 17546 21600 17552
rect 22008 17546 22060 17552
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21640 17264 21692 17270
rect 21546 17232 21602 17241
rect 21640 17206 21692 17212
rect 21546 17167 21548 17176
rect 21600 17167 21602 17176
rect 21548 17138 21600 17144
rect 21364 17060 21416 17066
rect 21364 17002 21416 17008
rect 21376 16250 21404 17002
rect 21546 16824 21602 16833
rect 21546 16759 21602 16768
rect 21560 16726 21588 16759
rect 21548 16720 21600 16726
rect 21548 16662 21600 16668
rect 21546 16280 21602 16289
rect 21364 16244 21416 16250
rect 21546 16215 21602 16224
rect 21364 16186 21416 16192
rect 21560 16182 21588 16215
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 21546 15464 21602 15473
rect 21546 15399 21548 15408
rect 21600 15399 21602 15408
rect 21548 15370 21600 15376
rect 21546 15056 21602 15065
rect 21546 14991 21548 15000
rect 21600 14991 21602 15000
rect 21548 14962 21600 14968
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21376 14074 21404 14418
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 21560 14249 21588 14282
rect 21546 14240 21602 14249
rect 21546 14175 21602 14184
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21548 13864 21600 13870
rect 21546 13832 21548 13841
rect 21600 13832 21602 13841
rect 21364 13796 21416 13802
rect 21546 13767 21602 13776
rect 21364 13738 21416 13744
rect 21376 12986 21404 13738
rect 21546 13424 21602 13433
rect 21546 13359 21548 13368
rect 21600 13359 21602 13368
rect 21548 13330 21600 13336
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21546 12880 21602 12889
rect 21546 12815 21548 12824
rect 21600 12815 21602 12824
rect 21548 12786 21600 12792
rect 21652 12434 21680 17206
rect 22020 12434 22048 17546
rect 21652 12406 21772 12434
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21456 12096 21508 12102
rect 21560 12073 21588 12106
rect 21456 12038 21508 12044
rect 21546 12064 21602 12073
rect 21468 11914 21496 12038
rect 21546 11999 21602 12008
rect 21468 11886 21588 11914
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21468 11218 21496 11698
rect 21560 11626 21588 11886
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21560 11257 21588 11562
rect 21546 11248 21602 11257
rect 21456 11212 21508 11218
rect 21546 11183 21602 11192
rect 21456 11154 21508 11160
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21376 10520 21404 11086
rect 21468 10849 21496 11154
rect 21454 10840 21510 10849
rect 21454 10775 21510 10784
rect 21456 10532 21508 10538
rect 21376 10492 21456 10520
rect 21456 10474 21508 10480
rect 21362 10024 21418 10033
rect 21362 9959 21364 9968
rect 21416 9959 21418 9968
rect 21364 9930 21416 9936
rect 21468 9489 21496 10474
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21546 9888 21602 9897
rect 21546 9823 21602 9832
rect 21560 9518 21588 9823
rect 21548 9512 21600 9518
rect 21454 9480 21510 9489
rect 21548 9454 21600 9460
rect 21454 9415 21510 9424
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21376 9110 21404 9318
rect 21364 9104 21416 9110
rect 21652 9081 21680 10066
rect 21364 9046 21416 9052
rect 21638 9072 21694 9081
rect 21548 9036 21600 9042
rect 21638 9007 21694 9016
rect 21548 8978 21600 8984
rect 21560 8673 21588 8978
rect 21744 8922 21772 12406
rect 21652 8894 21772 8922
rect 21928 12406 22048 12434
rect 21546 8664 21602 8673
rect 21546 8599 21602 8608
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 21560 8265 21588 8366
rect 21546 8256 21602 8265
rect 21546 8191 21602 8200
rect 21560 8090 21588 8191
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21284 7976 21404 8004
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21180 6112 21232 6118
rect 21086 6080 21142 6089
rect 21180 6054 21232 6060
rect 21086 6015 21142 6024
rect 21284 5522 21312 7822
rect 20824 4950 20944 4978
rect 21008 5494 21312 5522
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20824 4214 20852 4950
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20916 4282 20944 4626
rect 21008 4486 21036 5494
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21088 5160 21140 5166
rect 21284 5137 21312 5170
rect 21088 5102 21140 5108
rect 21270 5128 21326 5137
rect 21100 4672 21128 5102
rect 21270 5063 21326 5072
rect 21100 4644 21220 4672
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20812 4208 20864 4214
rect 20812 4150 20864 4156
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20640 3058 20668 3334
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20442 2544 20498 2553
rect 20442 2479 20498 2488
rect 20456 1465 20484 2479
rect 20442 1456 20498 1465
rect 20442 1391 20498 1400
rect 20640 800 20668 2858
rect 20732 1329 20760 4014
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20812 3120 20864 3126
rect 20916 3097 20944 3878
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 20996 3460 21048 3466
rect 20996 3402 21048 3408
rect 20812 3062 20864 3068
rect 20902 3088 20958 3097
rect 20824 2582 20852 3062
rect 20902 3023 20958 3032
rect 21008 2582 21036 3402
rect 20812 2576 20864 2582
rect 20812 2518 20864 2524
rect 20996 2576 21048 2582
rect 20996 2518 21048 2524
rect 21100 2446 21128 3470
rect 21192 3097 21220 4644
rect 21272 4072 21324 4078
rect 21270 4040 21272 4049
rect 21324 4040 21326 4049
rect 21270 3975 21326 3984
rect 21376 3670 21404 7976
rect 21546 7848 21602 7857
rect 21546 7783 21602 7792
rect 21560 7342 21588 7783
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21456 7200 21508 7206
rect 21454 7168 21456 7177
rect 21508 7168 21510 7177
rect 21454 7103 21510 7112
rect 21560 7002 21588 7278
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21548 6180 21600 6186
rect 21548 6122 21600 6128
rect 21456 5772 21508 5778
rect 21456 5714 21508 5720
rect 21468 5273 21496 5714
rect 21560 5681 21588 6122
rect 21546 5672 21602 5681
rect 21546 5607 21602 5616
rect 21548 5568 21600 5574
rect 21548 5510 21600 5516
rect 21454 5264 21510 5273
rect 21454 5199 21510 5208
rect 21456 5092 21508 5098
rect 21456 5034 21508 5040
rect 21468 4865 21496 5034
rect 21454 4856 21510 4865
rect 21454 4791 21510 4800
rect 21456 4684 21508 4690
rect 21456 4626 21508 4632
rect 21468 4457 21496 4626
rect 21454 4448 21510 4457
rect 21454 4383 21510 4392
rect 21456 4276 21508 4282
rect 21456 4218 21508 4224
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 21178 3088 21234 3097
rect 21178 3023 21234 3032
rect 21468 2938 21496 4218
rect 21560 4078 21588 5510
rect 21548 4072 21600 4078
rect 21548 4014 21600 4020
rect 21560 3641 21588 4014
rect 21546 3632 21602 3641
rect 21652 3602 21680 8894
rect 21824 7472 21876 7478
rect 21824 7414 21876 7420
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21546 3567 21602 3576
rect 21640 3596 21692 3602
rect 21640 3538 21692 3544
rect 21468 2910 21588 2938
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 20718 1320 20774 1329
rect 20718 1255 20774 1264
rect 2962 640 3018 649
rect 2962 575 3018 584
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20732 649 20760 1255
rect 21100 800 21128 2382
rect 21468 800 21496 2790
rect 21560 1873 21588 2910
rect 21744 2281 21772 5102
rect 21836 4826 21864 7414
rect 21928 5370 21956 12406
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 22006 10296 22062 10305
rect 22006 10231 22062 10240
rect 22020 9674 22048 10231
rect 22020 9646 22140 9674
rect 22006 6488 22062 6497
rect 22006 6423 22008 6432
rect 22060 6423 22062 6432
rect 22008 6394 22060 6400
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 21730 2272 21786 2281
rect 21730 2207 21786 2216
rect 21546 1864 21602 1873
rect 21546 1799 21602 1808
rect 21836 1057 21864 4558
rect 22112 3942 22140 9646
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 21916 3460 21968 3466
rect 21916 3402 21968 3408
rect 21822 1048 21878 1057
rect 21822 983 21878 992
rect 21928 800 21956 3402
rect 22204 2990 22232 10950
rect 22284 5296 22336 5302
rect 22284 5238 22336 5244
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 20718 640 20774 649
rect 20718 575 20774 584
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21914 0 21970 800
rect 22020 241 22048 2790
rect 22296 800 22324 5238
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22756 800 22784 3334
rect 22006 232 22062 241
rect 22006 167 22062 176
rect 22282 0 22338 800
rect 22742 0 22798 800
<< via2 >>
rect 1398 22616 1454 22672
rect 2962 22208 3018 22264
rect 1490 20204 1492 20224
rect 1492 20204 1544 20224
rect 1544 20204 1546 20224
rect 1490 20168 1546 20204
rect 1490 19660 1492 19680
rect 1492 19660 1544 19680
rect 1544 19660 1546 19680
rect 1490 19624 1546 19660
rect 1398 19252 1400 19272
rect 1400 19252 1452 19272
rect 1452 19252 1454 19272
rect 1398 19216 1454 19252
rect 1858 20596 1914 20632
rect 1858 20576 1860 20596
rect 1860 20576 1912 20596
rect 1912 20576 1914 20596
rect 2226 20984 2282 21040
rect 1398 18844 1400 18864
rect 1400 18844 1452 18864
rect 1452 18844 1454 18864
rect 1398 18808 1454 18844
rect 1950 19252 1952 19272
rect 1952 19252 2004 19272
rect 2004 19252 2006 19272
rect 1950 19216 2006 19252
rect 1858 18420 1914 18456
rect 1858 18400 1860 18420
rect 1860 18400 1912 18420
rect 1912 18400 1914 18420
rect 17498 22208 17554 22264
rect 2870 21800 2926 21856
rect 2778 21392 2834 21448
rect 2134 18808 2190 18864
rect 2042 18264 2098 18320
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 2778 19896 2834 19952
rect 2594 18672 2650 18728
rect 2502 18536 2558 18592
rect 3790 19352 3846 19408
rect 2410 17856 2466 17912
rect 1766 17604 1822 17640
rect 1766 17584 1768 17604
rect 1768 17584 1820 17604
rect 1820 17584 1822 17604
rect 1490 17176 1546 17232
rect 1490 16768 1546 16824
rect 1490 16224 1546 16280
rect 2962 17584 3018 17640
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4710 20204 4712 20224
rect 4712 20204 4764 20224
rect 4764 20204 4766 20224
rect 4710 20168 4766 20204
rect 3974 19216 4030 19272
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 3882 18572 3884 18592
rect 3884 18572 3936 18592
rect 3936 18572 3938 18592
rect 3882 18536 3938 18572
rect 3974 18128 4030 18184
rect 4342 19080 4398 19136
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4526 17876 4582 17912
rect 4526 17856 4528 17876
rect 4528 17856 4580 17876
rect 4580 17856 4582 17876
rect 1858 15816 1914 15872
rect 1398 15428 1454 15464
rect 1398 15408 1400 15428
rect 1400 15408 1452 15428
rect 1452 15408 1454 15428
rect 1398 15020 1454 15056
rect 1398 15000 1400 15020
rect 1400 15000 1452 15020
rect 1452 15000 1454 15020
rect 1858 14612 1914 14648
rect 1858 14592 1860 14612
rect 1860 14592 1912 14612
rect 1912 14592 1914 14612
rect 1490 14220 1492 14240
rect 1492 14220 1544 14240
rect 1544 14220 1546 14240
rect 1490 14184 1546 14220
rect 1766 13812 1768 13832
rect 1768 13812 1820 13832
rect 1820 13812 1822 13832
rect 1766 13776 1822 13812
rect 1398 13368 1454 13424
rect 1858 12824 1914 12880
rect 1398 12416 1454 12472
rect 1490 12008 1546 12064
rect 1582 11736 1638 11792
rect 1398 10784 1454 10840
rect 1490 10376 1546 10432
rect 1950 9288 2006 9344
rect 1766 8628 1822 8664
rect 1766 8608 1768 8628
rect 1768 8608 1820 8628
rect 1820 8608 1822 8628
rect 1858 8508 1860 8528
rect 1860 8508 1912 8528
rect 1912 8508 1914 8528
rect 1858 8472 1914 8508
rect 1674 8064 1730 8120
rect 1490 7792 1546 7848
rect 1490 6976 1546 7032
rect 1490 6860 1546 6896
rect 2134 7112 2190 7168
rect 1490 6840 1492 6860
rect 1492 6840 1544 6860
rect 1544 6840 1546 6860
rect 1122 6160 1178 6216
rect 938 5752 994 5808
rect 938 1808 994 1864
rect 1214 5616 1270 5672
rect 1306 5208 1362 5264
rect 1306 4392 1362 4448
rect 1306 4020 1308 4040
rect 1308 4020 1360 4040
rect 1360 4020 1362 4040
rect 1306 3984 1362 4020
rect 1490 6024 1546 6080
rect 1766 4936 1822 4992
rect 1582 3984 1638 4040
rect 1398 3596 1454 3632
rect 1398 3576 1400 3596
rect 1400 3576 1452 3596
rect 1452 3576 1454 3596
rect 1122 992 1178 1048
rect 2042 5072 2098 5128
rect 1766 3032 1822 3088
rect 2042 3032 2098 3088
rect 2410 7248 2466 7304
rect 2318 6996 2374 7032
rect 2318 6976 2320 6996
rect 2320 6976 2372 6996
rect 2372 6976 2374 6996
rect 2870 9152 2926 9208
rect 3330 13524 3386 13560
rect 3330 13504 3332 13524
rect 3332 13504 3384 13524
rect 3384 13504 3386 13524
rect 3882 16496 3938 16552
rect 3606 12688 3662 12744
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 3974 14356 3976 14376
rect 3976 14356 4028 14376
rect 4028 14356 4030 14376
rect 3974 14320 4030 14356
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 3974 13640 4030 13696
rect 4158 13640 4214 13696
rect 3882 12552 3938 12608
rect 3330 11212 3386 11248
rect 3330 11192 3332 11212
rect 3332 11192 3384 11212
rect 3384 11192 3386 11212
rect 3422 9868 3424 9888
rect 3424 9868 3476 9888
rect 3476 9868 3478 9888
rect 3422 9832 3478 9868
rect 4066 11600 4122 11656
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4710 13796 4766 13832
rect 4710 13776 4712 13796
rect 4712 13776 4764 13796
rect 4764 13776 4766 13796
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4250 11600 4306 11656
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 3238 9460 3240 9480
rect 3240 9460 3292 9480
rect 3292 9460 3294 9480
rect 3238 9424 3294 9460
rect 3146 9036 3202 9072
rect 3146 9016 3148 9036
rect 3148 9016 3200 9036
rect 3200 9016 3202 9036
rect 2962 7792 3018 7848
rect 3330 8900 3386 8936
rect 4250 10648 4306 10704
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 3330 8880 3332 8900
rect 3332 8880 3384 8900
rect 3384 8880 3386 8900
rect 3514 8200 3570 8256
rect 3238 7384 3294 7440
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4986 14220 4988 14240
rect 4988 14220 5040 14240
rect 5040 14220 5042 14240
rect 4986 14184 5042 14220
rect 5630 20168 5686 20224
rect 5446 18536 5502 18592
rect 5170 14220 5172 14240
rect 5172 14220 5224 14240
rect 5224 14220 5226 14240
rect 5170 14184 5226 14220
rect 5446 17856 5502 17912
rect 6366 20340 6368 20360
rect 6368 20340 6420 20360
rect 6420 20340 6422 20360
rect 6366 20304 6422 20340
rect 4894 8336 4950 8392
rect 3606 6704 3662 6760
rect 2870 6024 2926 6080
rect 2778 4800 2834 4856
rect 3238 6432 3294 6488
rect 2502 3460 2558 3496
rect 2502 3440 2504 3460
rect 2504 3440 2556 3460
rect 2556 3440 2558 3460
rect 2410 2796 2412 2816
rect 2412 2796 2464 2816
rect 2464 2796 2466 2816
rect 2410 2760 2466 2796
rect 1306 176 1362 232
rect 3238 5616 3294 5672
rect 3790 6432 3846 6488
rect 4158 7928 4214 7984
rect 4066 6840 4122 6896
rect 3790 5364 3846 5400
rect 5262 13776 5318 13832
rect 5354 13640 5410 13696
rect 5354 12960 5410 13016
rect 5538 13504 5594 13560
rect 5538 12280 5594 12336
rect 5354 12164 5410 12200
rect 5354 12144 5356 12164
rect 5356 12144 5408 12164
rect 5408 12144 5410 12164
rect 5262 11872 5318 11928
rect 5722 13504 5778 13560
rect 5906 13368 5962 13424
rect 5814 13096 5870 13152
rect 5630 10648 5686 10704
rect 5538 10532 5594 10568
rect 5538 10512 5540 10532
rect 5540 10512 5592 10532
rect 5592 10512 5594 10532
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4802 7520 4858 7576
rect 4250 6196 4252 6216
rect 4252 6196 4304 6216
rect 4304 6196 4306 6216
rect 4250 6160 4306 6196
rect 4158 5888 4214 5944
rect 3790 5344 3792 5364
rect 3792 5344 3844 5364
rect 3844 5344 3846 5364
rect 3698 5208 3754 5264
rect 4618 6840 4674 6896
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4802 6332 4804 6352
rect 4804 6332 4856 6352
rect 4856 6332 4858 6352
rect 4802 6296 4858 6332
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 3882 4800 3938 4856
rect 3238 2916 3294 2952
rect 3238 2896 3240 2916
rect 3240 2896 3292 2916
rect 3292 2896 3294 2916
rect 3790 3576 3846 3632
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4618 4120 4674 4176
rect 4434 3884 4436 3904
rect 4436 3884 4488 3904
rect 4488 3884 4490 3904
rect 4434 3848 4490 3884
rect 4710 3612 4712 3632
rect 4712 3612 4764 3632
rect 4764 3612 4766 3632
rect 4710 3576 4766 3612
rect 4250 1400 4306 1456
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 5906 12280 5962 12336
rect 6274 18400 6330 18456
rect 6182 14592 6238 14648
rect 6182 13776 6238 13832
rect 6090 11192 6146 11248
rect 5354 7520 5410 7576
rect 7010 19352 7066 19408
rect 6826 18400 6882 18456
rect 7286 19760 7342 19816
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 8206 19624 8262 19680
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7562 17720 7618 17776
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7746 17620 7748 17640
rect 7748 17620 7800 17640
rect 7800 17620 7802 17640
rect 7746 17584 7802 17620
rect 8206 17176 8262 17232
rect 7286 16904 7342 16960
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 6642 12688 6698 12744
rect 6550 12416 6606 12472
rect 6826 13640 6882 13696
rect 6918 13504 6974 13560
rect 6734 12280 6790 12336
rect 8574 19760 8630 19816
rect 8574 17484 8576 17504
rect 8576 17484 8628 17504
rect 8628 17484 8630 17504
rect 8574 17448 8630 17484
rect 8574 16496 8630 16552
rect 8482 16088 8538 16144
rect 5354 6840 5410 6896
rect 5538 6704 5594 6760
rect 5906 7112 5962 7168
rect 5630 6568 5686 6624
rect 5538 5908 5594 5944
rect 5538 5888 5540 5908
rect 5540 5888 5592 5908
rect 5592 5888 5594 5908
rect 6274 6976 6330 7032
rect 5998 6432 6054 6488
rect 4986 3884 4988 3904
rect 4988 3884 5040 3904
rect 5040 3884 5042 3904
rect 4986 3848 5042 3884
rect 4986 3712 5042 3768
rect 4802 2252 4804 2272
rect 4804 2252 4856 2272
rect 4856 2252 4858 2272
rect 4802 2216 4858 2252
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 5354 4256 5410 4312
rect 5354 3304 5410 3360
rect 5354 2760 5410 2816
rect 5814 5616 5870 5672
rect 5998 5616 6054 5672
rect 5814 4528 5870 4584
rect 5814 4392 5870 4448
rect 5722 3712 5778 3768
rect 6182 6704 6238 6760
rect 6182 6160 6238 6216
rect 6182 5772 6238 5808
rect 6182 5752 6184 5772
rect 6184 5752 6236 5772
rect 6236 5752 6238 5772
rect 6274 5480 6330 5536
rect 6274 4528 6330 4584
rect 6182 2760 6238 2816
rect 6458 10260 6514 10296
rect 6458 10240 6460 10260
rect 6460 10240 6512 10260
rect 6512 10240 6514 10260
rect 7010 12552 7066 12608
rect 6826 10104 6882 10160
rect 6826 9560 6882 9616
rect 6734 9288 6790 9344
rect 7010 9560 7066 9616
rect 7010 9460 7012 9480
rect 7012 9460 7064 9480
rect 7064 9460 7066 9480
rect 7010 9424 7066 9460
rect 6918 8064 6974 8120
rect 6642 6840 6698 6896
rect 6918 7520 6974 7576
rect 6918 7248 6974 7304
rect 6458 6160 6514 6216
rect 5538 2352 5594 2408
rect 6734 6160 6790 6216
rect 6734 5344 6790 5400
rect 7010 4664 7066 4720
rect 7562 14592 7618 14648
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7838 14884 7894 14920
rect 7838 14864 7840 14884
rect 7840 14864 7892 14884
rect 7892 14864 7894 14884
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7562 13368 7618 13424
rect 7562 12844 7618 12880
rect 7562 12824 7564 12844
rect 7564 12824 7616 12844
rect 7616 12824 7618 12844
rect 7378 12008 7434 12064
rect 7378 11464 7434 11520
rect 7378 11056 7434 11112
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 8206 12688 8262 12744
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 8114 12280 8170 12336
rect 8574 12960 8630 13016
rect 9126 19624 9182 19680
rect 8850 18536 8906 18592
rect 8666 12688 8722 12744
rect 8942 15816 8998 15872
rect 8850 13912 8906 13968
rect 8758 12552 8814 12608
rect 8850 12416 8906 12472
rect 8482 12280 8538 12336
rect 8390 12008 8446 12064
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7746 10784 7802 10840
rect 7562 10684 7564 10704
rect 7564 10684 7616 10704
rect 7616 10684 7618 10704
rect 7562 10648 7618 10684
rect 7562 10412 7564 10432
rect 7564 10412 7616 10432
rect 7616 10412 7618 10432
rect 7562 10376 7618 10412
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 8298 10920 8354 10976
rect 7930 9696 7986 9752
rect 8022 9424 8078 9480
rect 8298 9968 8354 10024
rect 8298 9424 8354 9480
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 8574 12008 8630 12064
rect 8390 8608 8446 8664
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 8758 11600 8814 11656
rect 8758 11500 8760 11520
rect 8760 11500 8812 11520
rect 8812 11500 8814 11520
rect 8758 11464 8814 11500
rect 8666 10920 8722 10976
rect 8850 10784 8906 10840
rect 8758 10376 8814 10432
rect 8758 7384 8814 7440
rect 7562 6704 7618 6760
rect 7378 6296 7434 6352
rect 7562 6296 7618 6352
rect 7194 5616 7250 5672
rect 7562 5752 7618 5808
rect 7746 6296 7802 6352
rect 8022 6160 8078 6216
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7470 5344 7526 5400
rect 7378 5072 7434 5128
rect 6734 2760 6790 2816
rect 7286 4936 7342 4992
rect 7286 4664 7342 4720
rect 7194 2508 7250 2544
rect 7194 2488 7196 2508
rect 7196 2488 7248 2508
rect 7248 2488 7250 2508
rect 8022 5480 8078 5536
rect 7930 5208 7986 5264
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 8482 6568 8538 6624
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 8666 5208 8722 5264
rect 8574 4392 8630 4448
rect 8758 4664 8814 4720
rect 8666 4120 8722 4176
rect 9218 18536 9274 18592
rect 9586 18164 9588 18184
rect 9588 18164 9640 18184
rect 9640 18164 9642 18184
rect 9586 18128 9642 18164
rect 9218 14048 9274 14104
rect 9126 12960 9182 13016
rect 9586 14884 9642 14920
rect 9586 14864 9588 14884
rect 9588 14864 9640 14884
rect 9640 14864 9642 14884
rect 9310 12960 9366 13016
rect 9218 12552 9274 12608
rect 9126 12416 9182 12472
rect 9034 11872 9090 11928
rect 9402 12416 9458 12472
rect 9218 10240 9274 10296
rect 9310 10104 9366 10160
rect 9218 9444 9274 9480
rect 9218 9424 9220 9444
rect 9220 9424 9272 9444
rect 9272 9424 9274 9444
rect 8942 6296 8998 6352
rect 8942 5480 8998 5536
rect 7470 3304 7526 3360
rect 7562 3032 7618 3088
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 8666 2896 8722 2952
rect 9310 9288 9366 9344
rect 9218 8608 9274 8664
rect 9310 8472 9366 8528
rect 9494 12008 9550 12064
rect 10046 20304 10102 20360
rect 9862 17448 9918 17504
rect 9770 17176 9826 17232
rect 9862 16496 9918 16552
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 9862 13676 9864 13696
rect 9864 13676 9916 13696
rect 9916 13676 9918 13696
rect 9862 13640 9918 13676
rect 9770 12416 9826 12472
rect 9494 11500 9496 11520
rect 9496 11500 9548 11520
rect 9548 11500 9550 11520
rect 9494 11464 9550 11500
rect 9678 11464 9734 11520
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 10414 16668 10416 16688
rect 10416 16668 10468 16688
rect 10468 16668 10470 16688
rect 10414 16632 10470 16668
rect 10138 13776 10194 13832
rect 10322 14728 10378 14784
rect 10414 14048 10470 14104
rect 11058 17584 11114 17640
rect 11058 16632 11114 16688
rect 11150 16496 11206 16552
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11334 17620 11336 17640
rect 11336 17620 11388 17640
rect 11388 17620 11390 17640
rect 11334 17584 11390 17620
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 10506 13776 10562 13832
rect 10230 12824 10286 12880
rect 10138 12552 10194 12608
rect 10046 11464 10102 11520
rect 9862 11328 9918 11384
rect 9770 10920 9826 10976
rect 9494 10376 9550 10432
rect 9494 9152 9550 9208
rect 9678 9152 9734 9208
rect 9402 8200 9458 8256
rect 9310 7928 9366 7984
rect 9126 7112 9182 7168
rect 9126 6432 9182 6488
rect 9126 6296 9182 6352
rect 9402 6604 9404 6624
rect 9404 6604 9456 6624
rect 9456 6604 9458 6624
rect 9402 6568 9458 6604
rect 9586 8744 9642 8800
rect 9678 7928 9734 7984
rect 10138 10376 10194 10432
rect 10138 8780 10140 8800
rect 10140 8780 10192 8800
rect 10192 8780 10194 8800
rect 10138 8744 10194 8780
rect 10046 8608 10102 8664
rect 10138 8336 10194 8392
rect 9954 7248 10010 7304
rect 9862 6704 9918 6760
rect 9678 6432 9734 6488
rect 9678 6024 9734 6080
rect 9678 5480 9734 5536
rect 9954 5888 10010 5944
rect 9954 4528 10010 4584
rect 9770 3188 9826 3224
rect 9770 3168 9772 3188
rect 9772 3168 9824 3188
rect 9824 3168 9826 3188
rect 9678 2760 9734 2816
rect 9586 2216 9642 2272
rect 10046 3440 10102 3496
rect 10782 14048 10838 14104
rect 10598 13504 10654 13560
rect 10506 12824 10562 12880
rect 10414 12008 10470 12064
rect 10598 11600 10654 11656
rect 10598 11464 10654 11520
rect 10506 11328 10562 11384
rect 10690 10920 10746 10976
rect 10598 10784 10654 10840
rect 10598 10376 10654 10432
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 10966 14320 11022 14376
rect 10874 13504 10930 13560
rect 11426 14476 11482 14512
rect 11426 14456 11428 14476
rect 11428 14456 11480 14476
rect 11480 14456 11482 14476
rect 11058 12960 11114 13016
rect 10966 12824 11022 12880
rect 10966 12588 10968 12608
rect 10968 12588 11020 12608
rect 11020 12588 11022 12608
rect 10966 12552 11022 12588
rect 10966 12416 11022 12472
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11334 13640 11390 13696
rect 11426 13504 11482 13560
rect 11426 13232 11482 13288
rect 19890 22616 19946 22672
rect 11978 15444 11980 15464
rect 11980 15444 12032 15464
rect 12032 15444 12034 15464
rect 11978 15408 12034 15444
rect 11886 15308 11888 15328
rect 11888 15308 11940 15328
rect 11940 15308 11942 15328
rect 11886 15272 11942 15308
rect 11978 15136 12034 15192
rect 12162 14728 12218 14784
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11610 12416 11666 12472
rect 11150 12008 11206 12064
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 13818 16768 13874 16824
rect 12346 15156 12402 15192
rect 12346 15136 12348 15156
rect 12348 15136 12400 15156
rect 12400 15136 12402 15156
rect 12346 14320 12402 14376
rect 12806 14048 12862 14104
rect 13450 15408 13506 15464
rect 13726 14184 13782 14240
rect 11794 11736 11850 11792
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11058 10240 11114 10296
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11058 8744 11114 8800
rect 10414 7656 10470 7712
rect 10322 6860 10378 6896
rect 10322 6840 10324 6860
rect 10324 6840 10376 6860
rect 10376 6840 10378 6860
rect 10598 7692 10600 7712
rect 10600 7692 10652 7712
rect 10652 7692 10654 7712
rect 10598 7656 10654 7692
rect 10598 7520 10654 7576
rect 10598 7248 10654 7304
rect 10598 7148 10600 7168
rect 10600 7148 10652 7168
rect 10652 7148 10654 7168
rect 10598 7112 10654 7148
rect 10506 6840 10562 6896
rect 10874 8200 10930 8256
rect 10598 5888 10654 5944
rect 10322 5072 10378 5128
rect 11702 9424 11758 9480
rect 12162 10920 12218 10976
rect 11978 10804 12034 10840
rect 11978 10784 11980 10804
rect 11980 10784 12032 10804
rect 12032 10784 12034 10804
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11150 7656 11206 7712
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11426 7248 11482 7304
rect 10874 6976 10930 7032
rect 10782 5480 10838 5536
rect 10322 2896 10378 2952
rect 10506 2488 10562 2544
rect 10966 6704 11022 6760
rect 11150 6976 11206 7032
rect 11426 6976 11482 7032
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11150 6432 11206 6488
rect 11426 6296 11482 6352
rect 11610 6160 11666 6216
rect 11518 5888 11574 5944
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11150 3576 11206 3632
rect 11058 3440 11114 3496
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11886 5888 11942 5944
rect 11794 4392 11850 4448
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11334 3032 11390 3088
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12162 9832 12218 9888
rect 12162 8744 12218 8800
rect 12346 11736 12402 11792
rect 13358 12824 13414 12880
rect 13450 12436 13506 12472
rect 13450 12416 13452 12436
rect 13452 12416 13504 12436
rect 13504 12416 13506 12436
rect 13174 11600 13230 11656
rect 12622 10920 12678 10976
rect 12254 7656 12310 7712
rect 12530 9832 12586 9888
rect 12438 9716 12494 9752
rect 12438 9696 12440 9716
rect 12440 9696 12492 9716
rect 12492 9696 12494 9716
rect 12622 9560 12678 9616
rect 12714 9424 12770 9480
rect 12622 9152 12678 9208
rect 12530 8880 12586 8936
rect 12346 6976 12402 7032
rect 12622 7792 12678 7848
rect 12162 6704 12218 6760
rect 12438 6840 12494 6896
rect 12162 5616 12218 5672
rect 12346 5908 12402 5944
rect 12530 6568 12586 6624
rect 12346 5888 12348 5908
rect 12348 5888 12400 5908
rect 12400 5888 12402 5908
rect 11886 3032 11942 3088
rect 13358 11056 13414 11112
rect 13174 10376 13230 10432
rect 12990 9560 13046 9616
rect 12990 9288 13046 9344
rect 12990 8064 13046 8120
rect 13266 8744 13322 8800
rect 13082 7692 13084 7712
rect 13084 7692 13136 7712
rect 13136 7692 13138 7712
rect 13082 7656 13138 7692
rect 12806 5752 12862 5808
rect 12162 3884 12164 3904
rect 12164 3884 12216 3904
rect 12216 3884 12218 3904
rect 12162 3848 12218 3884
rect 12346 4428 12348 4448
rect 12348 4428 12400 4448
rect 12400 4428 12402 4448
rect 12346 4392 12402 4428
rect 12438 3712 12494 3768
rect 13358 7520 13414 7576
rect 13266 6704 13322 6760
rect 13174 6160 13230 6216
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 14094 13096 14150 13152
rect 13818 7948 13874 7984
rect 13818 7928 13820 7948
rect 13820 7928 13872 7948
rect 13872 7928 13874 7948
rect 13358 5752 13414 5808
rect 13174 4936 13230 4992
rect 13542 4664 13598 4720
rect 12990 2760 13046 2816
rect 12806 2644 12862 2680
rect 12806 2624 12808 2644
rect 12808 2624 12860 2644
rect 12860 2624 12862 2644
rect 14094 9016 14150 9072
rect 13818 7520 13874 7576
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 16946 20052 17002 20088
rect 16946 20032 16948 20052
rect 16948 20032 17000 20052
rect 17000 20032 17002 20052
rect 17038 19760 17094 19816
rect 15474 17176 15530 17232
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14646 14728 14702 14784
rect 14554 13912 14610 13968
rect 14278 8064 14334 8120
rect 14002 6704 14058 6760
rect 14370 6160 14426 6216
rect 13634 2760 13690 2816
rect 14370 4972 14372 4992
rect 14372 4972 14424 4992
rect 14424 4972 14426 4992
rect 14370 4936 14426 4972
rect 14370 4664 14426 4720
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 15014 13404 15016 13424
rect 15016 13404 15068 13424
rect 15068 13404 15070 13424
rect 15014 13368 15070 13404
rect 14830 13096 14886 13152
rect 14830 12960 14886 13016
rect 15290 12960 15346 13016
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14830 11192 14886 11248
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14554 6604 14556 6624
rect 14556 6604 14608 6624
rect 14608 6604 14610 6624
rect 14554 6568 14610 6604
rect 14554 6296 14610 6352
rect 14554 5208 14610 5264
rect 15290 10784 15346 10840
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 15658 13776 15714 13832
rect 15474 11056 15530 11112
rect 16026 13912 16082 13968
rect 16118 13232 16174 13288
rect 15474 9560 15530 9616
rect 15474 8200 15530 8256
rect 15382 7792 15438 7848
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 16578 15136 16634 15192
rect 16394 12960 16450 13016
rect 16670 14048 16726 14104
rect 16670 12008 16726 12064
rect 16578 11056 16634 11112
rect 16302 8472 16358 8528
rect 15658 6296 15714 6352
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14738 4120 14794 4176
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 15842 4392 15898 4448
rect 16026 7828 16028 7848
rect 16028 7828 16080 7848
rect 16080 7828 16082 7848
rect 16026 7792 16082 7828
rect 16762 10920 16818 10976
rect 16118 4528 16174 4584
rect 15750 3848 15806 3904
rect 15382 3576 15438 3632
rect 16762 9460 16764 9480
rect 16764 9460 16816 9480
rect 16816 9460 16818 9480
rect 16762 9424 16818 9460
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18050 19352 18106 19408
rect 18510 20204 18512 20224
rect 18512 20204 18564 20224
rect 18564 20204 18566 20224
rect 18510 20168 18566 20204
rect 18786 20168 18842 20224
rect 18694 19896 18750 19952
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18418 19352 18474 19408
rect 19062 20032 19118 20088
rect 19246 19896 19302 19952
rect 19430 20168 19486 20224
rect 18694 18808 18750 18864
rect 18694 18692 18750 18728
rect 18694 18672 18696 18692
rect 18696 18672 18748 18692
rect 18748 18672 18750 18692
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18050 18264 18106 18320
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 17406 14184 17462 14240
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 20626 21392 20682 21448
rect 20258 20340 20260 20360
rect 20260 20340 20312 20360
rect 20312 20340 20314 20360
rect 20258 20304 20314 20340
rect 18786 14320 18842 14376
rect 17958 12824 18014 12880
rect 17038 8880 17094 8936
rect 17590 11872 17646 11928
rect 17774 12008 17830 12064
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18510 12280 18566 12336
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 17314 10648 17370 10704
rect 16854 7792 16910 7848
rect 16670 7284 16672 7304
rect 16672 7284 16724 7304
rect 16724 7284 16726 7304
rect 16670 7248 16726 7284
rect 16762 7112 16818 7168
rect 16578 6568 16634 6624
rect 16762 6704 16818 6760
rect 17130 8608 17186 8664
rect 17038 6976 17094 7032
rect 18878 11756 18934 11792
rect 18878 11736 18880 11756
rect 18880 11736 18932 11756
rect 18932 11736 18934 11756
rect 18786 11600 18842 11656
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18050 10512 18106 10568
rect 19154 11736 19210 11792
rect 20258 20032 20314 20088
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 17682 8880 17738 8936
rect 18050 9036 18106 9072
rect 18050 9016 18052 9036
rect 18052 9016 18104 9036
rect 18104 9016 18106 9036
rect 18234 8900 18290 8936
rect 18234 8880 18236 8900
rect 18236 8880 18288 8900
rect 18288 8880 18290 8900
rect 18142 8780 18144 8800
rect 18144 8780 18196 8800
rect 18196 8780 18198 8800
rect 18142 8744 18198 8780
rect 17590 7384 17646 7440
rect 17590 6568 17646 6624
rect 15382 2932 15384 2952
rect 15384 2932 15436 2952
rect 15436 2932 15438 2952
rect 15382 2896 15438 2932
rect 14370 2760 14426 2816
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18142 7520 18198 7576
rect 18418 6976 18474 7032
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18602 6296 18658 6352
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18142 4800 18198 4856
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18970 6840 19026 6896
rect 19062 6432 19118 6488
rect 19338 10240 19394 10296
rect 19430 9868 19432 9888
rect 19432 9868 19484 9888
rect 19484 9868 19486 9888
rect 19430 9832 19486 9868
rect 19338 8372 19340 8392
rect 19340 8372 19392 8392
rect 19392 8372 19394 8392
rect 19338 8336 19394 8372
rect 19246 7384 19302 7440
rect 20442 20984 20498 21040
rect 20810 20576 20866 20632
rect 20994 20032 21050 20088
rect 21270 21800 21326 21856
rect 21178 20168 21234 20224
rect 21362 20304 21418 20360
rect 21546 19624 21602 19680
rect 21454 19216 21510 19272
rect 21546 18828 21602 18864
rect 21546 18808 21548 18828
rect 21548 18808 21600 18828
rect 21600 18808 21602 18828
rect 21178 18400 21234 18456
rect 19246 6976 19302 7032
rect 18786 6160 18842 6216
rect 18234 4120 18290 4176
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 17866 2896 17922 2952
rect 17038 2488 17094 2544
rect 18510 2796 18512 2816
rect 18512 2796 18564 2816
rect 18564 2796 18566 2816
rect 18510 2760 18566 2796
rect 18786 3984 18842 4040
rect 18694 2488 18750 2544
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 19062 5788 19064 5808
rect 19064 5788 19116 5808
rect 19116 5788 19118 5808
rect 19062 5752 19118 5788
rect 19154 4528 19210 4584
rect 19154 4140 19210 4176
rect 19154 4120 19156 4140
rect 19156 4120 19208 4140
rect 19208 4120 19210 4140
rect 19522 3984 19578 4040
rect 19522 3884 19524 3904
rect 19524 3884 19576 3904
rect 19576 3884 19578 3904
rect 19522 3848 19578 3884
rect 20258 9560 20314 9616
rect 19890 6296 19946 6352
rect 20258 6432 20314 6488
rect 20166 6024 20222 6080
rect 19982 5208 20038 5264
rect 19430 2896 19486 2952
rect 19246 2624 19302 2680
rect 19982 4820 20038 4856
rect 19982 4800 19984 4820
rect 19984 4800 20036 4820
rect 20036 4800 20038 4820
rect 18970 2216 19026 2272
rect 18786 1264 18842 1320
rect 20166 2760 20222 2816
rect 20442 11636 20444 11656
rect 20444 11636 20496 11656
rect 20496 11636 20498 11656
rect 20442 11600 20498 11636
rect 21178 15816 21234 15872
rect 21178 14592 21234 14648
rect 20442 6432 20498 6488
rect 21178 12416 21234 12472
rect 21086 10376 21142 10432
rect 21178 10104 21234 10160
rect 20718 8608 20774 8664
rect 20810 7928 20866 7984
rect 20810 7828 20812 7848
rect 20812 7828 20864 7848
rect 20864 7828 20866 7848
rect 20810 7792 20866 7828
rect 20626 5752 20682 5808
rect 21546 17992 21602 18048
rect 21546 17604 21602 17640
rect 21546 17584 21548 17604
rect 21548 17584 21600 17604
rect 21600 17584 21602 17604
rect 21546 17196 21602 17232
rect 21546 17176 21548 17196
rect 21548 17176 21600 17196
rect 21600 17176 21602 17196
rect 21546 16768 21602 16824
rect 21546 16224 21602 16280
rect 21546 15428 21602 15464
rect 21546 15408 21548 15428
rect 21548 15408 21600 15428
rect 21600 15408 21602 15428
rect 21546 15020 21602 15056
rect 21546 15000 21548 15020
rect 21548 15000 21600 15020
rect 21600 15000 21602 15020
rect 21546 14184 21602 14240
rect 21546 13812 21548 13832
rect 21548 13812 21600 13832
rect 21600 13812 21602 13832
rect 21546 13776 21602 13812
rect 21546 13388 21602 13424
rect 21546 13368 21548 13388
rect 21548 13368 21600 13388
rect 21600 13368 21602 13388
rect 21546 12844 21602 12880
rect 21546 12824 21548 12844
rect 21548 12824 21600 12844
rect 21600 12824 21602 12844
rect 21546 12008 21602 12064
rect 21546 11192 21602 11248
rect 21454 10784 21510 10840
rect 21362 9988 21418 10024
rect 21362 9968 21364 9988
rect 21364 9968 21416 9988
rect 21416 9968 21418 9988
rect 21546 9832 21602 9888
rect 21454 9424 21510 9480
rect 21638 9016 21694 9072
rect 21546 8608 21602 8664
rect 21546 8200 21602 8256
rect 21086 6024 21142 6080
rect 21270 5072 21326 5128
rect 20442 2488 20498 2544
rect 20442 1400 20498 1456
rect 20902 3032 20958 3088
rect 21270 4020 21272 4040
rect 21272 4020 21324 4040
rect 21324 4020 21326 4040
rect 21270 3984 21326 4020
rect 21546 7792 21602 7848
rect 21454 7148 21456 7168
rect 21456 7148 21508 7168
rect 21508 7148 21510 7168
rect 21454 7112 21510 7148
rect 21546 5616 21602 5672
rect 21454 5208 21510 5264
rect 21454 4800 21510 4856
rect 21454 4392 21510 4448
rect 21178 3032 21234 3088
rect 21546 3576 21602 3632
rect 20718 1264 20774 1320
rect 2962 584 3018 640
rect 22006 10240 22062 10296
rect 22006 6452 22062 6488
rect 22006 6432 22008 6452
rect 22008 6432 22060 6452
rect 22060 6432 22062 6452
rect 21730 2216 21786 2272
rect 21546 1808 21602 1864
rect 21822 992 21878 1048
rect 20718 584 20774 640
rect 22006 176 22062 232
<< metal3 >>
rect 0 22674 800 22704
rect 1393 22674 1459 22677
rect 0 22672 1459 22674
rect 0 22616 1398 22672
rect 1454 22616 1459 22672
rect 0 22614 1459 22616
rect 0 22584 800 22614
rect 1393 22611 1459 22614
rect 19885 22674 19951 22677
rect 22200 22674 23000 22704
rect 19885 22672 23000 22674
rect 19885 22616 19890 22672
rect 19946 22616 23000 22672
rect 19885 22614 23000 22616
rect 19885 22611 19951 22614
rect 22200 22584 23000 22614
rect 0 22266 800 22296
rect 2957 22266 3023 22269
rect 0 22264 3023 22266
rect 0 22208 2962 22264
rect 3018 22208 3023 22264
rect 0 22206 3023 22208
rect 0 22176 800 22206
rect 2957 22203 3023 22206
rect 17493 22266 17559 22269
rect 22200 22266 23000 22296
rect 17493 22264 23000 22266
rect 17493 22208 17498 22264
rect 17554 22208 23000 22264
rect 17493 22206 23000 22208
rect 17493 22203 17559 22206
rect 22200 22176 23000 22206
rect 0 21858 800 21888
rect 2865 21858 2931 21861
rect 0 21856 2931 21858
rect 0 21800 2870 21856
rect 2926 21800 2931 21856
rect 0 21798 2931 21800
rect 0 21768 800 21798
rect 2865 21795 2931 21798
rect 21265 21858 21331 21861
rect 22200 21858 23000 21888
rect 21265 21856 23000 21858
rect 21265 21800 21270 21856
rect 21326 21800 23000 21856
rect 21265 21798 23000 21800
rect 21265 21795 21331 21798
rect 22200 21768 23000 21798
rect 0 21450 800 21480
rect 2773 21450 2839 21453
rect 0 21448 2839 21450
rect 0 21392 2778 21448
rect 2834 21392 2839 21448
rect 0 21390 2839 21392
rect 0 21360 800 21390
rect 2773 21387 2839 21390
rect 20621 21450 20687 21453
rect 22200 21450 23000 21480
rect 20621 21448 23000 21450
rect 20621 21392 20626 21448
rect 20682 21392 23000 21448
rect 20621 21390 23000 21392
rect 20621 21387 20687 21390
rect 22200 21360 23000 21390
rect 0 21042 800 21072
rect 2221 21042 2287 21045
rect 0 21040 2287 21042
rect 0 20984 2226 21040
rect 2282 20984 2287 21040
rect 0 20982 2287 20984
rect 0 20952 800 20982
rect 2221 20979 2287 20982
rect 20437 21042 20503 21045
rect 22200 21042 23000 21072
rect 20437 21040 23000 21042
rect 20437 20984 20442 21040
rect 20498 20984 23000 21040
rect 20437 20982 23000 20984
rect 20437 20979 20503 20982
rect 22200 20952 23000 20982
rect 4409 20704 4729 20705
rect 0 20634 800 20664
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 1853 20634 1919 20637
rect 0 20632 1919 20634
rect 0 20576 1858 20632
rect 1914 20576 1919 20632
rect 0 20574 1919 20576
rect 0 20544 800 20574
rect 1853 20571 1919 20574
rect 20805 20634 20871 20637
rect 22200 20634 23000 20664
rect 20805 20632 23000 20634
rect 20805 20576 20810 20632
rect 20866 20576 23000 20632
rect 20805 20574 23000 20576
rect 20805 20571 20871 20574
rect 22200 20544 23000 20574
rect 6361 20362 6427 20365
rect 10041 20362 10107 20365
rect 6361 20360 10107 20362
rect 6361 20304 6366 20360
rect 6422 20304 10046 20360
rect 10102 20304 10107 20360
rect 6361 20302 10107 20304
rect 6361 20299 6427 20302
rect 10041 20299 10107 20302
rect 20253 20362 20319 20365
rect 21357 20362 21423 20365
rect 20253 20360 21423 20362
rect 20253 20304 20258 20360
rect 20314 20304 21362 20360
rect 21418 20304 21423 20360
rect 20253 20302 21423 20304
rect 20253 20299 20319 20302
rect 21357 20299 21423 20302
rect 0 20226 800 20256
rect 1485 20226 1551 20229
rect 0 20224 1551 20226
rect 0 20168 1490 20224
rect 1546 20168 1551 20224
rect 0 20166 1551 20168
rect 0 20136 800 20166
rect 1485 20163 1551 20166
rect 4705 20226 4771 20229
rect 5625 20226 5691 20229
rect 4705 20224 5691 20226
rect 4705 20168 4710 20224
rect 4766 20168 5630 20224
rect 5686 20168 5691 20224
rect 4705 20166 5691 20168
rect 4705 20163 4771 20166
rect 5625 20163 5691 20166
rect 18505 20226 18571 20229
rect 18781 20226 18847 20229
rect 19425 20226 19491 20229
rect 18505 20224 19491 20226
rect 18505 20168 18510 20224
rect 18566 20168 18786 20224
rect 18842 20168 19430 20224
rect 19486 20168 19491 20224
rect 18505 20166 19491 20168
rect 18505 20163 18571 20166
rect 18781 20163 18847 20166
rect 19425 20163 19491 20166
rect 21173 20226 21239 20229
rect 22200 20226 23000 20256
rect 21173 20224 23000 20226
rect 21173 20168 21178 20224
rect 21234 20168 23000 20224
rect 21173 20166 23000 20168
rect 21173 20163 21239 20166
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 22200 20136 23000 20166
rect 14805 20095 15125 20096
rect 16941 20090 17007 20093
rect 19057 20090 19123 20093
rect 16941 20088 19123 20090
rect 16941 20032 16946 20088
rect 17002 20032 19062 20088
rect 19118 20032 19123 20088
rect 16941 20030 19123 20032
rect 16941 20027 17007 20030
rect 19057 20027 19123 20030
rect 20253 20090 20319 20093
rect 20989 20090 21055 20093
rect 20253 20088 21055 20090
rect 20253 20032 20258 20088
rect 20314 20032 20994 20088
rect 21050 20032 21055 20088
rect 20253 20030 21055 20032
rect 20253 20027 20319 20030
rect 20989 20027 21055 20030
rect 2773 19954 2839 19957
rect 18689 19954 18755 19957
rect 19241 19954 19307 19957
rect 2773 19952 18755 19954
rect 2773 19896 2778 19952
rect 2834 19896 18694 19952
rect 18750 19896 18755 19952
rect 2773 19894 18755 19896
rect 2773 19891 2839 19894
rect 18689 19891 18755 19894
rect 19198 19952 19307 19954
rect 19198 19896 19246 19952
rect 19302 19896 19307 19952
rect 19198 19891 19307 19896
rect 7281 19818 7347 19821
rect 8569 19818 8635 19821
rect 7281 19816 8635 19818
rect 7281 19760 7286 19816
rect 7342 19760 8574 19816
rect 8630 19760 8635 19816
rect 7281 19758 8635 19760
rect 7281 19755 7347 19758
rect 8569 19755 8635 19758
rect 17033 19818 17099 19821
rect 19198 19818 19258 19891
rect 17033 19816 19258 19818
rect 17033 19760 17038 19816
rect 17094 19760 19258 19816
rect 17033 19758 19258 19760
rect 17033 19755 17099 19758
rect 0 19682 800 19712
rect 1485 19682 1551 19685
rect 0 19680 1551 19682
rect 0 19624 1490 19680
rect 1546 19624 1551 19680
rect 0 19622 1551 19624
rect 0 19592 800 19622
rect 1485 19619 1551 19622
rect 8201 19682 8267 19685
rect 9121 19682 9187 19685
rect 8201 19680 9187 19682
rect 8201 19624 8206 19680
rect 8262 19624 9126 19680
rect 9182 19624 9187 19680
rect 8201 19622 9187 19624
rect 8201 19619 8267 19622
rect 9121 19619 9187 19622
rect 21541 19682 21607 19685
rect 22200 19682 23000 19712
rect 21541 19680 23000 19682
rect 21541 19624 21546 19680
rect 21602 19624 23000 19680
rect 21541 19622 23000 19624
rect 21541 19619 21607 19622
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 22200 19592 23000 19622
rect 18270 19551 18590 19552
rect 3785 19410 3851 19413
rect 7005 19410 7071 19413
rect 3785 19408 7071 19410
rect 3785 19352 3790 19408
rect 3846 19352 7010 19408
rect 7066 19352 7071 19408
rect 3785 19350 7071 19352
rect 3785 19347 3851 19350
rect 7005 19347 7071 19350
rect 18045 19410 18111 19413
rect 18413 19410 18479 19413
rect 18045 19408 18479 19410
rect 18045 19352 18050 19408
rect 18106 19352 18418 19408
rect 18474 19352 18479 19408
rect 18045 19350 18479 19352
rect 18045 19347 18111 19350
rect 18413 19347 18479 19350
rect 0 19274 800 19304
rect 1393 19274 1459 19277
rect 0 19272 1459 19274
rect 0 19216 1398 19272
rect 1454 19216 1459 19272
rect 0 19214 1459 19216
rect 0 19184 800 19214
rect 1393 19211 1459 19214
rect 1945 19274 2011 19277
rect 3969 19274 4035 19277
rect 1945 19272 4035 19274
rect 1945 19216 1950 19272
rect 2006 19216 3974 19272
rect 4030 19216 4035 19272
rect 1945 19214 4035 19216
rect 1945 19211 2011 19214
rect 3969 19211 4035 19214
rect 21449 19274 21515 19277
rect 22200 19274 23000 19304
rect 21449 19272 23000 19274
rect 21449 19216 21454 19272
rect 21510 19216 23000 19272
rect 21449 19214 23000 19216
rect 21449 19211 21515 19214
rect 22200 19184 23000 19214
rect 4337 19138 4403 19141
rect 7230 19138 7236 19140
rect 4337 19136 7236 19138
rect 4337 19080 4342 19136
rect 4398 19080 7236 19136
rect 4337 19078 7236 19080
rect 4337 19075 4403 19078
rect 7230 19076 7236 19078
rect 7300 19076 7306 19140
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 0 18866 800 18896
rect 1393 18866 1459 18869
rect 0 18864 1459 18866
rect 0 18808 1398 18864
rect 1454 18808 1459 18864
rect 0 18806 1459 18808
rect 0 18776 800 18806
rect 1393 18803 1459 18806
rect 2129 18866 2195 18869
rect 18689 18866 18755 18869
rect 2129 18864 18755 18866
rect 2129 18808 2134 18864
rect 2190 18808 18694 18864
rect 18750 18808 18755 18864
rect 2129 18806 18755 18808
rect 2129 18803 2195 18806
rect 18689 18803 18755 18806
rect 21541 18866 21607 18869
rect 22200 18866 23000 18896
rect 21541 18864 23000 18866
rect 21541 18808 21546 18864
rect 21602 18808 23000 18864
rect 21541 18806 23000 18808
rect 21541 18803 21607 18806
rect 22200 18776 23000 18806
rect 2589 18730 2655 18733
rect 18689 18730 18755 18733
rect 2589 18728 18755 18730
rect 2589 18672 2594 18728
rect 2650 18672 18694 18728
rect 18750 18672 18755 18728
rect 2589 18670 18755 18672
rect 2589 18667 2655 18670
rect 18689 18667 18755 18670
rect 2497 18594 2563 18597
rect 3877 18594 3943 18597
rect 2497 18592 3943 18594
rect 2497 18536 2502 18592
rect 2558 18536 3882 18592
rect 3938 18536 3943 18592
rect 2497 18534 3943 18536
rect 2497 18531 2563 18534
rect 3877 18531 3943 18534
rect 5441 18594 5507 18597
rect 8845 18594 8911 18597
rect 9213 18594 9279 18597
rect 5441 18592 9279 18594
rect 5441 18536 5446 18592
rect 5502 18536 8850 18592
rect 8906 18536 9218 18592
rect 9274 18536 9279 18592
rect 5441 18534 9279 18536
rect 5441 18531 5507 18534
rect 8845 18531 8911 18534
rect 9213 18531 9279 18534
rect 4409 18528 4729 18529
rect 0 18458 800 18488
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 1853 18458 1919 18461
rect 0 18456 1919 18458
rect 0 18400 1858 18456
rect 1914 18400 1919 18456
rect 0 18398 1919 18400
rect 0 18368 800 18398
rect 1853 18395 1919 18398
rect 6269 18458 6335 18461
rect 6821 18458 6887 18461
rect 6269 18456 6887 18458
rect 6269 18400 6274 18456
rect 6330 18400 6826 18456
rect 6882 18400 6887 18456
rect 6269 18398 6887 18400
rect 6269 18395 6335 18398
rect 6821 18395 6887 18398
rect 21173 18458 21239 18461
rect 22200 18458 23000 18488
rect 21173 18456 23000 18458
rect 21173 18400 21178 18456
rect 21234 18400 23000 18456
rect 21173 18398 23000 18400
rect 21173 18395 21239 18398
rect 22200 18368 23000 18398
rect 2037 18322 2103 18325
rect 18045 18322 18111 18325
rect 2037 18320 18111 18322
rect 2037 18264 2042 18320
rect 2098 18264 18050 18320
rect 18106 18264 18111 18320
rect 2037 18262 18111 18264
rect 2037 18259 2103 18262
rect 18045 18259 18111 18262
rect 3969 18186 4035 18189
rect 9581 18186 9647 18189
rect 3969 18184 9647 18186
rect 3969 18128 3974 18184
rect 4030 18128 9586 18184
rect 9642 18128 9647 18184
rect 3969 18126 9647 18128
rect 3969 18123 4035 18126
rect 9581 18123 9647 18126
rect 0 18050 800 18080
rect 1485 18050 1551 18053
rect 0 18048 1551 18050
rect 0 17992 1490 18048
rect 1546 17992 1551 18048
rect 0 17990 1551 17992
rect 0 17960 800 17990
rect 1485 17987 1551 17990
rect 21541 18050 21607 18053
rect 22200 18050 23000 18080
rect 21541 18048 23000 18050
rect 21541 17992 21546 18048
rect 21602 17992 23000 18048
rect 21541 17990 23000 17992
rect 21541 17987 21607 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22200 17960 23000 17990
rect 14805 17919 15125 17920
rect 2405 17914 2471 17917
rect 4521 17914 4587 17917
rect 5441 17914 5507 17917
rect 2405 17912 5507 17914
rect 2405 17856 2410 17912
rect 2466 17856 4526 17912
rect 4582 17856 5446 17912
rect 5502 17856 5507 17912
rect 2405 17854 5507 17856
rect 2405 17851 2471 17854
rect 4521 17851 4587 17854
rect 5441 17851 5507 17854
rect 7557 17778 7623 17781
rect 10542 17778 10548 17780
rect 7557 17776 10548 17778
rect 7557 17720 7562 17776
rect 7618 17720 10548 17776
rect 7557 17718 10548 17720
rect 7557 17715 7623 17718
rect 10542 17716 10548 17718
rect 10612 17716 10618 17780
rect 0 17642 800 17672
rect 1761 17642 1827 17645
rect 0 17640 1827 17642
rect 0 17584 1766 17640
rect 1822 17584 1827 17640
rect 0 17582 1827 17584
rect 0 17552 800 17582
rect 1761 17579 1827 17582
rect 2957 17642 3023 17645
rect 7741 17642 7807 17645
rect 11053 17642 11119 17645
rect 11329 17642 11395 17645
rect 2957 17640 8310 17642
rect 2957 17584 2962 17640
rect 3018 17584 7746 17640
rect 7802 17584 8310 17640
rect 2957 17582 8310 17584
rect 2957 17579 3023 17582
rect 7741 17579 7807 17582
rect 8250 17506 8310 17582
rect 11053 17640 11395 17642
rect 11053 17584 11058 17640
rect 11114 17584 11334 17640
rect 11390 17584 11395 17640
rect 11053 17582 11395 17584
rect 11053 17579 11119 17582
rect 11329 17579 11395 17582
rect 21541 17642 21607 17645
rect 22200 17642 23000 17672
rect 21541 17640 23000 17642
rect 21541 17584 21546 17640
rect 21602 17584 23000 17640
rect 21541 17582 23000 17584
rect 21541 17579 21607 17582
rect 22200 17552 23000 17582
rect 8569 17508 8635 17509
rect 8518 17506 8524 17508
rect 8250 17446 8524 17506
rect 8588 17506 8635 17508
rect 9857 17506 9923 17509
rect 9990 17506 9996 17508
rect 8588 17504 8680 17506
rect 8630 17448 8680 17504
rect 8518 17444 8524 17446
rect 8588 17446 8680 17448
rect 9857 17504 9996 17506
rect 9857 17448 9862 17504
rect 9918 17448 9996 17504
rect 9857 17446 9996 17448
rect 8588 17444 8635 17446
rect 8569 17443 8635 17444
rect 9857 17443 9923 17446
rect 9990 17444 9996 17446
rect 10060 17444 10066 17508
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 6862 17172 6868 17236
rect 6932 17234 6938 17236
rect 8201 17234 8267 17237
rect 6932 17232 8267 17234
rect 6932 17176 8206 17232
rect 8262 17176 8267 17232
rect 6932 17174 8267 17176
rect 6932 17172 6938 17174
rect 8201 17171 8267 17174
rect 9765 17234 9831 17237
rect 15469 17234 15535 17237
rect 9765 17232 15535 17234
rect 9765 17176 9770 17232
rect 9826 17176 15474 17232
rect 15530 17176 15535 17232
rect 9765 17174 15535 17176
rect 9765 17171 9831 17174
rect 15469 17171 15535 17174
rect 21541 17234 21607 17237
rect 22200 17234 23000 17264
rect 21541 17232 23000 17234
rect 21541 17176 21546 17232
rect 21602 17176 23000 17232
rect 21541 17174 23000 17176
rect 21541 17171 21607 17174
rect 22200 17144 23000 17174
rect 5942 16900 5948 16964
rect 6012 16962 6018 16964
rect 7281 16962 7347 16965
rect 6012 16960 7347 16962
rect 6012 16904 7286 16960
rect 7342 16904 7347 16960
rect 6012 16902 7347 16904
rect 6012 16900 6018 16902
rect 7281 16899 7347 16902
rect 7874 16896 8194 16897
rect 0 16826 800 16856
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 1485 16826 1551 16829
rect 0 16824 1551 16826
rect 0 16768 1490 16824
rect 1546 16768 1551 16824
rect 0 16766 1551 16768
rect 0 16736 800 16766
rect 1485 16763 1551 16766
rect 12566 16764 12572 16828
rect 12636 16826 12642 16828
rect 13813 16826 13879 16829
rect 12636 16824 13879 16826
rect 12636 16768 13818 16824
rect 13874 16768 13879 16824
rect 12636 16766 13879 16768
rect 12636 16764 12642 16766
rect 13813 16763 13879 16766
rect 21541 16826 21607 16829
rect 22200 16826 23000 16856
rect 21541 16824 23000 16826
rect 21541 16768 21546 16824
rect 21602 16768 23000 16824
rect 21541 16766 23000 16768
rect 21541 16763 21607 16766
rect 22200 16736 23000 16766
rect 10409 16690 10475 16693
rect 11053 16690 11119 16693
rect 10409 16688 11119 16690
rect 10409 16632 10414 16688
rect 10470 16632 11058 16688
rect 11114 16632 11119 16688
rect 10409 16630 11119 16632
rect 10409 16627 10475 16630
rect 11053 16627 11119 16630
rect 3877 16554 3943 16557
rect 8569 16554 8635 16557
rect 3877 16552 8635 16554
rect 3877 16496 3882 16552
rect 3938 16496 8574 16552
rect 8630 16496 8635 16552
rect 3877 16494 8635 16496
rect 3877 16491 3943 16494
rect 8569 16491 8635 16494
rect 9857 16554 9923 16557
rect 11145 16554 11211 16557
rect 9857 16552 11211 16554
rect 9857 16496 9862 16552
rect 9918 16496 11150 16552
rect 11206 16496 11211 16552
rect 9857 16494 11211 16496
rect 9857 16491 9923 16494
rect 11145 16491 11211 16494
rect 4409 16352 4729 16353
rect 0 16282 800 16312
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 1485 16282 1551 16285
rect 0 16280 1551 16282
rect 0 16224 1490 16280
rect 1546 16224 1551 16280
rect 0 16222 1551 16224
rect 0 16192 800 16222
rect 1485 16219 1551 16222
rect 21541 16282 21607 16285
rect 22200 16282 23000 16312
rect 21541 16280 23000 16282
rect 21541 16224 21546 16280
rect 21602 16224 23000 16280
rect 21541 16222 23000 16224
rect 21541 16219 21607 16222
rect 22200 16192 23000 16222
rect 8477 16146 8543 16149
rect 8702 16146 8708 16148
rect 8477 16144 8708 16146
rect 8477 16088 8482 16144
rect 8538 16088 8708 16144
rect 8477 16086 8708 16088
rect 8477 16083 8543 16086
rect 8702 16084 8708 16086
rect 8772 16084 8778 16148
rect 0 15874 800 15904
rect 1853 15874 1919 15877
rect 0 15872 1919 15874
rect 0 15816 1858 15872
rect 1914 15816 1919 15872
rect 0 15814 1919 15816
rect 0 15784 800 15814
rect 1853 15811 1919 15814
rect 8937 15874 9003 15877
rect 9254 15874 9260 15876
rect 8937 15872 9260 15874
rect 8937 15816 8942 15872
rect 8998 15816 9260 15872
rect 8937 15814 9260 15816
rect 8937 15811 9003 15814
rect 9254 15812 9260 15814
rect 9324 15812 9330 15876
rect 21173 15874 21239 15877
rect 22200 15874 23000 15904
rect 21173 15872 23000 15874
rect 21173 15816 21178 15872
rect 21234 15816 23000 15872
rect 21173 15814 23000 15816
rect 21173 15811 21239 15814
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 22200 15784 23000 15814
rect 14805 15743 15125 15744
rect 0 15466 800 15496
rect 1393 15466 1459 15469
rect 0 15464 1459 15466
rect 0 15408 1398 15464
rect 1454 15408 1459 15464
rect 0 15406 1459 15408
rect 0 15376 800 15406
rect 1393 15403 1459 15406
rect 11973 15466 12039 15469
rect 13445 15466 13511 15469
rect 11973 15464 13511 15466
rect 11973 15408 11978 15464
rect 12034 15408 13450 15464
rect 13506 15408 13511 15464
rect 11973 15406 13511 15408
rect 11973 15403 12039 15406
rect 13445 15403 13511 15406
rect 21541 15466 21607 15469
rect 22200 15466 23000 15496
rect 21541 15464 23000 15466
rect 21541 15408 21546 15464
rect 21602 15408 23000 15464
rect 21541 15406 23000 15408
rect 21541 15403 21607 15406
rect 22200 15376 23000 15406
rect 11881 15332 11947 15333
rect 11830 15268 11836 15332
rect 11900 15330 11947 15332
rect 11900 15328 11992 15330
rect 11942 15272 11992 15328
rect 11900 15270 11992 15272
rect 11900 15268 11947 15270
rect 11881 15267 11947 15268
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 11973 15196 12039 15197
rect 11973 15194 12020 15196
rect 11928 15192 12020 15194
rect 11928 15136 11978 15192
rect 11928 15134 12020 15136
rect 11973 15132 12020 15134
rect 12084 15132 12090 15196
rect 12341 15194 12407 15197
rect 16573 15194 16639 15197
rect 12341 15192 16639 15194
rect 12341 15136 12346 15192
rect 12402 15136 16578 15192
rect 16634 15136 16639 15192
rect 12341 15134 16639 15136
rect 11973 15131 12039 15132
rect 12341 15131 12407 15134
rect 16573 15131 16639 15134
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 21541 15058 21607 15061
rect 22200 15058 23000 15088
rect 21541 15056 23000 15058
rect 21541 15000 21546 15056
rect 21602 15000 23000 15056
rect 21541 14998 23000 15000
rect 21541 14995 21607 14998
rect 22200 14968 23000 14998
rect 7833 14922 7899 14925
rect 9581 14922 9647 14925
rect 7833 14920 9647 14922
rect 7833 14864 7838 14920
rect 7894 14864 9586 14920
rect 9642 14864 9647 14920
rect 7833 14862 9647 14864
rect 7833 14859 7899 14862
rect 9581 14859 9647 14862
rect 10174 14724 10180 14788
rect 10244 14786 10250 14788
rect 10317 14786 10383 14789
rect 10244 14784 10383 14786
rect 10244 14728 10322 14784
rect 10378 14728 10383 14784
rect 10244 14726 10383 14728
rect 10244 14724 10250 14726
rect 10317 14723 10383 14726
rect 12157 14786 12223 14789
rect 14641 14786 14707 14789
rect 12157 14784 14707 14786
rect 12157 14728 12162 14784
rect 12218 14728 14646 14784
rect 14702 14728 14707 14784
rect 12157 14726 14707 14728
rect 12157 14723 12223 14726
rect 14641 14723 14707 14726
rect 7874 14720 8194 14721
rect 0 14650 800 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 1853 14650 1919 14653
rect 0 14648 1919 14650
rect 0 14592 1858 14648
rect 1914 14592 1919 14648
rect 0 14590 1919 14592
rect 0 14560 800 14590
rect 1853 14587 1919 14590
rect 6177 14650 6243 14653
rect 7557 14650 7623 14653
rect 6177 14648 7623 14650
rect 6177 14592 6182 14648
rect 6238 14592 7562 14648
rect 7618 14592 7623 14648
rect 6177 14590 7623 14592
rect 6177 14587 6243 14590
rect 7557 14587 7623 14590
rect 21173 14650 21239 14653
rect 22200 14650 23000 14680
rect 21173 14648 23000 14650
rect 21173 14592 21178 14648
rect 21234 14592 23000 14648
rect 21173 14590 23000 14592
rect 21173 14587 21239 14590
rect 22200 14560 23000 14590
rect 6678 14452 6684 14516
rect 6748 14514 6754 14516
rect 11421 14514 11487 14517
rect 6748 14512 11487 14514
rect 6748 14456 11426 14512
rect 11482 14456 11487 14512
rect 6748 14454 11487 14456
rect 6748 14452 6754 14454
rect 11421 14451 11487 14454
rect 3969 14378 4035 14381
rect 10961 14378 11027 14381
rect 3969 14376 11027 14378
rect 3969 14320 3974 14376
rect 4030 14320 10966 14376
rect 11022 14320 11027 14376
rect 3969 14318 11027 14320
rect 3969 14315 4035 14318
rect 10961 14315 11027 14318
rect 12341 14378 12407 14381
rect 18781 14378 18847 14381
rect 12341 14376 18847 14378
rect 12341 14320 12346 14376
rect 12402 14320 18786 14376
rect 18842 14320 18847 14376
rect 12341 14318 18847 14320
rect 12341 14315 12407 14318
rect 18781 14315 18847 14318
rect 0 14242 800 14272
rect 1485 14242 1551 14245
rect 0 14240 1551 14242
rect 0 14184 1490 14240
rect 1546 14184 1551 14240
rect 0 14182 1551 14184
rect 0 14152 800 14182
rect 1485 14179 1551 14182
rect 4838 14180 4844 14244
rect 4908 14242 4914 14244
rect 4981 14242 5047 14245
rect 4908 14240 5047 14242
rect 4908 14184 4986 14240
rect 5042 14184 5047 14240
rect 4908 14182 5047 14184
rect 4908 14180 4914 14182
rect 4981 14179 5047 14182
rect 5165 14242 5231 14245
rect 8886 14242 8892 14244
rect 5165 14240 8892 14242
rect 5165 14184 5170 14240
rect 5226 14184 8892 14240
rect 5165 14182 8892 14184
rect 5165 14179 5231 14182
rect 8886 14180 8892 14182
rect 8956 14180 8962 14244
rect 13721 14242 13787 14245
rect 17401 14242 17467 14245
rect 13721 14240 17467 14242
rect 13721 14184 13726 14240
rect 13782 14184 17406 14240
rect 17462 14184 17467 14240
rect 13721 14182 17467 14184
rect 13721 14179 13787 14182
rect 17401 14179 17467 14182
rect 21541 14242 21607 14245
rect 22200 14242 23000 14272
rect 21541 14240 23000 14242
rect 21541 14184 21546 14240
rect 21602 14184 23000 14240
rect 21541 14182 23000 14184
rect 21541 14179 21607 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 22200 14152 23000 14182
rect 18270 14111 18590 14112
rect 9213 14106 9279 14109
rect 10409 14106 10475 14109
rect 10777 14106 10843 14109
rect 9213 14104 9322 14106
rect 9213 14048 9218 14104
rect 9274 14048 9322 14104
rect 9213 14043 9322 14048
rect 10409 14104 10843 14106
rect 10409 14048 10414 14104
rect 10470 14048 10782 14104
rect 10838 14048 10843 14104
rect 10409 14046 10843 14048
rect 10409 14043 10475 14046
rect 10777 14043 10843 14046
rect 12382 14044 12388 14108
rect 12452 14106 12458 14108
rect 12801 14106 12867 14109
rect 16665 14106 16731 14109
rect 12452 14104 12867 14106
rect 12452 14048 12806 14104
rect 12862 14048 12867 14104
rect 12452 14046 12867 14048
rect 12452 14044 12458 14046
rect 12801 14043 12867 14046
rect 14414 14104 16731 14106
rect 14414 14048 16670 14104
rect 16726 14048 16731 14104
rect 14414 14046 16731 14048
rect 5942 13908 5948 13972
rect 6012 13970 6018 13972
rect 8845 13970 8911 13973
rect 6012 13968 8911 13970
rect 6012 13912 8850 13968
rect 8906 13912 8911 13968
rect 6012 13910 8911 13912
rect 6012 13908 6018 13910
rect 8845 13907 8911 13910
rect 0 13834 800 13864
rect 1761 13834 1827 13837
rect 0 13832 1827 13834
rect 0 13776 1766 13832
rect 1822 13776 1827 13832
rect 0 13774 1827 13776
rect 0 13744 800 13774
rect 1761 13771 1827 13774
rect 4705 13834 4771 13837
rect 5257 13834 5323 13837
rect 6177 13834 6243 13837
rect 4705 13832 6243 13834
rect 4705 13776 4710 13832
rect 4766 13776 5262 13832
rect 5318 13776 6182 13832
rect 6238 13776 6243 13832
rect 4705 13774 6243 13776
rect 4705 13771 4771 13774
rect 5257 13771 5323 13774
rect 6177 13771 6243 13774
rect 3969 13698 4035 13701
rect 4153 13698 4219 13701
rect 5349 13698 5415 13701
rect 6821 13698 6887 13701
rect 3969 13696 6887 13698
rect 3969 13640 3974 13696
rect 4030 13640 4158 13696
rect 4214 13640 5354 13696
rect 5410 13640 6826 13696
rect 6882 13640 6887 13696
rect 3969 13638 6887 13640
rect 3969 13635 4035 13638
rect 4153 13635 4219 13638
rect 5349 13635 5415 13638
rect 6821 13635 6887 13638
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 3325 13562 3391 13565
rect 5533 13562 5599 13565
rect 3325 13560 5599 13562
rect 3325 13504 3330 13560
rect 3386 13504 5538 13560
rect 5594 13504 5599 13560
rect 3325 13502 5599 13504
rect 3325 13499 3391 13502
rect 5533 13499 5599 13502
rect 5717 13562 5783 13565
rect 6913 13562 6979 13565
rect 5717 13560 6979 13562
rect 5717 13504 5722 13560
rect 5778 13504 6918 13560
rect 6974 13504 6979 13560
rect 5717 13502 6979 13504
rect 5717 13499 5783 13502
rect 6913 13499 6979 13502
rect 0 13426 800 13456
rect 1393 13426 1459 13429
rect 5901 13428 5967 13429
rect 5901 13426 5948 13428
rect 0 13424 1459 13426
rect 0 13368 1398 13424
rect 1454 13368 1459 13424
rect 0 13366 1459 13368
rect 5856 13424 5948 13426
rect 5856 13368 5906 13424
rect 5856 13366 5948 13368
rect 0 13336 800 13366
rect 1393 13363 1459 13366
rect 5901 13364 5948 13366
rect 6012 13364 6018 13428
rect 7557 13426 7623 13429
rect 9262 13426 9322 14043
rect 10542 13908 10548 13972
rect 10612 13970 10618 13972
rect 14414 13970 14474 14046
rect 16665 14043 16731 14046
rect 10612 13910 14474 13970
rect 14549 13970 14615 13973
rect 16021 13970 16087 13973
rect 14549 13968 16087 13970
rect 14549 13912 14554 13968
rect 14610 13912 16026 13968
rect 16082 13912 16087 13968
rect 14549 13910 16087 13912
rect 10612 13908 10618 13910
rect 14549 13907 14615 13910
rect 16021 13907 16087 13910
rect 10133 13832 10199 13837
rect 10133 13776 10138 13832
rect 10194 13776 10199 13832
rect 10133 13771 10199 13776
rect 10501 13834 10567 13837
rect 15653 13834 15719 13837
rect 10501 13832 15719 13834
rect 10501 13776 10506 13832
rect 10562 13776 15658 13832
rect 15714 13776 15719 13832
rect 10501 13774 15719 13776
rect 10501 13771 10567 13774
rect 15653 13771 15719 13774
rect 21541 13834 21607 13837
rect 22200 13834 23000 13864
rect 21541 13832 23000 13834
rect 21541 13776 21546 13832
rect 21602 13776 23000 13832
rect 21541 13774 23000 13776
rect 21541 13771 21607 13774
rect 9857 13700 9923 13701
rect 9806 13636 9812 13700
rect 9876 13698 9923 13700
rect 9876 13696 9968 13698
rect 9918 13640 9968 13696
rect 9876 13638 9968 13640
rect 9876 13636 9923 13638
rect 9857 13635 9923 13636
rect 10136 13562 10196 13771
rect 22200 13744 23000 13774
rect 11329 13698 11395 13701
rect 14590 13698 14596 13700
rect 11329 13696 14596 13698
rect 11329 13640 11334 13696
rect 11390 13640 14596 13696
rect 11329 13638 14596 13640
rect 11329 13635 11395 13638
rect 14590 13636 14596 13638
rect 14660 13636 14666 13700
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 10593 13562 10659 13565
rect 10136 13560 10659 13562
rect 10136 13504 10598 13560
rect 10654 13504 10659 13560
rect 10136 13502 10659 13504
rect 10593 13499 10659 13502
rect 10869 13562 10935 13565
rect 11421 13562 11487 13565
rect 10869 13560 11487 13562
rect 10869 13504 10874 13560
rect 10930 13504 11426 13560
rect 11482 13504 11487 13560
rect 10869 13502 11487 13504
rect 10869 13499 10935 13502
rect 11421 13499 11487 13502
rect 15009 13426 15075 13429
rect 7557 13424 15075 13426
rect 7557 13368 7562 13424
rect 7618 13368 15014 13424
rect 15070 13368 15075 13424
rect 7557 13366 15075 13368
rect 5901 13363 5967 13364
rect 7557 13363 7623 13366
rect 15009 13363 15075 13366
rect 21541 13426 21607 13429
rect 22200 13426 23000 13456
rect 21541 13424 23000 13426
rect 21541 13368 21546 13424
rect 21602 13368 23000 13424
rect 21541 13366 23000 13368
rect 21541 13363 21607 13366
rect 22200 13336 23000 13366
rect 11421 13290 11487 13293
rect 16113 13290 16179 13293
rect 8158 13288 16179 13290
rect 8158 13232 11426 13288
rect 11482 13232 16118 13288
rect 16174 13232 16179 13288
rect 8158 13230 16179 13232
rect 5809 13154 5875 13157
rect 8158 13154 8218 13230
rect 11421 13227 11487 13230
rect 16113 13227 16179 13230
rect 5809 13152 8218 13154
rect 5809 13096 5814 13152
rect 5870 13096 8218 13152
rect 5809 13094 8218 13096
rect 14089 13154 14155 13157
rect 14222 13154 14228 13156
rect 14089 13152 14228 13154
rect 14089 13096 14094 13152
rect 14150 13096 14228 13152
rect 14089 13094 14228 13096
rect 5809 13091 5875 13094
rect 14089 13091 14155 13094
rect 14222 13092 14228 13094
rect 14292 13154 14298 13156
rect 14825 13154 14891 13157
rect 14292 13152 14891 13154
rect 14292 13096 14830 13152
rect 14886 13096 14891 13152
rect 14292 13094 14891 13096
rect 14292 13092 14298 13094
rect 14825 13091 14891 13094
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 5349 13018 5415 13021
rect 8569 13018 8635 13021
rect 9121 13020 9187 13021
rect 9070 13018 9076 13020
rect 5349 13016 8635 13018
rect 5349 12960 5354 13016
rect 5410 12960 8574 13016
rect 8630 12960 8635 13016
rect 5349 12958 8635 12960
rect 9030 12958 9076 13018
rect 9140 13016 9187 13020
rect 9182 12960 9187 13016
rect 5349 12955 5415 12958
rect 8569 12955 8635 12958
rect 9070 12956 9076 12958
rect 9140 12956 9187 12960
rect 9121 12955 9187 12956
rect 9305 13018 9371 13021
rect 11053 13018 11119 13021
rect 9305 13016 11119 13018
rect 9305 12960 9310 13016
rect 9366 12960 11058 13016
rect 11114 12960 11119 13016
rect 9305 12958 11119 12960
rect 9305 12955 9371 12958
rect 11053 12955 11119 12958
rect 14825 13018 14891 13021
rect 15285 13018 15351 13021
rect 16389 13018 16455 13021
rect 14825 13016 16455 13018
rect 14825 12960 14830 13016
rect 14886 12960 15290 13016
rect 15346 12960 16394 13016
rect 16450 12960 16455 13016
rect 14825 12958 16455 12960
rect 14825 12955 14891 12958
rect 15285 12955 15351 12958
rect 16389 12955 16455 12958
rect 0 12882 800 12912
rect 1853 12882 1919 12885
rect 0 12880 1919 12882
rect 0 12824 1858 12880
rect 1914 12824 1919 12880
rect 0 12822 1919 12824
rect 0 12792 800 12822
rect 1853 12819 1919 12822
rect 7557 12882 7623 12885
rect 10225 12882 10291 12885
rect 7557 12880 10291 12882
rect 7557 12824 7562 12880
rect 7618 12824 10230 12880
rect 10286 12824 10291 12880
rect 7557 12822 10291 12824
rect 7557 12819 7623 12822
rect 10225 12819 10291 12822
rect 10501 12882 10567 12885
rect 10961 12884 11027 12885
rect 10501 12880 10610 12882
rect 10501 12824 10506 12880
rect 10562 12824 10610 12880
rect 10501 12819 10610 12824
rect 10910 12820 10916 12884
rect 10980 12882 11027 12884
rect 13353 12882 13419 12885
rect 17953 12882 18019 12885
rect 10980 12880 11072 12882
rect 11022 12824 11072 12880
rect 10980 12822 11072 12824
rect 13353 12880 18019 12882
rect 13353 12824 13358 12880
rect 13414 12824 17958 12880
rect 18014 12824 18019 12880
rect 13353 12822 18019 12824
rect 10980 12820 11027 12822
rect 10961 12819 11027 12820
rect 13353 12819 13419 12822
rect 17953 12819 18019 12822
rect 21541 12882 21607 12885
rect 22200 12882 23000 12912
rect 21541 12880 23000 12882
rect 21541 12824 21546 12880
rect 21602 12824 23000 12880
rect 21541 12822 23000 12824
rect 21541 12819 21607 12822
rect 3601 12746 3667 12749
rect 6637 12748 6703 12749
rect 6637 12746 6684 12748
rect 3601 12744 6684 12746
rect 6748 12746 6754 12748
rect 8201 12746 8267 12749
rect 8334 12746 8340 12748
rect 3601 12688 3606 12744
rect 3662 12688 6642 12744
rect 3601 12686 6684 12688
rect 3601 12683 3667 12686
rect 6637 12684 6684 12686
rect 6748 12686 6830 12746
rect 8201 12744 8340 12746
rect 8201 12688 8206 12744
rect 8262 12688 8340 12744
rect 8201 12686 8340 12688
rect 6748 12684 6754 12686
rect 6637 12683 6703 12684
rect 8201 12683 8267 12686
rect 8334 12684 8340 12686
rect 8404 12684 8410 12748
rect 8661 12746 8727 12749
rect 10358 12746 10364 12748
rect 8661 12744 10364 12746
rect 8661 12688 8666 12744
rect 8722 12688 10364 12744
rect 8661 12686 10364 12688
rect 8661 12683 8727 12686
rect 10358 12684 10364 12686
rect 10428 12684 10434 12748
rect 3877 12610 3943 12613
rect 7005 12610 7071 12613
rect 3877 12608 7071 12610
rect 3877 12552 3882 12608
rect 3938 12552 7010 12608
rect 7066 12552 7071 12608
rect 3877 12550 7071 12552
rect 3877 12547 3943 12550
rect 7005 12547 7071 12550
rect 8753 12610 8819 12613
rect 9213 12610 9279 12613
rect 8753 12608 9279 12610
rect 8753 12552 8758 12608
rect 8814 12552 9218 12608
rect 9274 12552 9279 12608
rect 8753 12550 9279 12552
rect 8753 12547 8819 12550
rect 9213 12547 9279 12550
rect 9438 12548 9444 12612
rect 9508 12610 9514 12612
rect 10133 12610 10199 12613
rect 10550 12610 10610 12819
rect 22200 12792 23000 12822
rect 9508 12608 10610 12610
rect 9508 12552 10138 12608
rect 10194 12552 10610 12608
rect 9508 12550 10610 12552
rect 10961 12610 11027 12613
rect 10961 12608 11530 12610
rect 10961 12552 10966 12608
rect 11022 12552 11530 12608
rect 10961 12550 11530 12552
rect 9508 12548 9514 12550
rect 10133 12547 10199 12550
rect 10961 12547 11027 12550
rect 7874 12544 8194 12545
rect 0 12474 800 12504
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 1393 12474 1459 12477
rect 0 12472 1459 12474
rect 0 12416 1398 12472
rect 1454 12416 1459 12472
rect 0 12414 1459 12416
rect 0 12384 800 12414
rect 1393 12411 1459 12414
rect 6545 12474 6611 12477
rect 6678 12474 6684 12476
rect 6545 12472 6684 12474
rect 6545 12416 6550 12472
rect 6606 12416 6684 12472
rect 6545 12414 6684 12416
rect 6545 12411 6611 12414
rect 6678 12412 6684 12414
rect 6748 12412 6754 12476
rect 8845 12474 8911 12477
rect 8296 12472 8911 12474
rect 8296 12416 8850 12472
rect 8906 12416 8911 12472
rect 8296 12414 8911 12416
rect 5533 12340 5599 12341
rect 5533 12338 5580 12340
rect 5488 12336 5580 12338
rect 5488 12280 5538 12336
rect 5488 12278 5580 12280
rect 5533 12276 5580 12278
rect 5644 12276 5650 12340
rect 5758 12276 5764 12340
rect 5828 12338 5834 12340
rect 5901 12338 5967 12341
rect 6729 12340 6795 12341
rect 6678 12338 6684 12340
rect 5828 12336 5967 12338
rect 5828 12280 5906 12336
rect 5962 12280 5967 12336
rect 5828 12278 5967 12280
rect 6638 12278 6684 12338
rect 6748 12336 6795 12340
rect 6790 12280 6795 12336
rect 5828 12276 5834 12278
rect 5533 12275 5599 12276
rect 5901 12275 5967 12278
rect 6678 12276 6684 12278
rect 6748 12276 6795 12280
rect 6729 12275 6795 12276
rect 8109 12338 8175 12341
rect 8296 12338 8356 12414
rect 8845 12411 8911 12414
rect 9121 12474 9187 12477
rect 9397 12474 9463 12477
rect 9121 12472 9463 12474
rect 9121 12416 9126 12472
rect 9182 12416 9402 12472
rect 9458 12416 9463 12472
rect 9121 12414 9463 12416
rect 9121 12411 9187 12414
rect 9397 12411 9463 12414
rect 9765 12474 9831 12477
rect 10961 12474 11027 12477
rect 9765 12472 11027 12474
rect 9765 12416 9770 12472
rect 9826 12416 10966 12472
rect 11022 12416 11027 12472
rect 9765 12414 11027 12416
rect 11470 12474 11530 12550
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 11605 12474 11671 12477
rect 13445 12474 13511 12477
rect 11470 12472 11671 12474
rect 11470 12416 11610 12472
rect 11666 12416 11671 12472
rect 11470 12414 11671 12416
rect 9765 12411 9831 12414
rect 10961 12411 11027 12414
rect 11605 12411 11671 12414
rect 12252 12472 13511 12474
rect 12252 12416 13450 12472
rect 13506 12416 13511 12472
rect 12252 12414 13511 12416
rect 8109 12336 8356 12338
rect 8109 12280 8114 12336
rect 8170 12280 8356 12336
rect 8109 12278 8356 12280
rect 8477 12338 8543 12341
rect 9070 12338 9076 12340
rect 8477 12336 9076 12338
rect 8477 12280 8482 12336
rect 8538 12280 9076 12336
rect 8477 12278 9076 12280
rect 8109 12275 8175 12278
rect 8477 12275 8543 12278
rect 9070 12276 9076 12278
rect 9140 12276 9146 12340
rect 9806 12276 9812 12340
rect 9876 12338 9882 12340
rect 12252 12338 12312 12414
rect 13445 12411 13511 12414
rect 21173 12474 21239 12477
rect 22200 12474 23000 12504
rect 21173 12472 23000 12474
rect 21173 12416 21178 12472
rect 21234 12416 23000 12472
rect 21173 12414 23000 12416
rect 21173 12411 21239 12414
rect 22200 12384 23000 12414
rect 9876 12278 12312 12338
rect 9876 12276 9882 12278
rect 12382 12276 12388 12340
rect 12452 12338 12458 12340
rect 18505 12338 18571 12341
rect 12452 12336 18571 12338
rect 12452 12280 18510 12336
rect 18566 12280 18571 12336
rect 12452 12278 18571 12280
rect 12452 12276 12458 12278
rect 18505 12275 18571 12278
rect 5349 12202 5415 12205
rect 12750 12202 12756 12204
rect 5349 12200 12756 12202
rect 5349 12144 5354 12200
rect 5410 12144 12756 12200
rect 5349 12142 12756 12144
rect 5349 12139 5415 12142
rect 12750 12140 12756 12142
rect 12820 12140 12826 12204
rect 0 12066 800 12096
rect 1485 12066 1551 12069
rect 0 12064 1551 12066
rect 0 12008 1490 12064
rect 1546 12008 1551 12064
rect 0 12006 1551 12008
rect 0 11976 800 12006
rect 1485 12003 1551 12006
rect 7373 12066 7439 12069
rect 8385 12066 8451 12069
rect 7373 12064 8451 12066
rect 7373 12008 7378 12064
rect 7434 12008 8390 12064
rect 8446 12008 8451 12064
rect 7373 12006 8451 12008
rect 7373 12003 7439 12006
rect 8385 12003 8451 12006
rect 8569 12066 8635 12069
rect 9489 12066 9555 12069
rect 10409 12068 10475 12069
rect 10358 12066 10364 12068
rect 8569 12064 9555 12066
rect 8569 12008 8574 12064
rect 8630 12008 9494 12064
rect 9550 12008 9555 12064
rect 8569 12006 9555 12008
rect 10318 12006 10364 12066
rect 10428 12064 10475 12068
rect 10470 12008 10475 12064
rect 8569 12003 8635 12006
rect 9489 12003 9555 12006
rect 10358 12004 10364 12006
rect 10428 12004 10475 12008
rect 10910 12004 10916 12068
rect 10980 12066 10986 12068
rect 11145 12066 11211 12069
rect 10980 12064 11211 12066
rect 10980 12008 11150 12064
rect 11206 12008 11211 12064
rect 10980 12006 11211 12008
rect 12758 12066 12818 12140
rect 16665 12066 16731 12069
rect 17769 12066 17835 12069
rect 12758 12064 17835 12066
rect 12758 12008 16670 12064
rect 16726 12008 17774 12064
rect 17830 12008 17835 12064
rect 12758 12006 17835 12008
rect 10980 12004 10986 12006
rect 10409 12003 10475 12004
rect 11145 12003 11211 12006
rect 16665 12003 16731 12006
rect 17769 12003 17835 12006
rect 21541 12066 21607 12069
rect 22200 12066 23000 12096
rect 21541 12064 23000 12066
rect 21541 12008 21546 12064
rect 21602 12008 23000 12064
rect 21541 12006 23000 12008
rect 21541 12003 21607 12006
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 22200 11976 23000 12006
rect 18270 11935 18590 11936
rect 5257 11930 5323 11933
rect 9029 11930 9095 11933
rect 17585 11930 17651 11933
rect 5257 11928 9095 11930
rect 5257 11872 5262 11928
rect 5318 11872 9034 11928
rect 9090 11872 9095 11928
rect 5257 11870 9095 11872
rect 5257 11867 5323 11870
rect 9029 11867 9095 11870
rect 11976 11928 17651 11930
rect 11976 11872 17590 11928
rect 17646 11872 17651 11928
rect 11976 11870 17651 11872
rect 1577 11794 1643 11797
rect 11789 11794 11855 11797
rect 1577 11792 11855 11794
rect 1577 11736 1582 11792
rect 1638 11736 11794 11792
rect 11850 11736 11855 11792
rect 1577 11734 11855 11736
rect 1577 11731 1643 11734
rect 11789 11731 11855 11734
rect 0 11658 800 11688
rect 4061 11658 4127 11661
rect 0 11656 4127 11658
rect 0 11600 4066 11656
rect 4122 11600 4127 11656
rect 0 11598 4127 11600
rect 0 11568 800 11598
rect 4061 11595 4127 11598
rect 4245 11658 4311 11661
rect 8753 11658 8819 11661
rect 4245 11656 8819 11658
rect 4245 11600 4250 11656
rect 4306 11600 8758 11656
rect 8814 11600 8819 11656
rect 4245 11598 8819 11600
rect 4245 11595 4311 11598
rect 8753 11595 8819 11598
rect 9990 11596 9996 11660
rect 10060 11658 10066 11660
rect 10593 11658 10659 11661
rect 11976 11658 12036 11870
rect 17585 11867 17651 11870
rect 12341 11794 12407 11797
rect 18873 11794 18939 11797
rect 19149 11794 19215 11797
rect 12341 11792 19215 11794
rect 12341 11736 12346 11792
rect 12402 11736 18878 11792
rect 18934 11736 19154 11792
rect 19210 11736 19215 11792
rect 12341 11734 19215 11736
rect 12341 11731 12407 11734
rect 18873 11731 18939 11734
rect 19149 11731 19215 11734
rect 10060 11656 12036 11658
rect 10060 11600 10598 11656
rect 10654 11600 12036 11656
rect 10060 11598 12036 11600
rect 13169 11658 13235 11661
rect 18781 11658 18847 11661
rect 13169 11656 18847 11658
rect 13169 11600 13174 11656
rect 13230 11600 18786 11656
rect 18842 11600 18847 11656
rect 13169 11598 18847 11600
rect 10060 11596 10066 11598
rect 10593 11595 10659 11598
rect 13169 11595 13235 11598
rect 18781 11595 18847 11598
rect 20437 11658 20503 11661
rect 22200 11658 23000 11688
rect 20437 11656 23000 11658
rect 20437 11600 20442 11656
rect 20498 11600 23000 11656
rect 20437 11598 23000 11600
rect 20437 11595 20503 11598
rect 22200 11568 23000 11598
rect 7373 11524 7439 11525
rect 7373 11522 7420 11524
rect 7328 11520 7420 11522
rect 7328 11464 7378 11520
rect 7328 11462 7420 11464
rect 7373 11460 7420 11462
rect 7484 11460 7490 11524
rect 8753 11522 8819 11525
rect 9489 11522 9555 11525
rect 9673 11524 9739 11525
rect 8753 11520 9555 11522
rect 8753 11464 8758 11520
rect 8814 11464 9494 11520
rect 9550 11464 9555 11520
rect 8753 11462 9555 11464
rect 7373 11459 7439 11460
rect 8753 11459 8819 11462
rect 9489 11459 9555 11462
rect 9622 11460 9628 11524
rect 9692 11522 9739 11524
rect 10041 11522 10107 11525
rect 10593 11522 10659 11525
rect 9692 11520 9784 11522
rect 9734 11464 9784 11520
rect 9692 11462 9784 11464
rect 10041 11520 10659 11522
rect 10041 11464 10046 11520
rect 10102 11464 10598 11520
rect 10654 11464 10659 11520
rect 10041 11462 10659 11464
rect 9692 11460 9739 11462
rect 9673 11459 9739 11460
rect 10041 11459 10107 11462
rect 10593 11459 10659 11462
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 9857 11386 9923 11389
rect 10501 11386 10567 11389
rect 9857 11384 10567 11386
rect 9857 11328 9862 11384
rect 9918 11328 10506 11384
rect 10562 11328 10567 11384
rect 9857 11326 10567 11328
rect 9857 11323 9923 11326
rect 10501 11323 10567 11326
rect 0 11250 800 11280
rect 3325 11250 3391 11253
rect 0 11248 3391 11250
rect 0 11192 3330 11248
rect 3386 11192 3391 11248
rect 0 11190 3391 11192
rect 0 11160 800 11190
rect 3325 11187 3391 11190
rect 6085 11250 6151 11253
rect 14825 11250 14891 11253
rect 6085 11248 14891 11250
rect 6085 11192 6090 11248
rect 6146 11192 14830 11248
rect 14886 11192 14891 11248
rect 6085 11190 14891 11192
rect 6085 11187 6151 11190
rect 14825 11187 14891 11190
rect 21541 11250 21607 11253
rect 22200 11250 23000 11280
rect 21541 11248 23000 11250
rect 21541 11192 21546 11248
rect 21602 11192 23000 11248
rect 21541 11190 23000 11192
rect 21541 11187 21607 11190
rect 22200 11160 23000 11190
rect 7373 11114 7439 11117
rect 13353 11114 13419 11117
rect 7373 11112 13419 11114
rect 7373 11056 7378 11112
rect 7434 11056 13358 11112
rect 13414 11056 13419 11112
rect 7373 11054 13419 11056
rect 7373 11051 7439 11054
rect 13353 11051 13419 11054
rect 15469 11114 15535 11117
rect 16573 11114 16639 11117
rect 15469 11112 16639 11114
rect 15469 11056 15474 11112
rect 15530 11056 16578 11112
rect 16634 11056 16639 11112
rect 15469 11054 16639 11056
rect 15469 11051 15535 11054
rect 16573 11051 16639 11054
rect 8293 10978 8359 10981
rect 8661 10978 8727 10981
rect 8293 10976 8727 10978
rect 8293 10920 8298 10976
rect 8354 10920 8666 10976
rect 8722 10920 8727 10976
rect 8293 10918 8727 10920
rect 8293 10915 8359 10918
rect 8661 10915 8727 10918
rect 9622 10916 9628 10980
rect 9692 10978 9698 10980
rect 9765 10978 9831 10981
rect 9692 10976 9831 10978
rect 9692 10920 9770 10976
rect 9826 10920 9831 10976
rect 9692 10918 9831 10920
rect 9692 10916 9698 10918
rect 9765 10915 9831 10918
rect 10174 10916 10180 10980
rect 10244 10978 10250 10980
rect 10685 10978 10751 10981
rect 10244 10976 10751 10978
rect 10244 10920 10690 10976
rect 10746 10920 10751 10976
rect 10244 10918 10751 10920
rect 10244 10916 10250 10918
rect 10685 10915 10751 10918
rect 12157 10978 12223 10981
rect 12617 10978 12683 10981
rect 16757 10978 16823 10981
rect 12157 10976 16823 10978
rect 12157 10920 12162 10976
rect 12218 10920 12622 10976
rect 12678 10920 16762 10976
rect 16818 10920 16823 10976
rect 12157 10918 16823 10920
rect 12157 10915 12223 10918
rect 12617 10915 12683 10918
rect 16757 10915 16823 10918
rect 4409 10912 4729 10913
rect 0 10842 800 10872
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 1393 10842 1459 10845
rect 0 10840 1459 10842
rect 0 10784 1398 10840
rect 1454 10784 1459 10840
rect 0 10782 1459 10784
rect 0 10752 800 10782
rect 1393 10779 1459 10782
rect 6678 10780 6684 10844
rect 6748 10842 6754 10844
rect 7741 10842 7807 10845
rect 8845 10842 8911 10845
rect 10593 10842 10659 10845
rect 6748 10840 8310 10842
rect 6748 10784 7746 10840
rect 7802 10784 8310 10840
rect 6748 10782 8310 10784
rect 6748 10780 6754 10782
rect 7741 10779 7807 10782
rect 4245 10706 4311 10709
rect 5625 10708 5691 10709
rect 4838 10706 4844 10708
rect 4245 10704 4844 10706
rect 4245 10648 4250 10704
rect 4306 10648 4844 10704
rect 4245 10646 4844 10648
rect 4245 10643 4311 10646
rect 4838 10644 4844 10646
rect 4908 10644 4914 10708
rect 5574 10706 5580 10708
rect 5498 10646 5580 10706
rect 5644 10706 5691 10708
rect 7046 10706 7052 10708
rect 5644 10704 7052 10706
rect 5686 10648 7052 10704
rect 5574 10644 5580 10646
rect 5644 10646 7052 10648
rect 5644 10644 5691 10646
rect 7046 10644 7052 10646
rect 7116 10706 7122 10708
rect 7557 10706 7623 10709
rect 7116 10704 7623 10706
rect 7116 10648 7562 10704
rect 7618 10648 7623 10704
rect 7116 10646 7623 10648
rect 8250 10706 8310 10782
rect 8845 10840 10659 10842
rect 8845 10784 8850 10840
rect 8906 10784 10598 10840
rect 10654 10784 10659 10840
rect 8845 10782 10659 10784
rect 8845 10779 8911 10782
rect 10593 10779 10659 10782
rect 11973 10842 12039 10845
rect 15285 10842 15351 10845
rect 11973 10840 15351 10842
rect 11973 10784 11978 10840
rect 12034 10784 15290 10840
rect 15346 10784 15351 10840
rect 11973 10782 15351 10784
rect 11973 10779 12039 10782
rect 15285 10779 15351 10782
rect 21449 10842 21515 10845
rect 22200 10842 23000 10872
rect 21449 10840 23000 10842
rect 21449 10784 21454 10840
rect 21510 10784 23000 10840
rect 21449 10782 23000 10784
rect 21449 10779 21515 10782
rect 22200 10752 23000 10782
rect 17309 10706 17375 10709
rect 8250 10704 17375 10706
rect 8250 10648 17314 10704
rect 17370 10648 17375 10704
rect 8250 10646 17375 10648
rect 7116 10644 7122 10646
rect 5625 10643 5691 10644
rect 7557 10643 7623 10646
rect 17309 10643 17375 10646
rect 5533 10570 5599 10573
rect 18045 10570 18111 10573
rect 5533 10568 18111 10570
rect 5533 10512 5538 10568
rect 5594 10512 18050 10568
rect 18106 10512 18111 10568
rect 5533 10510 18111 10512
rect 5533 10507 5599 10510
rect 0 10434 800 10464
rect 1485 10434 1551 10437
rect 0 10432 1551 10434
rect 0 10376 1490 10432
rect 1546 10376 1551 10432
rect 0 10374 1551 10376
rect 0 10344 800 10374
rect 1485 10371 1551 10374
rect 6456 10301 6516 10510
rect 18045 10507 18111 10510
rect 7557 10436 7623 10437
rect 7230 10372 7236 10436
rect 7300 10434 7306 10436
rect 7557 10434 7604 10436
rect 7300 10432 7604 10434
rect 7668 10434 7674 10436
rect 8753 10434 8819 10437
rect 9489 10434 9555 10437
rect 7300 10376 7562 10432
rect 7300 10374 7604 10376
rect 7300 10372 7306 10374
rect 7557 10372 7604 10374
rect 7668 10374 7750 10434
rect 8753 10432 9555 10434
rect 8753 10376 8758 10432
rect 8814 10376 9494 10432
rect 9550 10376 9555 10432
rect 8753 10374 9555 10376
rect 7668 10372 7674 10374
rect 7557 10371 7623 10372
rect 8753 10371 8819 10374
rect 9489 10371 9555 10374
rect 9806 10372 9812 10436
rect 9876 10434 9882 10436
rect 10133 10434 10199 10437
rect 9876 10432 10199 10434
rect 9876 10376 10138 10432
rect 10194 10376 10199 10432
rect 9876 10374 10199 10376
rect 9876 10372 9882 10374
rect 10133 10371 10199 10374
rect 10593 10434 10659 10437
rect 11830 10434 11836 10436
rect 10593 10432 11836 10434
rect 10593 10376 10598 10432
rect 10654 10376 11836 10432
rect 10593 10374 11836 10376
rect 10593 10371 10659 10374
rect 11830 10372 11836 10374
rect 11900 10434 11906 10436
rect 13169 10434 13235 10437
rect 11900 10432 13235 10434
rect 11900 10376 13174 10432
rect 13230 10376 13235 10432
rect 11900 10374 13235 10376
rect 11900 10372 11906 10374
rect 13169 10371 13235 10374
rect 21081 10434 21147 10437
rect 22200 10434 23000 10464
rect 21081 10432 23000 10434
rect 21081 10376 21086 10432
rect 21142 10376 23000 10432
rect 21081 10374 23000 10376
rect 21081 10371 21147 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 22200 10344 23000 10374
rect 14805 10303 15125 10304
rect 6453 10296 6519 10301
rect 6453 10240 6458 10296
rect 6514 10240 6519 10296
rect 6453 10235 6519 10240
rect 9213 10298 9279 10301
rect 11053 10298 11119 10301
rect 19333 10298 19399 10301
rect 22001 10298 22067 10301
rect 9213 10296 12082 10298
rect 9213 10240 9218 10296
rect 9274 10240 11058 10296
rect 11114 10240 12082 10296
rect 9213 10238 12082 10240
rect 9213 10235 9279 10238
rect 11053 10235 11119 10238
rect 6821 10162 6887 10165
rect 9305 10162 9371 10165
rect 12022 10162 12082 10238
rect 19333 10296 22067 10298
rect 19333 10240 19338 10296
rect 19394 10240 22006 10296
rect 22062 10240 22067 10296
rect 19333 10238 22067 10240
rect 19333 10235 19399 10238
rect 22001 10235 22067 10238
rect 21173 10162 21239 10165
rect 6821 10160 11898 10162
rect 6821 10104 6826 10160
rect 6882 10104 9310 10160
rect 9366 10104 11898 10160
rect 6821 10102 11898 10104
rect 12022 10160 21239 10162
rect 12022 10104 21178 10160
rect 21234 10104 21239 10160
rect 12022 10102 21239 10104
rect 6821 10099 6887 10102
rect 9305 10099 9371 10102
rect 8293 10026 8359 10029
rect 8702 10026 8708 10028
rect 8293 10024 8708 10026
rect 8293 9968 8298 10024
rect 8354 9968 8708 10024
rect 8293 9966 8708 9968
rect 8293 9963 8359 9966
rect 8702 9964 8708 9966
rect 8772 9964 8778 10028
rect 0 9890 800 9920
rect 3417 9890 3483 9893
rect 0 9888 3483 9890
rect 0 9832 3422 9888
rect 3478 9832 3483 9888
rect 0 9830 3483 9832
rect 0 9800 800 9830
rect 3417 9827 3483 9830
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 7925 9754 7991 9757
rect 8518 9754 8524 9756
rect 7925 9752 8524 9754
rect 7925 9696 7930 9752
rect 7986 9696 8524 9752
rect 7925 9694 8524 9696
rect 7925 9691 7991 9694
rect 8518 9692 8524 9694
rect 8588 9754 8594 9756
rect 11838 9754 11898 10102
rect 21173 10099 21239 10102
rect 21357 10026 21423 10029
rect 12758 10024 21423 10026
rect 12758 9968 21362 10024
rect 21418 9968 21423 10024
rect 12758 9966 21423 9968
rect 12157 9890 12223 9893
rect 12525 9890 12591 9893
rect 12157 9888 12591 9890
rect 12157 9832 12162 9888
rect 12218 9832 12530 9888
rect 12586 9832 12591 9888
rect 12157 9830 12591 9832
rect 12157 9827 12223 9830
rect 12525 9827 12591 9830
rect 12433 9754 12499 9757
rect 12758 9754 12818 9966
rect 21357 9963 21423 9966
rect 19425 9890 19491 9893
rect 21541 9890 21607 9893
rect 22200 9890 23000 9920
rect 19425 9888 23000 9890
rect 19425 9832 19430 9888
rect 19486 9832 21546 9888
rect 21602 9832 23000 9888
rect 19425 9830 23000 9832
rect 19425 9827 19491 9830
rect 21541 9827 21607 9830
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 22200 9800 23000 9830
rect 18270 9759 18590 9760
rect 8588 9694 11162 9754
rect 11838 9752 12499 9754
rect 11838 9696 12438 9752
rect 12494 9696 12499 9752
rect 11838 9694 12499 9696
rect 8588 9692 8594 9694
rect 6494 9556 6500 9620
rect 6564 9618 6570 9620
rect 6821 9618 6887 9621
rect 6564 9616 6887 9618
rect 6564 9560 6826 9616
rect 6882 9560 6887 9616
rect 6564 9558 6887 9560
rect 6564 9556 6570 9558
rect 6821 9555 6887 9558
rect 7005 9618 7071 9621
rect 9806 9618 9812 9620
rect 7005 9616 9812 9618
rect 7005 9560 7010 9616
rect 7066 9560 9812 9616
rect 7005 9558 9812 9560
rect 7005 9555 7071 9558
rect 9806 9556 9812 9558
rect 9876 9556 9882 9620
rect 11102 9618 11162 9694
rect 12433 9691 12499 9694
rect 12574 9694 12818 9754
rect 12574 9621 12634 9694
rect 12574 9618 12683 9621
rect 11102 9616 12683 9618
rect 11102 9560 12622 9616
rect 12678 9560 12683 9616
rect 11102 9558 12683 9560
rect 12617 9555 12683 9558
rect 12985 9618 13051 9621
rect 15469 9618 15535 9621
rect 12985 9616 15535 9618
rect 12985 9560 12990 9616
rect 13046 9560 15474 9616
rect 15530 9560 15535 9616
rect 12985 9558 15535 9560
rect 12985 9555 13051 9558
rect 15469 9555 15535 9558
rect 20253 9618 20319 9621
rect 20478 9618 20484 9620
rect 20253 9616 20484 9618
rect 20253 9560 20258 9616
rect 20314 9560 20484 9616
rect 20253 9558 20484 9560
rect 20253 9555 20319 9558
rect 20478 9556 20484 9558
rect 20548 9556 20554 9620
rect 0 9482 800 9512
rect 3233 9482 3299 9485
rect 0 9480 3299 9482
rect 0 9424 3238 9480
rect 3294 9424 3299 9480
rect 0 9422 3299 9424
rect 0 9392 800 9422
rect 3233 9419 3299 9422
rect 5758 9420 5764 9484
rect 5828 9482 5834 9484
rect 7005 9482 7071 9485
rect 5828 9480 7071 9482
rect 5828 9424 7010 9480
rect 7066 9424 7071 9480
rect 5828 9422 7071 9424
rect 5828 9420 5834 9422
rect 7005 9419 7071 9422
rect 7230 9420 7236 9484
rect 7300 9482 7306 9484
rect 8017 9482 8083 9485
rect 7300 9480 8083 9482
rect 7300 9424 8022 9480
rect 8078 9424 8083 9480
rect 7300 9422 8083 9424
rect 7300 9420 7306 9422
rect 8017 9419 8083 9422
rect 8293 9482 8359 9485
rect 9213 9482 9279 9485
rect 8293 9480 9279 9482
rect 8293 9424 8298 9480
rect 8354 9424 9218 9480
rect 9274 9424 9279 9480
rect 8293 9422 9279 9424
rect 8293 9419 8359 9422
rect 9213 9419 9279 9422
rect 10174 9420 10180 9484
rect 10244 9482 10250 9484
rect 11697 9482 11763 9485
rect 10244 9480 11763 9482
rect 10244 9424 11702 9480
rect 11758 9424 11763 9480
rect 10244 9422 11763 9424
rect 10244 9420 10250 9422
rect 11697 9419 11763 9422
rect 12709 9482 12775 9485
rect 16757 9482 16823 9485
rect 12709 9480 16823 9482
rect 12709 9424 12714 9480
rect 12770 9424 16762 9480
rect 16818 9424 16823 9480
rect 12709 9422 16823 9424
rect 12709 9419 12775 9422
rect 16757 9419 16823 9422
rect 21449 9482 21515 9485
rect 22200 9482 23000 9512
rect 21449 9480 23000 9482
rect 21449 9424 21454 9480
rect 21510 9424 23000 9480
rect 21449 9422 23000 9424
rect 21449 9419 21515 9422
rect 22200 9392 23000 9422
rect 1945 9346 2011 9349
rect 6729 9346 6795 9349
rect 1945 9344 6795 9346
rect 1945 9288 1950 9344
rect 2006 9288 6734 9344
rect 6790 9288 6795 9344
rect 1945 9286 6795 9288
rect 1945 9283 2011 9286
rect 6729 9283 6795 9286
rect 9305 9346 9371 9349
rect 12985 9346 13051 9349
rect 9305 9344 14658 9346
rect 9305 9288 9310 9344
rect 9366 9288 12990 9344
rect 13046 9288 14658 9344
rect 9305 9286 14658 9288
rect 9305 9283 9371 9286
rect 12985 9283 13051 9286
rect 2865 9210 2931 9213
rect 2998 9210 3004 9212
rect 2865 9208 3004 9210
rect 2865 9152 2870 9208
rect 2926 9152 3004 9208
rect 2865 9150 3004 9152
rect 2865 9147 2931 9150
rect 2998 9148 3004 9150
rect 3068 9148 3074 9212
rect 0 9074 800 9104
rect 3141 9074 3207 9077
rect 0 9072 3207 9074
rect 0 9016 3146 9072
rect 3202 9016 3207 9072
rect 0 9014 3207 9016
rect 6732 9074 6792 9283
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 9254 9148 9260 9212
rect 9324 9210 9330 9212
rect 9489 9210 9555 9213
rect 9324 9208 9555 9210
rect 9324 9152 9494 9208
rect 9550 9152 9555 9208
rect 9324 9150 9555 9152
rect 9324 9148 9330 9150
rect 9489 9147 9555 9150
rect 9673 9210 9739 9213
rect 12198 9210 12204 9212
rect 9673 9208 12204 9210
rect 9673 9152 9678 9208
rect 9734 9152 12204 9208
rect 9673 9150 12204 9152
rect 9673 9147 9739 9150
rect 12198 9148 12204 9150
rect 12268 9148 12274 9212
rect 12617 9210 12683 9213
rect 13118 9210 13124 9212
rect 12617 9208 13124 9210
rect 12617 9152 12622 9208
rect 12678 9152 13124 9208
rect 12617 9150 13124 9152
rect 12617 9147 12683 9150
rect 13118 9148 13124 9150
rect 13188 9148 13194 9212
rect 14089 9074 14155 9077
rect 6732 9072 14155 9074
rect 6732 9016 14094 9072
rect 14150 9016 14155 9072
rect 6732 9014 14155 9016
rect 14598 9074 14658 9286
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 18045 9074 18111 9077
rect 14598 9072 18111 9074
rect 14598 9016 18050 9072
rect 18106 9016 18111 9072
rect 14598 9014 18111 9016
rect 0 8984 800 9014
rect 3141 9011 3207 9014
rect 14089 9011 14155 9014
rect 18045 9011 18111 9014
rect 21633 9074 21699 9077
rect 22200 9074 23000 9104
rect 21633 9072 23000 9074
rect 21633 9016 21638 9072
rect 21694 9016 23000 9072
rect 21633 9014 23000 9016
rect 21633 9011 21699 9014
rect 22200 8984 23000 9014
rect 3325 8938 3391 8941
rect 12525 8938 12591 8941
rect 17033 8938 17099 8941
rect 17677 8938 17743 8941
rect 18229 8938 18295 8941
rect 3325 8936 12450 8938
rect 3325 8880 3330 8936
rect 3386 8880 12450 8936
rect 3325 8878 12450 8880
rect 3325 8875 3391 8878
rect 9581 8802 9647 8805
rect 10133 8802 10199 8805
rect 4800 8800 9647 8802
rect 4800 8744 9586 8800
rect 9642 8744 9647 8800
rect 4800 8742 9647 8744
rect 4409 8736 4729 8737
rect 0 8666 800 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 1761 8666 1827 8669
rect 0 8664 1827 8666
rect 0 8608 1766 8664
rect 1822 8608 1827 8664
rect 0 8606 1827 8608
rect 0 8576 800 8606
rect 1761 8603 1827 8606
rect 1853 8530 1919 8533
rect 4800 8530 4860 8742
rect 9581 8739 9647 8742
rect 9768 8800 10199 8802
rect 9768 8744 10138 8800
rect 10194 8744 10199 8800
rect 9768 8742 10199 8744
rect 8385 8666 8451 8669
rect 9213 8666 9279 8669
rect 9768 8666 9828 8742
rect 10133 8739 10199 8742
rect 10358 8740 10364 8804
rect 10428 8802 10434 8804
rect 11053 8802 11119 8805
rect 10428 8800 11119 8802
rect 10428 8744 11058 8800
rect 11114 8744 11119 8800
rect 10428 8742 11119 8744
rect 10428 8740 10434 8742
rect 11053 8739 11119 8742
rect 12157 8800 12223 8805
rect 12157 8744 12162 8800
rect 12218 8744 12223 8800
rect 12157 8739 12223 8744
rect 12390 8802 12450 8878
rect 12525 8936 18295 8938
rect 12525 8880 12530 8936
rect 12586 8880 17038 8936
rect 17094 8880 17682 8936
rect 17738 8880 18234 8936
rect 18290 8880 18295 8936
rect 12525 8878 18295 8880
rect 12525 8875 12591 8878
rect 17033 8875 17099 8878
rect 17677 8875 17743 8878
rect 18229 8875 18295 8878
rect 12566 8802 12572 8804
rect 12390 8742 12572 8802
rect 12566 8740 12572 8742
rect 12636 8740 12642 8804
rect 13261 8802 13327 8805
rect 18137 8802 18203 8805
rect 13261 8800 18203 8802
rect 13261 8744 13266 8800
rect 13322 8744 18142 8800
rect 18198 8744 18203 8800
rect 13261 8742 18203 8744
rect 13261 8739 13327 8742
rect 18137 8739 18203 8742
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 8385 8664 9828 8666
rect 8385 8608 8390 8664
rect 8446 8608 9218 8664
rect 9274 8608 9828 8664
rect 8385 8606 9828 8608
rect 10041 8666 10107 8669
rect 10726 8666 10732 8668
rect 10041 8664 10732 8666
rect 10041 8608 10046 8664
rect 10102 8608 10732 8664
rect 10041 8606 10732 8608
rect 8385 8603 8451 8606
rect 9213 8603 9279 8606
rect 10041 8603 10107 8606
rect 10726 8604 10732 8606
rect 10796 8604 10802 8668
rect 12160 8666 12220 8739
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 12934 8666 12940 8668
rect 12160 8606 12940 8666
rect 12934 8604 12940 8606
rect 13004 8666 13010 8668
rect 17125 8666 17191 8669
rect 20713 8666 20779 8669
rect 13004 8664 17191 8666
rect 13004 8608 17130 8664
rect 17186 8608 17191 8664
rect 13004 8606 17191 8608
rect 13004 8604 13010 8606
rect 17125 8603 17191 8606
rect 20670 8664 20779 8666
rect 20670 8608 20718 8664
rect 20774 8608 20779 8664
rect 20670 8603 20779 8608
rect 21541 8666 21607 8669
rect 22200 8666 23000 8696
rect 21541 8664 23000 8666
rect 21541 8608 21546 8664
rect 21602 8608 23000 8664
rect 21541 8606 23000 8608
rect 21541 8603 21607 8606
rect 1853 8528 4860 8530
rect 1853 8472 1858 8528
rect 1914 8472 4860 8528
rect 1853 8470 4860 8472
rect 9305 8530 9371 8533
rect 16297 8530 16363 8533
rect 9305 8528 16363 8530
rect 9305 8472 9310 8528
rect 9366 8472 16302 8528
rect 16358 8472 16363 8528
rect 9305 8470 16363 8472
rect 1853 8467 1919 8470
rect 9305 8467 9371 8470
rect 16297 8467 16363 8470
rect 4889 8394 4955 8397
rect 10133 8394 10199 8397
rect 19333 8394 19399 8397
rect 4889 8392 10199 8394
rect 4889 8336 4894 8392
rect 4950 8336 10138 8392
rect 10194 8336 10199 8392
rect 4889 8334 10199 8336
rect 4889 8331 4955 8334
rect 10133 8331 10199 8334
rect 10366 8392 19399 8394
rect 10366 8336 19338 8392
rect 19394 8336 19399 8392
rect 10366 8334 19399 8336
rect 0 8258 800 8288
rect 3509 8258 3575 8261
rect 9397 8258 9463 8261
rect 10366 8258 10426 8334
rect 19333 8331 19399 8334
rect 0 8256 3575 8258
rect 0 8200 3514 8256
rect 3570 8200 3575 8256
rect 0 8198 3575 8200
rect 0 8168 800 8198
rect 3509 8195 3575 8198
rect 8296 8256 10426 8258
rect 8296 8200 9402 8256
rect 9458 8200 10426 8256
rect 8296 8198 10426 8200
rect 10869 8258 10935 8261
rect 14222 8258 14228 8260
rect 10869 8256 14228 8258
rect 10869 8200 10874 8256
rect 10930 8200 14228 8256
rect 10869 8198 14228 8200
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 1669 8122 1735 8125
rect 6913 8122 6979 8125
rect 1669 8120 6979 8122
rect 1669 8064 1674 8120
rect 1730 8064 6918 8120
rect 6974 8064 6979 8120
rect 1669 8062 6979 8064
rect 1669 8059 1735 8062
rect 6913 8059 6979 8062
rect 4153 7986 4219 7989
rect 8296 7986 8356 8198
rect 9397 8195 9463 8198
rect 10869 8195 10935 8198
rect 14222 8196 14228 8198
rect 14292 8196 14298 8260
rect 15469 8258 15535 8261
rect 20670 8258 20730 8603
rect 22200 8576 23000 8606
rect 15469 8256 20730 8258
rect 15469 8200 15474 8256
rect 15530 8200 20730 8256
rect 15469 8198 20730 8200
rect 21541 8258 21607 8261
rect 22200 8258 23000 8288
rect 21541 8256 23000 8258
rect 21541 8200 21546 8256
rect 21602 8200 23000 8256
rect 21541 8198 23000 8200
rect 15469 8195 15535 8198
rect 21541 8195 21607 8198
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 22200 8168 23000 8198
rect 14805 8127 15125 8128
rect 8702 8060 8708 8124
rect 8772 8122 8778 8124
rect 12985 8122 13051 8125
rect 8772 8120 13051 8122
rect 8772 8064 12990 8120
rect 13046 8064 13051 8120
rect 8772 8062 13051 8064
rect 8772 8060 8778 8062
rect 12985 8059 13051 8062
rect 14273 8122 14339 8125
rect 14406 8122 14412 8124
rect 14273 8120 14412 8122
rect 14273 8064 14278 8120
rect 14334 8064 14412 8120
rect 14273 8062 14412 8064
rect 14273 8059 14339 8062
rect 14406 8060 14412 8062
rect 14476 8060 14482 8124
rect 4153 7984 8356 7986
rect 4153 7928 4158 7984
rect 4214 7928 8356 7984
rect 4153 7926 8356 7928
rect 4153 7923 4219 7926
rect 9070 7924 9076 7988
rect 9140 7986 9146 7988
rect 9305 7986 9371 7989
rect 9140 7984 9371 7986
rect 9140 7928 9310 7984
rect 9366 7928 9371 7984
rect 9140 7926 9371 7928
rect 9140 7924 9146 7926
rect 9305 7923 9371 7926
rect 9673 7986 9739 7989
rect 13813 7986 13879 7989
rect 20805 7986 20871 7989
rect 9673 7984 13738 7986
rect 9673 7928 9678 7984
rect 9734 7928 13738 7984
rect 9673 7926 13738 7928
rect 9673 7923 9739 7926
rect 0 7850 800 7880
rect 1485 7850 1551 7853
rect 0 7848 1551 7850
rect 0 7792 1490 7848
rect 1546 7792 1551 7848
rect 0 7790 1551 7792
rect 0 7760 800 7790
rect 1485 7787 1551 7790
rect 2957 7850 3023 7853
rect 9438 7850 9444 7852
rect 2957 7848 9444 7850
rect 2957 7792 2962 7848
rect 3018 7792 9444 7848
rect 2957 7790 9444 7792
rect 2957 7787 3023 7790
rect 9438 7788 9444 7790
rect 9508 7788 9514 7852
rect 9622 7788 9628 7852
rect 9692 7850 9698 7852
rect 12617 7850 12683 7853
rect 9692 7848 12683 7850
rect 9692 7792 12622 7848
rect 12678 7792 12683 7848
rect 9692 7790 12683 7792
rect 13678 7850 13738 7926
rect 13813 7984 20871 7986
rect 13813 7928 13818 7984
rect 13874 7928 20810 7984
rect 20866 7928 20871 7984
rect 13813 7926 20871 7928
rect 13813 7923 13879 7926
rect 20805 7923 20871 7926
rect 15377 7850 15443 7853
rect 16021 7850 16087 7853
rect 13678 7848 16087 7850
rect 13678 7792 15382 7848
rect 15438 7792 16026 7848
rect 16082 7792 16087 7848
rect 13678 7790 16087 7792
rect 9692 7788 9698 7790
rect 12617 7787 12683 7790
rect 15377 7787 15443 7790
rect 16021 7787 16087 7790
rect 16849 7850 16915 7853
rect 20805 7850 20871 7853
rect 16849 7848 20871 7850
rect 16849 7792 16854 7848
rect 16910 7792 20810 7848
rect 20866 7792 20871 7848
rect 16849 7790 20871 7792
rect 16849 7787 16915 7790
rect 20805 7787 20871 7790
rect 21541 7850 21607 7853
rect 22200 7850 23000 7880
rect 21541 7848 23000 7850
rect 21541 7792 21546 7848
rect 21602 7792 23000 7848
rect 21541 7790 23000 7792
rect 21541 7787 21607 7790
rect 22200 7760 23000 7790
rect 9254 7652 9260 7716
rect 9324 7714 9330 7716
rect 10409 7714 10475 7717
rect 10593 7716 10659 7717
rect 9324 7712 10475 7714
rect 9324 7656 10414 7712
rect 10470 7656 10475 7712
rect 9324 7654 10475 7656
rect 9324 7652 9330 7654
rect 10409 7651 10475 7654
rect 10542 7652 10548 7716
rect 10612 7714 10659 7716
rect 10612 7712 10704 7714
rect 10654 7656 10704 7712
rect 10612 7654 10704 7656
rect 10612 7652 10659 7654
rect 10910 7652 10916 7716
rect 10980 7714 10986 7716
rect 11145 7714 11211 7717
rect 10980 7712 11211 7714
rect 10980 7656 11150 7712
rect 11206 7656 11211 7712
rect 10980 7654 11211 7656
rect 10980 7652 10986 7654
rect 10593 7651 10659 7652
rect 11145 7651 11211 7654
rect 12249 7714 12315 7717
rect 13077 7714 13143 7717
rect 12249 7712 13143 7714
rect 12249 7656 12254 7712
rect 12310 7656 13082 7712
rect 13138 7656 13143 7712
rect 12249 7654 13143 7656
rect 12249 7651 12315 7654
rect 13077 7651 13143 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 4797 7578 4863 7581
rect 5349 7578 5415 7581
rect 6913 7580 6979 7581
rect 4797 7576 5415 7578
rect 4797 7520 4802 7576
rect 4858 7520 5354 7576
rect 5410 7520 5415 7576
rect 4797 7518 5415 7520
rect 4797 7515 4863 7518
rect 5349 7515 5415 7518
rect 6862 7516 6868 7580
rect 6932 7578 6979 7580
rect 10593 7578 10659 7581
rect 13353 7580 13419 7581
rect 13302 7578 13308 7580
rect 6932 7576 10659 7578
rect 6974 7520 10598 7576
rect 10654 7520 10659 7576
rect 6932 7518 10659 7520
rect 13262 7518 13308 7578
rect 13372 7576 13419 7580
rect 13414 7520 13419 7576
rect 6932 7516 6979 7518
rect 6913 7515 6979 7516
rect 10593 7515 10659 7518
rect 13302 7516 13308 7518
rect 13372 7516 13419 7520
rect 13353 7515 13419 7516
rect 13813 7578 13879 7581
rect 14590 7578 14596 7580
rect 13813 7576 14596 7578
rect 13813 7520 13818 7576
rect 13874 7520 14596 7576
rect 13813 7518 14596 7520
rect 13813 7515 13879 7518
rect 14590 7516 14596 7518
rect 14660 7578 14666 7580
rect 18137 7578 18203 7581
rect 14660 7576 18203 7578
rect 14660 7520 18142 7576
rect 18198 7520 18203 7576
rect 14660 7518 18203 7520
rect 14660 7516 14666 7518
rect 18137 7515 18203 7518
rect 0 7442 800 7472
rect 3233 7442 3299 7445
rect 0 7440 3299 7442
rect 0 7384 3238 7440
rect 3294 7384 3299 7440
rect 0 7382 3299 7384
rect 0 7352 800 7382
rect 3233 7379 3299 7382
rect 3918 7380 3924 7444
rect 3988 7442 3994 7444
rect 8518 7442 8524 7444
rect 3988 7382 8524 7442
rect 3988 7380 3994 7382
rect 8518 7380 8524 7382
rect 8588 7380 8594 7444
rect 8753 7442 8819 7445
rect 17585 7442 17651 7445
rect 8753 7440 17651 7442
rect 8753 7384 8758 7440
rect 8814 7384 17590 7440
rect 17646 7384 17651 7440
rect 8753 7382 17651 7384
rect 8753 7379 8819 7382
rect 17585 7379 17651 7382
rect 19241 7442 19307 7445
rect 22200 7442 23000 7472
rect 19241 7440 23000 7442
rect 19241 7384 19246 7440
rect 19302 7384 23000 7440
rect 19241 7382 23000 7384
rect 19241 7379 19307 7382
rect 22200 7352 23000 7382
rect 2405 7306 2471 7309
rect 6913 7306 6979 7309
rect 9949 7306 10015 7309
rect 2405 7304 10015 7306
rect 2405 7248 2410 7304
rect 2466 7248 6918 7304
rect 6974 7248 9954 7304
rect 10010 7248 10015 7304
rect 2405 7246 10015 7248
rect 2405 7243 2471 7246
rect 6913 7243 6979 7246
rect 9949 7243 10015 7246
rect 10593 7306 10659 7309
rect 11421 7306 11487 7309
rect 10593 7304 11487 7306
rect 10593 7248 10598 7304
rect 10654 7248 11426 7304
rect 11482 7248 11487 7304
rect 10593 7246 11487 7248
rect 10593 7243 10659 7246
rect 11421 7243 11487 7246
rect 12198 7244 12204 7308
rect 12268 7306 12274 7308
rect 16665 7306 16731 7309
rect 12268 7304 16731 7306
rect 12268 7248 16670 7304
rect 16726 7248 16731 7304
rect 12268 7246 16731 7248
rect 12268 7244 12274 7246
rect 16665 7243 16731 7246
rect 2129 7170 2195 7173
rect 5901 7170 5967 7173
rect 2129 7168 5967 7170
rect 2129 7112 2134 7168
rect 2190 7112 5906 7168
rect 5962 7112 5967 7168
rect 2129 7110 5967 7112
rect 2129 7107 2195 7110
rect 5901 7107 5967 7110
rect 9121 7170 9187 7173
rect 9622 7170 9628 7172
rect 9121 7168 9628 7170
rect 9121 7112 9126 7168
rect 9182 7112 9628 7168
rect 9121 7110 9628 7112
rect 9121 7107 9187 7110
rect 9622 7108 9628 7110
rect 9692 7108 9698 7172
rect 9806 7108 9812 7172
rect 9876 7170 9882 7172
rect 10593 7170 10659 7173
rect 12198 7170 12204 7172
rect 9876 7168 12204 7170
rect 9876 7112 10598 7168
rect 10654 7112 12204 7168
rect 9876 7110 12204 7112
rect 9876 7108 9882 7110
rect 10593 7107 10659 7110
rect 12198 7108 12204 7110
rect 12268 7108 12274 7172
rect 16757 7170 16823 7173
rect 21449 7170 21515 7173
rect 16757 7168 21515 7170
rect 16757 7112 16762 7168
rect 16818 7112 21454 7168
rect 21510 7112 21515 7168
rect 16757 7110 21515 7112
rect 16757 7107 16823 7110
rect 21449 7107 21515 7110
rect 7874 7104 8194 7105
rect 0 7034 800 7064
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 1485 7034 1551 7037
rect 0 7032 1551 7034
rect 0 6976 1490 7032
rect 1546 6976 1551 7032
rect 0 6974 1551 6976
rect 0 6944 800 6974
rect 1485 6971 1551 6974
rect 2313 7034 2379 7037
rect 6269 7034 6335 7037
rect 10869 7034 10935 7037
rect 11145 7034 11211 7037
rect 2313 7032 5412 7034
rect 2313 6976 2318 7032
rect 2374 6976 5412 7032
rect 2313 6974 5412 6976
rect 2313 6971 2379 6974
rect 5352 6901 5412 6974
rect 6269 7032 7804 7034
rect 6269 6976 6274 7032
rect 6330 6976 7804 7032
rect 6269 6974 7804 6976
rect 6269 6971 6335 6974
rect 1485 6898 1551 6901
rect 4061 6898 4127 6901
rect 1485 6896 4127 6898
rect 1485 6840 1490 6896
rect 1546 6840 4066 6896
rect 4122 6840 4127 6896
rect 1485 6838 4127 6840
rect 1485 6835 1551 6838
rect 4061 6835 4127 6838
rect 4613 6898 4679 6901
rect 4838 6898 4844 6900
rect 4613 6896 4844 6898
rect 4613 6840 4618 6896
rect 4674 6840 4844 6896
rect 4613 6838 4844 6840
rect 4613 6835 4679 6838
rect 4838 6836 4844 6838
rect 4908 6836 4914 6900
rect 5349 6896 5415 6901
rect 5349 6840 5354 6896
rect 5410 6840 5415 6896
rect 5349 6835 5415 6840
rect 6494 6836 6500 6900
rect 6564 6898 6570 6900
rect 6637 6898 6703 6901
rect 6564 6896 6703 6898
rect 6564 6840 6642 6896
rect 6698 6840 6703 6896
rect 6564 6838 6703 6840
rect 7744 6898 7804 6974
rect 8342 7032 11211 7034
rect 8342 6976 10874 7032
rect 10930 6976 11150 7032
rect 11206 6976 11211 7032
rect 8342 6974 11211 6976
rect 8342 6898 8402 6974
rect 10869 6971 10935 6974
rect 11145 6971 11211 6974
rect 11421 7034 11487 7037
rect 12341 7034 12407 7037
rect 17033 7034 17099 7037
rect 18413 7034 18479 7037
rect 11421 7032 12036 7034
rect 11421 6976 11426 7032
rect 11482 6976 12036 7032
rect 11421 6974 12036 6976
rect 11421 6971 11487 6974
rect 7744 6838 8402 6898
rect 6564 6836 6570 6838
rect 6637 6835 6703 6838
rect 10174 6836 10180 6900
rect 10244 6898 10250 6900
rect 10317 6898 10383 6901
rect 10244 6896 10383 6898
rect 10244 6840 10322 6896
rect 10378 6840 10383 6896
rect 10244 6838 10383 6840
rect 10244 6836 10250 6838
rect 10317 6835 10383 6838
rect 10501 6898 10567 6901
rect 11830 6898 11836 6900
rect 10501 6896 11836 6898
rect 10501 6840 10506 6896
rect 10562 6840 11836 6896
rect 10501 6838 11836 6840
rect 10501 6835 10567 6838
rect 11830 6836 11836 6838
rect 11900 6836 11906 6900
rect 11976 6898 12036 6974
rect 12341 7032 14658 7034
rect 12341 6976 12346 7032
rect 12402 6976 14658 7032
rect 12341 6974 14658 6976
rect 12341 6971 12407 6974
rect 12433 6898 12499 6901
rect 11976 6896 12499 6898
rect 11976 6840 12438 6896
rect 12494 6840 12499 6896
rect 11976 6838 12499 6840
rect 14598 6898 14658 6974
rect 17033 7032 18479 7034
rect 17033 6976 17038 7032
rect 17094 6976 18418 7032
rect 18474 6976 18479 7032
rect 17033 6974 18479 6976
rect 17033 6971 17099 6974
rect 18413 6971 18479 6974
rect 19241 7034 19307 7037
rect 22200 7034 23000 7064
rect 19241 7032 23000 7034
rect 19241 6976 19246 7032
rect 19302 6976 23000 7032
rect 19241 6974 23000 6976
rect 19241 6971 19307 6974
rect 22200 6944 23000 6974
rect 18965 6898 19031 6901
rect 14598 6896 19031 6898
rect 14598 6840 18970 6896
rect 19026 6840 19031 6896
rect 14598 6838 19031 6840
rect 12433 6835 12499 6838
rect 18965 6835 19031 6838
rect 3601 6762 3667 6765
rect 5533 6762 5599 6765
rect 3601 6760 5599 6762
rect 3601 6704 3606 6760
rect 3662 6704 5538 6760
rect 5594 6704 5599 6760
rect 3601 6702 5599 6704
rect 3601 6699 3667 6702
rect 5533 6699 5599 6702
rect 6177 6762 6243 6765
rect 7557 6762 7623 6765
rect 6177 6760 7623 6762
rect 6177 6704 6182 6760
rect 6238 6704 7562 6760
rect 7618 6704 7623 6760
rect 6177 6702 7623 6704
rect 6177 6699 6243 6702
rect 7557 6699 7623 6702
rect 9857 6762 9923 6765
rect 10174 6762 10180 6764
rect 9857 6760 10180 6762
rect 9857 6704 9862 6760
rect 9918 6704 10180 6760
rect 9857 6702 10180 6704
rect 9857 6699 9923 6702
rect 10174 6700 10180 6702
rect 10244 6700 10250 6764
rect 10961 6762 11027 6765
rect 12157 6762 12223 6765
rect 13261 6762 13327 6765
rect 10961 6760 13327 6762
rect 10961 6704 10966 6760
rect 11022 6704 12162 6760
rect 12218 6704 13266 6760
rect 13322 6704 13327 6760
rect 10961 6702 13327 6704
rect 10961 6699 11027 6702
rect 12157 6699 12223 6702
rect 13261 6699 13327 6702
rect 13997 6762 14063 6765
rect 16757 6762 16823 6765
rect 13997 6760 16823 6762
rect 13997 6704 14002 6760
rect 14058 6704 16762 6760
rect 16818 6704 16823 6760
rect 13997 6702 16823 6704
rect 13997 6699 14063 6702
rect 16757 6699 16823 6702
rect 5625 6626 5691 6629
rect 8477 6626 8543 6629
rect 9397 6628 9463 6629
rect 9397 6626 9444 6628
rect 5625 6624 8543 6626
rect 5625 6568 5630 6624
rect 5686 6568 8482 6624
rect 8538 6568 8543 6624
rect 5625 6566 8543 6568
rect 9352 6624 9444 6626
rect 9352 6568 9402 6624
rect 9352 6566 9444 6568
rect 5625 6563 5691 6566
rect 8477 6563 8543 6566
rect 9397 6564 9444 6566
rect 9508 6564 9514 6628
rect 12525 6626 12591 6629
rect 14549 6626 14615 6629
rect 16573 6626 16639 6629
rect 17585 6626 17651 6629
rect 12525 6624 17651 6626
rect 12525 6568 12530 6624
rect 12586 6568 14554 6624
rect 14610 6568 16578 6624
rect 16634 6568 17590 6624
rect 17646 6568 17651 6624
rect 12525 6566 17651 6568
rect 9397 6563 9463 6564
rect 12525 6563 12591 6566
rect 14549 6563 14615 6566
rect 16573 6563 16639 6566
rect 17585 6563 17651 6566
rect 4409 6560 4729 6561
rect 0 6490 800 6520
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 3233 6490 3299 6493
rect 0 6488 3299 6490
rect 0 6432 3238 6488
rect 3294 6432 3299 6488
rect 0 6430 3299 6432
rect 0 6400 800 6430
rect 3233 6427 3299 6430
rect 3785 6488 3851 6493
rect 3785 6432 3790 6488
rect 3846 6432 3851 6488
rect 3785 6427 3851 6432
rect 5993 6490 6059 6493
rect 9121 6490 9187 6493
rect 5993 6488 9187 6490
rect 5993 6432 5998 6488
rect 6054 6432 9126 6488
rect 9182 6432 9187 6488
rect 5993 6430 9187 6432
rect 5993 6427 6059 6430
rect 9121 6427 9187 6430
rect 9673 6490 9739 6493
rect 11145 6490 11211 6493
rect 9673 6488 11211 6490
rect 9673 6432 9678 6488
rect 9734 6432 11150 6488
rect 11206 6432 11211 6488
rect 9673 6430 11211 6432
rect 9673 6427 9739 6430
rect 11145 6427 11211 6430
rect 19057 6490 19123 6493
rect 20253 6490 20319 6493
rect 19057 6488 20319 6490
rect 19057 6432 19062 6488
rect 19118 6432 20258 6488
rect 20314 6432 20319 6488
rect 19057 6430 20319 6432
rect 19057 6427 19123 6430
rect 20253 6427 20319 6430
rect 20437 6490 20503 6493
rect 22001 6490 22067 6493
rect 22200 6490 23000 6520
rect 20437 6488 23000 6490
rect 20437 6432 20442 6488
rect 20498 6432 22006 6488
rect 22062 6432 23000 6488
rect 20437 6430 23000 6432
rect 20437 6427 20503 6430
rect 22001 6427 22067 6430
rect 3788 6354 3848 6427
rect 22200 6400 23000 6430
rect 4797 6354 4863 6357
rect 7373 6354 7439 6357
rect 3788 6352 4863 6354
rect 3788 6296 4802 6352
rect 4858 6296 4863 6352
rect 3788 6294 4863 6296
rect 4797 6291 4863 6294
rect 6502 6352 7439 6354
rect 6502 6296 7378 6352
rect 7434 6296 7439 6352
rect 6502 6294 7439 6296
rect 6502 6221 6562 6294
rect 7373 6291 7439 6294
rect 7557 6354 7623 6357
rect 7741 6354 7807 6357
rect 8937 6356 9003 6357
rect 7557 6352 7807 6354
rect 7557 6296 7562 6352
rect 7618 6296 7746 6352
rect 7802 6296 7807 6352
rect 7557 6294 7807 6296
rect 7557 6291 7623 6294
rect 7741 6291 7807 6294
rect 8886 6292 8892 6356
rect 8956 6354 9003 6356
rect 9121 6354 9187 6357
rect 10358 6354 10364 6356
rect 8956 6352 9048 6354
rect 8998 6296 9048 6352
rect 8956 6294 9048 6296
rect 9121 6352 10364 6354
rect 9121 6296 9126 6352
rect 9182 6296 10364 6352
rect 9121 6294 10364 6296
rect 8956 6292 9003 6294
rect 8937 6291 9003 6292
rect 9121 6291 9187 6294
rect 10358 6292 10364 6294
rect 10428 6354 10434 6356
rect 11421 6354 11487 6357
rect 10428 6352 11487 6354
rect 10428 6296 11426 6352
rect 11482 6296 11487 6352
rect 10428 6294 11487 6296
rect 10428 6292 10434 6294
rect 11421 6291 11487 6294
rect 14549 6354 14615 6357
rect 15653 6354 15719 6357
rect 14549 6352 15719 6354
rect 14549 6296 14554 6352
rect 14610 6296 15658 6352
rect 15714 6296 15719 6352
rect 14549 6294 15719 6296
rect 14549 6291 14615 6294
rect 15653 6291 15719 6294
rect 18597 6354 18663 6357
rect 19885 6354 19951 6357
rect 18597 6352 19951 6354
rect 18597 6296 18602 6352
rect 18658 6296 19890 6352
rect 19946 6296 19951 6352
rect 18597 6294 19951 6296
rect 18597 6291 18663 6294
rect 19885 6291 19951 6294
rect 1117 6218 1183 6221
rect 4245 6218 4311 6221
rect 6177 6218 6243 6221
rect 1117 6216 6243 6218
rect 1117 6160 1122 6216
rect 1178 6160 4250 6216
rect 4306 6160 6182 6216
rect 6238 6160 6243 6216
rect 1117 6158 6243 6160
rect 1117 6155 1183 6158
rect 4245 6155 4311 6158
rect 6177 6155 6243 6158
rect 6453 6216 6562 6221
rect 6453 6160 6458 6216
rect 6514 6160 6562 6216
rect 6453 6158 6562 6160
rect 6729 6218 6795 6221
rect 8017 6218 8083 6221
rect 9990 6218 9996 6220
rect 6729 6216 9996 6218
rect 6729 6160 6734 6216
rect 6790 6160 8022 6216
rect 8078 6160 9996 6216
rect 6729 6158 9996 6160
rect 6453 6155 6519 6158
rect 6729 6155 6795 6158
rect 8017 6155 8083 6158
rect 9990 6156 9996 6158
rect 10060 6156 10066 6220
rect 10174 6156 10180 6220
rect 10244 6218 10250 6220
rect 11605 6218 11671 6221
rect 10244 6216 11671 6218
rect 10244 6160 11610 6216
rect 11666 6160 11671 6216
rect 10244 6158 11671 6160
rect 10244 6156 10250 6158
rect 0 6082 800 6112
rect 1485 6082 1551 6085
rect 0 6080 1551 6082
rect 0 6024 1490 6080
rect 1546 6024 1551 6080
rect 0 6022 1551 6024
rect 0 5992 800 6022
rect 1485 6019 1551 6022
rect 2865 6082 2931 6085
rect 2865 6080 7804 6082
rect 2865 6024 2870 6080
rect 2926 6024 7804 6080
rect 2865 6022 7804 6024
rect 2865 6019 2931 6022
rect 4153 5946 4219 5949
rect 5533 5946 5599 5949
rect 4153 5944 5599 5946
rect 4153 5888 4158 5944
rect 4214 5888 5538 5944
rect 5594 5888 5599 5944
rect 4153 5886 5599 5888
rect 4153 5883 4219 5886
rect 5533 5883 5599 5886
rect 933 5810 999 5813
rect 6177 5810 6243 5813
rect 7557 5810 7623 5813
rect 933 5808 7623 5810
rect 933 5752 938 5808
rect 994 5752 6182 5808
rect 6238 5752 7562 5808
rect 7618 5752 7623 5808
rect 933 5750 7623 5752
rect 7744 5810 7804 6022
rect 9673 6080 9739 6085
rect 9673 6024 9678 6080
rect 9734 6024 9739 6080
rect 9673 6019 9739 6024
rect 9998 6082 10058 6156
rect 11605 6155 11671 6158
rect 12198 6156 12204 6220
rect 12268 6218 12274 6220
rect 13169 6218 13235 6221
rect 12268 6216 13235 6218
rect 12268 6160 13174 6216
rect 13230 6160 13235 6216
rect 12268 6158 13235 6160
rect 12268 6156 12274 6158
rect 13169 6155 13235 6158
rect 14365 6216 14431 6221
rect 14365 6160 14370 6216
rect 14426 6160 14431 6216
rect 14365 6155 14431 6160
rect 18781 6220 18847 6221
rect 18781 6216 18828 6220
rect 18892 6218 18898 6220
rect 18781 6160 18786 6216
rect 18781 6156 18828 6160
rect 18892 6158 18938 6218
rect 18892 6156 18898 6158
rect 18781 6155 18847 6156
rect 14368 6082 14428 6155
rect 9998 6022 14428 6082
rect 20161 6082 20227 6085
rect 21081 6082 21147 6085
rect 22200 6082 23000 6112
rect 20161 6080 23000 6082
rect 20161 6024 20166 6080
rect 20222 6024 21086 6080
rect 21142 6024 23000 6080
rect 20161 6022 23000 6024
rect 20161 6019 20227 6022
rect 21081 6019 21147 6022
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 9676 5946 9736 6019
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 22200 5992 23000 6022
rect 14805 5951 15125 5952
rect 9949 5946 10015 5949
rect 9676 5944 10015 5946
rect 9676 5888 9954 5944
rect 10010 5888 10015 5944
rect 9676 5886 10015 5888
rect 9949 5883 10015 5886
rect 10593 5946 10659 5949
rect 11513 5946 11579 5949
rect 10593 5944 11579 5946
rect 10593 5888 10598 5944
rect 10654 5888 11518 5944
rect 11574 5888 11579 5944
rect 10593 5886 11579 5888
rect 10593 5883 10659 5886
rect 11513 5883 11579 5886
rect 11881 5946 11947 5949
rect 12341 5948 12407 5949
rect 12014 5946 12020 5948
rect 11881 5944 12020 5946
rect 11881 5888 11886 5944
rect 11942 5888 12020 5944
rect 11881 5886 12020 5888
rect 11881 5883 11947 5886
rect 12014 5884 12020 5886
rect 12084 5884 12090 5948
rect 12341 5946 12388 5948
rect 12296 5944 12388 5946
rect 12296 5888 12346 5944
rect 12296 5886 12388 5888
rect 12341 5884 12388 5886
rect 12452 5884 12458 5948
rect 12341 5883 12407 5884
rect 11094 5810 11100 5812
rect 7744 5750 11100 5810
rect 933 5747 999 5750
rect 6177 5747 6243 5750
rect 7557 5747 7623 5750
rect 11094 5748 11100 5750
rect 11164 5748 11170 5812
rect 11830 5748 11836 5812
rect 11900 5810 11906 5812
rect 12801 5810 12867 5813
rect 11900 5808 12867 5810
rect 11900 5752 12806 5808
rect 12862 5752 12867 5808
rect 11900 5750 12867 5752
rect 11900 5748 11906 5750
rect 12801 5747 12867 5750
rect 13353 5810 13419 5813
rect 19057 5810 19123 5813
rect 13353 5808 19123 5810
rect 13353 5752 13358 5808
rect 13414 5752 19062 5808
rect 19118 5752 19123 5808
rect 13353 5750 19123 5752
rect 13353 5747 13419 5750
rect 19057 5747 19123 5750
rect 20478 5748 20484 5812
rect 20548 5810 20554 5812
rect 20621 5810 20687 5813
rect 20548 5808 20687 5810
rect 20548 5752 20626 5808
rect 20682 5752 20687 5808
rect 20548 5750 20687 5752
rect 20548 5748 20554 5750
rect 20621 5747 20687 5750
rect 0 5674 800 5704
rect 1209 5674 1275 5677
rect 0 5672 1275 5674
rect 0 5616 1214 5672
rect 1270 5616 1275 5672
rect 0 5614 1275 5616
rect 0 5584 800 5614
rect 1209 5611 1275 5614
rect 2998 5612 3004 5676
rect 3068 5674 3074 5676
rect 3233 5674 3299 5677
rect 5809 5674 5875 5677
rect 3068 5672 5875 5674
rect 3068 5616 3238 5672
rect 3294 5616 5814 5672
rect 5870 5616 5875 5672
rect 3068 5614 5875 5616
rect 3068 5612 3074 5614
rect 3233 5611 3299 5614
rect 5809 5611 5875 5614
rect 5993 5674 6059 5677
rect 7189 5674 7255 5677
rect 5993 5672 7255 5674
rect 5993 5616 5998 5672
rect 6054 5616 7194 5672
rect 7250 5616 7255 5672
rect 5993 5614 7255 5616
rect 5993 5611 6059 5614
rect 7189 5611 7255 5614
rect 7414 5612 7420 5676
rect 7484 5674 7490 5676
rect 12157 5674 12223 5677
rect 7484 5672 12223 5674
rect 7484 5616 12162 5672
rect 12218 5616 12223 5672
rect 7484 5614 12223 5616
rect 7484 5612 7490 5614
rect 6269 5538 6335 5541
rect 7422 5538 7482 5612
rect 12157 5611 12223 5614
rect 21541 5674 21607 5677
rect 22200 5674 23000 5704
rect 21541 5672 23000 5674
rect 21541 5616 21546 5672
rect 21602 5616 23000 5672
rect 21541 5614 23000 5616
rect 21541 5611 21607 5614
rect 22200 5584 23000 5614
rect 6269 5536 7482 5538
rect 6269 5480 6274 5536
rect 6330 5480 7482 5536
rect 6269 5478 7482 5480
rect 8017 5538 8083 5541
rect 8937 5538 9003 5541
rect 8017 5536 9003 5538
rect 8017 5480 8022 5536
rect 8078 5480 8942 5536
rect 8998 5480 9003 5536
rect 8017 5478 9003 5480
rect 6269 5475 6335 5478
rect 8017 5475 8083 5478
rect 8937 5475 9003 5478
rect 9673 5538 9739 5541
rect 10777 5540 10843 5541
rect 9806 5538 9812 5540
rect 9673 5536 9812 5538
rect 9673 5480 9678 5536
rect 9734 5480 9812 5536
rect 9673 5478 9812 5480
rect 9673 5475 9739 5478
rect 9806 5476 9812 5478
rect 9876 5476 9882 5540
rect 10726 5476 10732 5540
rect 10796 5538 10843 5540
rect 10796 5536 10888 5538
rect 10838 5480 10888 5536
rect 10796 5478 10888 5480
rect 10796 5476 10843 5478
rect 10777 5475 10843 5476
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 3785 5402 3851 5405
rect 6729 5404 6795 5405
rect 3918 5402 3924 5404
rect 3785 5400 3924 5402
rect 3785 5344 3790 5400
rect 3846 5344 3924 5400
rect 3785 5342 3924 5344
rect 3785 5339 3851 5342
rect 3918 5340 3924 5342
rect 3988 5340 3994 5404
rect 6678 5340 6684 5404
rect 6748 5402 6795 5404
rect 6748 5400 6840 5402
rect 6790 5344 6840 5400
rect 6748 5342 6840 5344
rect 6748 5340 6795 5342
rect 7230 5340 7236 5404
rect 7300 5402 7306 5404
rect 7465 5402 7531 5405
rect 7300 5400 9690 5402
rect 7300 5344 7470 5400
rect 7526 5344 9690 5400
rect 7300 5342 9690 5344
rect 7300 5340 7306 5342
rect 6729 5339 6795 5340
rect 7465 5339 7531 5342
rect 0 5266 800 5296
rect 1301 5266 1367 5269
rect 0 5264 1367 5266
rect 0 5208 1306 5264
rect 1362 5208 1367 5264
rect 0 5206 1367 5208
rect 0 5176 800 5206
rect 1301 5203 1367 5206
rect 3693 5266 3759 5269
rect 7925 5266 7991 5269
rect 3693 5264 7991 5266
rect 3693 5208 3698 5264
rect 3754 5208 7930 5264
rect 7986 5208 7991 5264
rect 3693 5206 7991 5208
rect 3693 5203 3759 5206
rect 7925 5203 7991 5206
rect 8518 5204 8524 5268
rect 8588 5266 8594 5268
rect 8661 5266 8727 5269
rect 8588 5264 8727 5266
rect 8588 5208 8666 5264
rect 8722 5208 8727 5264
rect 8588 5206 8727 5208
rect 9630 5266 9690 5342
rect 14549 5266 14615 5269
rect 9630 5264 14615 5266
rect 9630 5208 14554 5264
rect 14610 5208 14615 5264
rect 9630 5206 14615 5208
rect 8588 5204 8594 5206
rect 8661 5203 8727 5206
rect 14549 5203 14615 5206
rect 19977 5266 20043 5269
rect 21449 5266 21515 5269
rect 22200 5266 23000 5296
rect 19977 5264 23000 5266
rect 19977 5208 19982 5264
rect 20038 5208 21454 5264
rect 21510 5208 23000 5264
rect 19977 5206 23000 5208
rect 19977 5203 20043 5206
rect 21449 5203 21515 5206
rect 22200 5176 23000 5206
rect 2037 5130 2103 5133
rect 7373 5130 7439 5133
rect 2037 5128 7439 5130
rect 2037 5072 2042 5128
rect 2098 5072 7378 5128
rect 7434 5072 7439 5128
rect 2037 5070 7439 5072
rect 2037 5067 2103 5070
rect 7373 5067 7439 5070
rect 10317 5130 10383 5133
rect 21265 5130 21331 5133
rect 10317 5128 21331 5130
rect 10317 5072 10322 5128
rect 10378 5072 21270 5128
rect 21326 5072 21331 5128
rect 10317 5070 21331 5072
rect 10317 5067 10383 5070
rect 21265 5067 21331 5070
rect 1761 4994 1827 4997
rect 7281 4994 7347 4997
rect 13169 4996 13235 4997
rect 13118 4994 13124 4996
rect 1761 4992 7347 4994
rect 1761 4936 1766 4992
rect 1822 4936 7286 4992
rect 7342 4936 7347 4992
rect 1761 4934 7347 4936
rect 13078 4934 13124 4994
rect 13188 4992 13235 4996
rect 13230 4936 13235 4992
rect 1761 4931 1827 4934
rect 7281 4931 7347 4934
rect 13118 4932 13124 4934
rect 13188 4932 13235 4936
rect 13169 4931 13235 4932
rect 14365 4996 14431 4997
rect 14365 4992 14412 4996
rect 14476 4994 14482 4996
rect 14365 4936 14370 4992
rect 14365 4932 14412 4936
rect 14476 4934 14522 4994
rect 14476 4932 14482 4934
rect 14365 4931 14431 4932
rect 7874 4928 8194 4929
rect 0 4858 800 4888
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 2773 4858 2839 4861
rect 3877 4858 3943 4861
rect 11830 4858 11836 4860
rect 0 4856 3943 4858
rect 0 4800 2778 4856
rect 2834 4800 3882 4856
rect 3938 4800 3943 4856
rect 0 4798 3943 4800
rect 0 4768 800 4798
rect 2773 4795 2839 4798
rect 3877 4795 3943 4798
rect 9630 4798 11836 4858
rect 7005 4724 7071 4725
rect 7005 4722 7052 4724
rect 6960 4720 7052 4722
rect 6960 4664 7010 4720
rect 6960 4662 7052 4664
rect 7005 4660 7052 4662
rect 7116 4660 7122 4724
rect 7281 4722 7347 4725
rect 8753 4722 8819 4725
rect 7281 4720 8819 4722
rect 7281 4664 7286 4720
rect 7342 4664 8758 4720
rect 8814 4664 8819 4720
rect 7281 4662 8819 4664
rect 7005 4659 7071 4660
rect 7281 4659 7347 4662
rect 8753 4659 8819 4662
rect 5809 4586 5875 4589
rect 6269 4586 6335 4589
rect 9630 4586 9690 4798
rect 11830 4796 11836 4798
rect 11900 4796 11906 4860
rect 18137 4858 18203 4861
rect 19977 4858 20043 4861
rect 18137 4856 20043 4858
rect 18137 4800 18142 4856
rect 18198 4800 19982 4856
rect 20038 4800 20043 4856
rect 18137 4798 20043 4800
rect 18137 4795 18203 4798
rect 19977 4795 20043 4798
rect 21449 4858 21515 4861
rect 22200 4858 23000 4888
rect 21449 4856 23000 4858
rect 21449 4800 21454 4856
rect 21510 4800 23000 4856
rect 21449 4798 23000 4800
rect 21449 4795 21515 4798
rect 22200 4768 23000 4798
rect 12566 4660 12572 4724
rect 12636 4722 12642 4724
rect 13537 4722 13603 4725
rect 14365 4722 14431 4725
rect 12636 4720 14431 4722
rect 12636 4664 13542 4720
rect 13598 4664 14370 4720
rect 14426 4664 14431 4720
rect 12636 4662 14431 4664
rect 12636 4660 12642 4662
rect 13537 4659 13603 4662
rect 14365 4659 14431 4662
rect 5809 4584 9690 4586
rect 5809 4528 5814 4584
rect 5870 4528 6274 4584
rect 6330 4528 9690 4584
rect 5809 4526 9690 4528
rect 9949 4586 10015 4589
rect 16113 4586 16179 4589
rect 9949 4584 16179 4586
rect 9949 4528 9954 4584
rect 10010 4528 16118 4584
rect 16174 4528 16179 4584
rect 9949 4526 16179 4528
rect 5809 4523 5875 4526
rect 6269 4523 6335 4526
rect 9949 4523 10015 4526
rect 16113 4523 16179 4526
rect 19149 4586 19215 4589
rect 19149 4584 19258 4586
rect 19149 4528 19154 4584
rect 19210 4528 19258 4584
rect 19149 4523 19258 4528
rect 0 4450 800 4480
rect 1301 4450 1367 4453
rect 0 4448 1367 4450
rect 0 4392 1306 4448
rect 1362 4392 1367 4448
rect 0 4390 1367 4392
rect 0 4360 800 4390
rect 1301 4387 1367 4390
rect 5809 4450 5875 4453
rect 8569 4450 8635 4453
rect 5809 4448 8635 4450
rect 5809 4392 5814 4448
rect 5870 4392 8574 4448
rect 8630 4392 8635 4448
rect 5809 4390 8635 4392
rect 5809 4387 5875 4390
rect 8569 4387 8635 4390
rect 11789 4450 11855 4453
rect 12341 4450 12407 4453
rect 15837 4450 15903 4453
rect 11789 4448 15903 4450
rect 11789 4392 11794 4448
rect 11850 4392 12346 4448
rect 12402 4392 15842 4448
rect 15898 4392 15903 4448
rect 11789 4390 15903 4392
rect 19198 4450 19258 4523
rect 21449 4450 21515 4453
rect 22200 4450 23000 4480
rect 19198 4448 23000 4450
rect 19198 4392 21454 4448
rect 21510 4392 23000 4448
rect 19198 4390 23000 4392
rect 11789 4387 11855 4390
rect 12341 4387 12407 4390
rect 15837 4387 15903 4390
rect 21449 4387 21515 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 22200 4360 23000 4390
rect 18270 4319 18590 4320
rect 5349 4314 5415 4317
rect 7598 4314 7604 4316
rect 5349 4312 7604 4314
rect 5349 4256 5354 4312
rect 5410 4256 7604 4312
rect 5349 4254 7604 4256
rect 5349 4251 5415 4254
rect 7598 4252 7604 4254
rect 7668 4314 7674 4316
rect 7668 4254 8954 4314
rect 7668 4252 7674 4254
rect 4613 4178 4679 4181
rect 8661 4178 8727 4181
rect 4613 4176 8727 4178
rect 4613 4120 4618 4176
rect 4674 4120 8666 4176
rect 8722 4120 8727 4176
rect 4613 4118 8727 4120
rect 8894 4178 8954 4254
rect 14733 4178 14799 4181
rect 8894 4176 14799 4178
rect 8894 4120 14738 4176
rect 14794 4120 14799 4176
rect 8894 4118 14799 4120
rect 4613 4115 4679 4118
rect 8661 4115 8727 4118
rect 14733 4115 14799 4118
rect 18229 4178 18295 4181
rect 19149 4178 19215 4181
rect 18229 4176 19215 4178
rect 18229 4120 18234 4176
rect 18290 4120 19154 4176
rect 19210 4120 19215 4176
rect 18229 4118 19215 4120
rect 18229 4115 18295 4118
rect 19149 4115 19215 4118
rect 0 4042 800 4072
rect 1301 4042 1367 4045
rect 0 4040 1367 4042
rect 0 3984 1306 4040
rect 1362 3984 1367 4040
rect 0 3982 1367 3984
rect 0 3952 800 3982
rect 1301 3979 1367 3982
rect 1577 4042 1643 4045
rect 18781 4042 18847 4045
rect 19517 4042 19583 4045
rect 1577 4040 12450 4042
rect 1577 3984 1582 4040
rect 1638 3984 12450 4040
rect 1577 3982 12450 3984
rect 1577 3979 1643 3982
rect 4429 3906 4495 3909
rect 4838 3906 4844 3908
rect 4429 3904 4844 3906
rect 4429 3848 4434 3904
rect 4490 3848 4844 3904
rect 4429 3846 4844 3848
rect 4429 3843 4495 3846
rect 4838 3844 4844 3846
rect 4908 3844 4914 3908
rect 4981 3906 5047 3909
rect 5758 3906 5764 3908
rect 4981 3904 5764 3906
rect 4981 3848 4986 3904
rect 5042 3848 5764 3904
rect 4981 3846 5764 3848
rect 4981 3843 5047 3846
rect 5758 3844 5764 3846
rect 5828 3844 5834 3908
rect 12014 3906 12020 3908
rect 9630 3846 12020 3906
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 4981 3770 5047 3773
rect 5717 3770 5783 3773
rect 4981 3768 5783 3770
rect 4981 3712 4986 3768
rect 5042 3712 5722 3768
rect 5778 3712 5783 3768
rect 4981 3710 5783 3712
rect 4981 3707 5047 3710
rect 5717 3707 5783 3710
rect 0 3634 800 3664
rect 1393 3634 1459 3637
rect 0 3632 1459 3634
rect 0 3576 1398 3632
rect 1454 3576 1459 3632
rect 0 3574 1459 3576
rect 0 3544 800 3574
rect 1393 3571 1459 3574
rect 3785 3634 3851 3637
rect 4705 3634 4771 3637
rect 3785 3632 4771 3634
rect 3785 3576 3790 3632
rect 3846 3576 4710 3632
rect 4766 3576 4771 3632
rect 3785 3574 4771 3576
rect 3785 3571 3851 3574
rect 4705 3571 4771 3574
rect 2497 3498 2563 3501
rect 9630 3498 9690 3846
rect 12014 3844 12020 3846
rect 12084 3906 12090 3908
rect 12157 3906 12223 3909
rect 12084 3904 12223 3906
rect 12084 3848 12162 3904
rect 12218 3848 12223 3904
rect 12084 3846 12223 3848
rect 12390 3906 12450 3982
rect 18781 4040 19583 4042
rect 18781 3984 18786 4040
rect 18842 3984 19522 4040
rect 19578 3984 19583 4040
rect 18781 3982 19583 3984
rect 18781 3979 18847 3982
rect 19517 3979 19583 3982
rect 21265 4042 21331 4045
rect 22200 4042 23000 4072
rect 21265 4040 23000 4042
rect 21265 3984 21270 4040
rect 21326 3984 23000 4040
rect 21265 3982 23000 3984
rect 21265 3979 21331 3982
rect 22200 3952 23000 3982
rect 13302 3906 13308 3908
rect 12390 3846 13308 3906
rect 12084 3844 12090 3846
rect 12157 3843 12223 3846
rect 13302 3844 13308 3846
rect 13372 3844 13378 3908
rect 15745 3906 15811 3909
rect 19517 3906 19583 3909
rect 15745 3904 19583 3906
rect 15745 3848 15750 3904
rect 15806 3848 19522 3904
rect 19578 3848 19583 3904
rect 15745 3846 19583 3848
rect 15745 3843 15811 3846
rect 19517 3843 19583 3846
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 11094 3708 11100 3772
rect 11164 3770 11170 3772
rect 12433 3770 12499 3773
rect 11164 3768 12499 3770
rect 11164 3712 12438 3768
rect 12494 3712 12499 3768
rect 11164 3710 12499 3712
rect 11164 3708 11170 3710
rect 12433 3707 12499 3710
rect 11145 3634 11211 3637
rect 15377 3634 15443 3637
rect 11145 3632 15443 3634
rect 11145 3576 11150 3632
rect 11206 3576 15382 3632
rect 15438 3576 15443 3632
rect 11145 3574 15443 3576
rect 11145 3571 11211 3574
rect 15377 3571 15443 3574
rect 21541 3634 21607 3637
rect 22200 3634 23000 3664
rect 21541 3632 23000 3634
rect 21541 3576 21546 3632
rect 21602 3576 23000 3632
rect 21541 3574 23000 3576
rect 21541 3571 21607 3574
rect 22200 3544 23000 3574
rect 10041 3500 10107 3501
rect 9990 3498 9996 3500
rect 2497 3496 9690 3498
rect 2497 3440 2502 3496
rect 2558 3440 9690 3496
rect 2497 3438 9690 3440
rect 9950 3438 9996 3498
rect 10060 3496 10107 3500
rect 11053 3498 11119 3501
rect 10102 3440 10107 3496
rect 2497 3435 2563 3438
rect 9990 3436 9996 3438
rect 10060 3436 10107 3440
rect 10041 3435 10107 3436
rect 10550 3496 11119 3498
rect 10550 3440 11058 3496
rect 11114 3440 11119 3496
rect 10550 3438 11119 3440
rect 5349 3362 5415 3365
rect 7465 3362 7531 3365
rect 10550 3362 10610 3438
rect 11053 3435 11119 3438
rect 5349 3360 10610 3362
rect 5349 3304 5354 3360
rect 5410 3304 7470 3360
rect 7526 3304 10610 3360
rect 5349 3302 10610 3304
rect 5349 3299 5415 3302
rect 7465 3299 7531 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 9765 3226 9831 3229
rect 10174 3226 10180 3228
rect 9765 3224 10180 3226
rect 9765 3168 9770 3224
rect 9826 3168 10180 3224
rect 9765 3166 10180 3168
rect 9765 3163 9831 3166
rect 10174 3164 10180 3166
rect 10244 3164 10250 3228
rect 0 3090 800 3120
rect 1761 3090 1827 3093
rect 0 3088 1827 3090
rect 0 3032 1766 3088
rect 1822 3032 1827 3088
rect 0 3030 1827 3032
rect 0 3000 800 3030
rect 1761 3027 1827 3030
rect 2037 3090 2103 3093
rect 7557 3090 7623 3093
rect 9622 3090 9628 3092
rect 2037 3088 9628 3090
rect 2037 3032 2042 3088
rect 2098 3032 7562 3088
rect 7618 3032 9628 3088
rect 2037 3030 9628 3032
rect 2037 3027 2103 3030
rect 7557 3027 7623 3030
rect 9622 3028 9628 3030
rect 9692 3028 9698 3092
rect 10910 3028 10916 3092
rect 10980 3090 10986 3092
rect 11329 3090 11395 3093
rect 10980 3088 11395 3090
rect 10980 3032 11334 3088
rect 11390 3032 11395 3088
rect 10980 3030 11395 3032
rect 10980 3028 10986 3030
rect 11329 3027 11395 3030
rect 11881 3090 11947 3093
rect 20897 3090 20963 3093
rect 11881 3088 20963 3090
rect 11881 3032 11886 3088
rect 11942 3032 20902 3088
rect 20958 3032 20963 3088
rect 11881 3030 20963 3032
rect 11881 3027 11947 3030
rect 20897 3027 20963 3030
rect 21173 3090 21239 3093
rect 22200 3090 23000 3120
rect 21173 3088 23000 3090
rect 21173 3032 21178 3088
rect 21234 3032 23000 3088
rect 21173 3030 23000 3032
rect 21173 3027 21239 3030
rect 22200 3000 23000 3030
rect 3233 2954 3299 2957
rect 8661 2954 8727 2957
rect 3233 2952 8727 2954
rect 3233 2896 3238 2952
rect 3294 2896 8666 2952
rect 8722 2896 8727 2952
rect 3233 2894 8727 2896
rect 3233 2891 3299 2894
rect 8661 2891 8727 2894
rect 10317 2954 10383 2957
rect 12934 2954 12940 2956
rect 10317 2952 12940 2954
rect 10317 2896 10322 2952
rect 10378 2896 12940 2952
rect 10317 2894 12940 2896
rect 10317 2891 10383 2894
rect 12934 2892 12940 2894
rect 13004 2954 13010 2956
rect 15377 2954 15443 2957
rect 13004 2952 15443 2954
rect 13004 2896 15382 2952
rect 15438 2896 15443 2952
rect 13004 2894 15443 2896
rect 13004 2892 13010 2894
rect 15377 2891 15443 2894
rect 17861 2954 17927 2957
rect 19425 2954 19491 2957
rect 17861 2952 19491 2954
rect 17861 2896 17866 2952
rect 17922 2896 19430 2952
rect 19486 2896 19491 2952
rect 17861 2894 19491 2896
rect 17861 2891 17927 2894
rect 19425 2891 19491 2894
rect 2405 2818 2471 2821
rect 5349 2818 5415 2821
rect 2405 2816 5415 2818
rect 2405 2760 2410 2816
rect 2466 2760 5354 2816
rect 5410 2760 5415 2816
rect 2405 2758 5415 2760
rect 2405 2755 2471 2758
rect 5349 2755 5415 2758
rect 6177 2818 6243 2821
rect 6494 2818 6500 2820
rect 6177 2816 6500 2818
rect 6177 2760 6182 2816
rect 6238 2760 6500 2816
rect 6177 2758 6500 2760
rect 6177 2755 6243 2758
rect 6494 2756 6500 2758
rect 6564 2756 6570 2820
rect 6729 2818 6795 2821
rect 6862 2818 6868 2820
rect 6729 2816 6868 2818
rect 6729 2760 6734 2816
rect 6790 2760 6868 2816
rect 6729 2758 6868 2760
rect 6729 2755 6795 2758
rect 6862 2756 6868 2758
rect 6932 2756 6938 2820
rect 9438 2756 9444 2820
rect 9508 2818 9514 2820
rect 9673 2818 9739 2821
rect 9508 2816 9739 2818
rect 9508 2760 9678 2816
rect 9734 2760 9739 2816
rect 9508 2758 9739 2760
rect 9508 2756 9514 2758
rect 9673 2755 9739 2758
rect 12985 2818 13051 2821
rect 13629 2818 13695 2821
rect 12985 2816 13695 2818
rect 12985 2760 12990 2816
rect 13046 2760 13634 2816
rect 13690 2760 13695 2816
rect 12985 2758 13695 2760
rect 12985 2755 13051 2758
rect 13629 2755 13695 2758
rect 14222 2756 14228 2820
rect 14292 2818 14298 2820
rect 14365 2818 14431 2821
rect 14292 2816 14431 2818
rect 14292 2760 14370 2816
rect 14426 2760 14431 2816
rect 14292 2758 14431 2760
rect 14292 2756 14298 2758
rect 14365 2755 14431 2758
rect 18505 2818 18571 2821
rect 18822 2818 18828 2820
rect 18505 2816 18828 2818
rect 18505 2760 18510 2816
rect 18566 2760 18828 2816
rect 18505 2758 18828 2760
rect 18505 2755 18571 2758
rect 18822 2756 18828 2758
rect 18892 2756 18898 2820
rect 20161 2818 20227 2821
rect 20118 2816 20227 2818
rect 20118 2760 20166 2816
rect 20222 2760 20227 2816
rect 20118 2755 20227 2760
rect 7874 2752 8194 2753
rect 0 2682 800 2712
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 12801 2684 12867 2685
rect 6494 2682 6500 2684
rect 0 2622 6500 2682
rect 0 2592 800 2622
rect 6494 2620 6500 2622
rect 6564 2620 6570 2684
rect 12750 2620 12756 2684
rect 12820 2682 12867 2684
rect 19241 2682 19307 2685
rect 20118 2682 20178 2755
rect 22200 2682 23000 2712
rect 12820 2680 12912 2682
rect 12862 2624 12912 2680
rect 12820 2622 12912 2624
rect 19241 2680 23000 2682
rect 19241 2624 19246 2680
rect 19302 2624 23000 2680
rect 19241 2622 23000 2624
rect 12820 2620 12867 2622
rect 12801 2619 12867 2620
rect 19241 2619 19307 2622
rect 22200 2592 23000 2622
rect 7189 2546 7255 2549
rect 10501 2548 10567 2549
rect 8518 2546 8524 2548
rect 7189 2544 8524 2546
rect 7189 2488 7194 2544
rect 7250 2488 8524 2544
rect 7189 2486 8524 2488
rect 7189 2483 7255 2486
rect 8518 2484 8524 2486
rect 8588 2484 8594 2548
rect 10501 2546 10548 2548
rect 10420 2544 10548 2546
rect 10612 2546 10618 2548
rect 17033 2546 17099 2549
rect 10612 2544 17099 2546
rect 10420 2488 10506 2544
rect 10612 2488 17038 2544
rect 17094 2488 17099 2544
rect 10420 2486 10548 2488
rect 10501 2484 10548 2486
rect 10612 2486 17099 2488
rect 10612 2484 10618 2486
rect 10501 2483 10567 2484
rect 17033 2483 17099 2486
rect 18689 2546 18755 2549
rect 20437 2546 20503 2549
rect 18689 2544 20503 2546
rect 18689 2488 18694 2544
rect 18750 2488 20442 2544
rect 20498 2488 20503 2544
rect 18689 2486 20503 2488
rect 18689 2483 18755 2486
rect 20437 2483 20503 2486
rect 5533 2410 5599 2413
rect 4156 2408 5599 2410
rect 4156 2352 5538 2408
rect 5594 2352 5599 2408
rect 4156 2350 5599 2352
rect 0 2274 800 2304
rect 4156 2274 4216 2350
rect 5533 2347 5599 2350
rect 0 2214 4216 2274
rect 4797 2274 4863 2277
rect 9581 2274 9647 2277
rect 4797 2272 9647 2274
rect 4797 2216 4802 2272
rect 4858 2216 9586 2272
rect 9642 2216 9647 2272
rect 4797 2214 9647 2216
rect 0 2184 800 2214
rect 4797 2211 4863 2214
rect 9581 2211 9647 2214
rect 18965 2274 19031 2277
rect 21725 2274 21791 2277
rect 22200 2274 23000 2304
rect 18965 2272 23000 2274
rect 18965 2216 18970 2272
rect 19026 2216 21730 2272
rect 21786 2216 23000 2272
rect 18965 2214 23000 2216
rect 18965 2211 19031 2214
rect 21725 2211 21791 2214
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 22200 2184 23000 2214
rect 18270 2143 18590 2144
rect 0 1866 800 1896
rect 933 1866 999 1869
rect 0 1864 999 1866
rect 0 1808 938 1864
rect 994 1808 999 1864
rect 0 1806 999 1808
rect 0 1776 800 1806
rect 933 1803 999 1806
rect 21541 1866 21607 1869
rect 22200 1866 23000 1896
rect 21541 1864 23000 1866
rect 21541 1808 21546 1864
rect 21602 1808 23000 1864
rect 21541 1806 23000 1808
rect 21541 1803 21607 1806
rect 22200 1776 23000 1806
rect 0 1458 800 1488
rect 4245 1458 4311 1461
rect 0 1456 4311 1458
rect 0 1400 4250 1456
rect 4306 1400 4311 1456
rect 0 1398 4311 1400
rect 0 1368 800 1398
rect 4245 1395 4311 1398
rect 20437 1458 20503 1461
rect 22200 1458 23000 1488
rect 20437 1456 23000 1458
rect 20437 1400 20442 1456
rect 20498 1400 23000 1456
rect 20437 1398 23000 1400
rect 20437 1395 20503 1398
rect 22200 1368 23000 1398
rect 18781 1322 18847 1325
rect 20713 1322 20779 1325
rect 18781 1320 20779 1322
rect 18781 1264 18786 1320
rect 18842 1264 20718 1320
rect 20774 1264 20779 1320
rect 18781 1262 20779 1264
rect 18781 1259 18847 1262
rect 20713 1259 20779 1262
rect 0 1050 800 1080
rect 1117 1050 1183 1053
rect 0 1048 1183 1050
rect 0 992 1122 1048
rect 1178 992 1183 1048
rect 0 990 1183 992
rect 0 960 800 990
rect 1117 987 1183 990
rect 21817 1050 21883 1053
rect 22200 1050 23000 1080
rect 21817 1048 23000 1050
rect 21817 992 21822 1048
rect 21878 992 23000 1048
rect 21817 990 23000 992
rect 21817 987 21883 990
rect 22200 960 23000 990
rect 0 642 800 672
rect 2957 642 3023 645
rect 0 640 3023 642
rect 0 584 2962 640
rect 3018 584 3023 640
rect 0 582 3023 584
rect 0 552 800 582
rect 2957 579 3023 582
rect 20713 642 20779 645
rect 22200 642 23000 672
rect 20713 640 23000 642
rect 20713 584 20718 640
rect 20774 584 23000 640
rect 20713 582 23000 584
rect 20713 579 20779 582
rect 22200 552 23000 582
rect 0 234 800 264
rect 1301 234 1367 237
rect 0 232 1367 234
rect 0 176 1306 232
rect 1362 176 1367 232
rect 0 174 1367 176
rect 0 144 800 174
rect 1301 171 1367 174
rect 22001 234 22067 237
rect 22200 234 23000 264
rect 22001 232 23000 234
rect 22001 176 22006 232
rect 22062 176 23000 232
rect 22001 174 23000 176
rect 22001 171 22067 174
rect 22200 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7236 19076 7300 19140
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 10548 17716 10612 17780
rect 8524 17504 8588 17508
rect 8524 17448 8574 17504
rect 8574 17448 8588 17504
rect 8524 17444 8588 17448
rect 9996 17444 10060 17508
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 6868 17172 6932 17236
rect 5948 16900 6012 16964
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 12572 16764 12636 16828
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 8708 16084 8772 16148
rect 9260 15812 9324 15876
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 11836 15328 11900 15332
rect 11836 15272 11886 15328
rect 11886 15272 11900 15328
rect 11836 15268 11900 15272
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 12020 15192 12084 15196
rect 12020 15136 12034 15192
rect 12034 15136 12084 15192
rect 12020 15132 12084 15136
rect 10180 14724 10244 14788
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 6684 14452 6748 14516
rect 4844 14180 4908 14244
rect 8892 14180 8956 14244
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 12388 14044 12452 14108
rect 5948 13908 6012 13972
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 5948 13424 6012 13428
rect 5948 13368 5962 13424
rect 5962 13368 6012 13424
rect 5948 13364 6012 13368
rect 10548 13908 10612 13972
rect 9812 13696 9876 13700
rect 9812 13640 9862 13696
rect 9862 13640 9876 13696
rect 9812 13636 9876 13640
rect 14596 13636 14660 13700
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 14228 13092 14292 13156
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 9076 13016 9140 13020
rect 9076 12960 9126 13016
rect 9126 12960 9140 13016
rect 9076 12956 9140 12960
rect 10916 12880 10980 12884
rect 10916 12824 10966 12880
rect 10966 12824 10980 12880
rect 10916 12820 10980 12824
rect 6684 12744 6748 12748
rect 6684 12688 6698 12744
rect 6698 12688 6748 12744
rect 6684 12684 6748 12688
rect 8340 12684 8404 12748
rect 10364 12684 10428 12748
rect 9444 12548 9508 12612
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 6684 12412 6748 12476
rect 5580 12336 5644 12340
rect 5580 12280 5594 12336
rect 5594 12280 5644 12336
rect 5580 12276 5644 12280
rect 5764 12276 5828 12340
rect 6684 12336 6748 12340
rect 6684 12280 6734 12336
rect 6734 12280 6748 12336
rect 6684 12276 6748 12280
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 9076 12276 9140 12340
rect 9812 12276 9876 12340
rect 12388 12276 12452 12340
rect 12756 12140 12820 12204
rect 10364 12064 10428 12068
rect 10364 12008 10414 12064
rect 10414 12008 10428 12064
rect 10364 12004 10428 12008
rect 10916 12004 10980 12068
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 9996 11596 10060 11660
rect 7420 11520 7484 11524
rect 7420 11464 7434 11520
rect 7434 11464 7484 11520
rect 7420 11460 7484 11464
rect 9628 11520 9692 11524
rect 9628 11464 9678 11520
rect 9678 11464 9692 11520
rect 9628 11460 9692 11464
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 9628 10916 9692 10980
rect 10180 10916 10244 10980
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 6684 10780 6748 10844
rect 4844 10644 4908 10708
rect 5580 10704 5644 10708
rect 5580 10648 5630 10704
rect 5630 10648 5644 10704
rect 5580 10644 5644 10648
rect 7052 10644 7116 10708
rect 7236 10372 7300 10436
rect 7604 10432 7668 10436
rect 7604 10376 7618 10432
rect 7618 10376 7668 10432
rect 7604 10372 7668 10376
rect 9812 10372 9876 10436
rect 11836 10372 11900 10436
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 8708 9964 8772 10028
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 8524 9692 8588 9756
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 6500 9556 6564 9620
rect 9812 9556 9876 9620
rect 20484 9556 20548 9620
rect 5764 9420 5828 9484
rect 7236 9420 7300 9484
rect 10180 9420 10244 9484
rect 3004 9148 3068 9212
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 9260 9148 9324 9212
rect 12204 9148 12268 9212
rect 13124 9148 13188 9212
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 10364 8740 10428 8804
rect 12572 8740 12636 8804
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 10732 8604 10796 8668
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 12940 8604 13004 8668
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14228 8196 14292 8260
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 8708 8060 8772 8124
rect 14412 8060 14476 8124
rect 9076 7924 9140 7988
rect 9444 7788 9508 7852
rect 9628 7788 9692 7852
rect 9260 7652 9324 7716
rect 10548 7712 10612 7716
rect 10548 7656 10598 7712
rect 10598 7656 10612 7712
rect 10548 7652 10612 7656
rect 10916 7652 10980 7716
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 6868 7576 6932 7580
rect 6868 7520 6918 7576
rect 6918 7520 6932 7576
rect 6868 7516 6932 7520
rect 13308 7576 13372 7580
rect 13308 7520 13358 7576
rect 13358 7520 13372 7576
rect 13308 7516 13372 7520
rect 14596 7516 14660 7580
rect 3924 7380 3988 7444
rect 8524 7380 8588 7444
rect 12204 7244 12268 7308
rect 9628 7108 9692 7172
rect 9812 7108 9876 7172
rect 12204 7108 12268 7172
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4844 6836 4908 6900
rect 6500 6836 6564 6900
rect 10180 6836 10244 6900
rect 11836 6836 11900 6900
rect 10180 6700 10244 6764
rect 9444 6624 9508 6628
rect 9444 6568 9458 6624
rect 9458 6568 9508 6624
rect 9444 6564 9508 6568
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 8892 6352 8956 6356
rect 8892 6296 8942 6352
rect 8942 6296 8956 6352
rect 8892 6292 8956 6296
rect 10364 6292 10428 6356
rect 9996 6156 10060 6220
rect 10180 6156 10244 6220
rect 12204 6156 12268 6220
rect 18828 6216 18892 6220
rect 18828 6160 18842 6216
rect 18842 6160 18892 6216
rect 18828 6156 18892 6160
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 12020 5884 12084 5948
rect 12388 5944 12452 5948
rect 12388 5888 12402 5944
rect 12402 5888 12452 5944
rect 12388 5884 12452 5888
rect 11100 5748 11164 5812
rect 11836 5748 11900 5812
rect 20484 5748 20548 5812
rect 3004 5612 3068 5676
rect 7420 5612 7484 5676
rect 9812 5476 9876 5540
rect 10732 5536 10796 5540
rect 10732 5480 10782 5536
rect 10782 5480 10796 5536
rect 10732 5476 10796 5480
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 3924 5340 3988 5404
rect 6684 5400 6748 5404
rect 6684 5344 6734 5400
rect 6734 5344 6748 5400
rect 6684 5340 6748 5344
rect 7236 5340 7300 5404
rect 8524 5204 8588 5268
rect 13124 4992 13188 4996
rect 13124 4936 13174 4992
rect 13174 4936 13188 4992
rect 13124 4932 13188 4936
rect 14412 4992 14476 4996
rect 14412 4936 14426 4992
rect 14426 4936 14476 4992
rect 14412 4932 14476 4936
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 7052 4720 7116 4724
rect 7052 4664 7066 4720
rect 7066 4664 7116 4720
rect 7052 4660 7116 4664
rect 11836 4796 11900 4860
rect 12572 4660 12636 4724
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7604 4252 7668 4316
rect 4844 3844 4908 3908
rect 5764 3844 5828 3908
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 12020 3844 12084 3908
rect 13308 3844 13372 3908
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 11100 3708 11164 3772
rect 9996 3496 10060 3500
rect 9996 3440 10046 3496
rect 10046 3440 10060 3496
rect 9996 3436 10060 3440
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 10180 3164 10244 3228
rect 9628 3028 9692 3092
rect 10916 3028 10980 3092
rect 12940 2892 13004 2956
rect 6500 2756 6564 2820
rect 6868 2756 6932 2820
rect 9444 2756 9508 2820
rect 14228 2756 14292 2820
rect 18828 2756 18892 2820
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 6500 2620 6564 2684
rect 12756 2680 12820 2684
rect 12756 2624 12806 2680
rect 12806 2624 12820 2680
rect 12756 2620 12820 2624
rect 8524 2484 8588 2548
rect 10548 2544 10612 2548
rect 10548 2488 10562 2544
rect 10562 2488 10612 2544
rect 10548 2484 10612 2488
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7235 19140 7301 19141
rect 7235 19076 7236 19140
rect 7300 19076 7301 19140
rect 7235 19075 7301 19076
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 6867 17236 6933 17237
rect 6867 17172 6868 17236
rect 6932 17172 6933 17236
rect 6867 17171 6933 17172
rect 5947 16964 6013 16965
rect 5947 16900 5948 16964
rect 6012 16900 6013 16964
rect 5947 16899 6013 16900
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4843 14244 4909 14245
rect 4843 14180 4844 14244
rect 4908 14180 4909 14244
rect 4843 14179 4909 14180
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4846 10709 4906 14179
rect 5950 13973 6010 16899
rect 6683 14516 6749 14517
rect 6683 14452 6684 14516
rect 6748 14452 6749 14516
rect 6683 14451 6749 14452
rect 5947 13972 6013 13973
rect 5947 13908 5948 13972
rect 6012 13908 6013 13972
rect 5947 13907 6013 13908
rect 5950 13429 6010 13907
rect 5947 13428 6013 13429
rect 5947 13364 5948 13428
rect 6012 13364 6013 13428
rect 5947 13363 6013 13364
rect 6686 12749 6746 14451
rect 6683 12748 6749 12749
rect 6683 12684 6684 12748
rect 6748 12684 6749 12748
rect 6683 12683 6749 12684
rect 6683 12476 6749 12477
rect 6683 12412 6684 12476
rect 6748 12412 6749 12476
rect 6683 12411 6749 12412
rect 6686 12341 6746 12411
rect 5579 12340 5645 12341
rect 5579 12276 5580 12340
rect 5644 12276 5645 12340
rect 5579 12275 5645 12276
rect 5763 12340 5829 12341
rect 5763 12276 5764 12340
rect 5828 12276 5829 12340
rect 5763 12275 5829 12276
rect 6683 12340 6749 12341
rect 6683 12276 6684 12340
rect 6748 12276 6749 12340
rect 6683 12275 6749 12276
rect 5582 10709 5642 12275
rect 4843 10708 4909 10709
rect 4843 10644 4844 10708
rect 4908 10644 4909 10708
rect 4843 10643 4909 10644
rect 5579 10708 5645 10709
rect 5579 10644 5580 10708
rect 5644 10644 5645 10708
rect 5579 10643 5645 10644
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 3003 9212 3069 9213
rect 3003 9148 3004 9212
rect 3068 9148 3069 9212
rect 3003 9147 3069 9148
rect 3006 5677 3066 9147
rect 4409 8736 4729 9760
rect 5766 9485 5826 12275
rect 6683 10844 6749 10845
rect 6683 10780 6684 10844
rect 6748 10780 6749 10844
rect 6683 10779 6749 10780
rect 6499 9620 6565 9621
rect 6499 9556 6500 9620
rect 6564 9556 6565 9620
rect 6499 9555 6565 9556
rect 5763 9484 5829 9485
rect 5763 9420 5764 9484
rect 5828 9420 5829 9484
rect 5763 9419 5829 9420
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 3923 7444 3989 7445
rect 3923 7380 3924 7444
rect 3988 7380 3989 7444
rect 3923 7379 3989 7380
rect 3003 5676 3069 5677
rect 3003 5612 3004 5676
rect 3068 5612 3069 5676
rect 3003 5611 3069 5612
rect 3926 5405 3986 7379
rect 4409 6560 4729 7584
rect 4843 6900 4909 6901
rect 4843 6836 4844 6900
rect 4908 6836 4909 6900
rect 4843 6835 4909 6836
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 3923 5404 3989 5405
rect 3923 5340 3924 5404
rect 3988 5340 3989 5404
rect 3923 5339 3989 5340
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4846 3909 4906 6835
rect 5766 3909 5826 9419
rect 6502 6901 6562 9555
rect 6499 6900 6565 6901
rect 6499 6836 6500 6900
rect 6564 6836 6565 6900
rect 6499 6835 6565 6836
rect 6686 5405 6746 10779
rect 6870 7581 6930 17171
rect 7051 10708 7117 10709
rect 7051 10644 7052 10708
rect 7116 10644 7117 10708
rect 7051 10643 7117 10644
rect 6867 7580 6933 7581
rect 6867 7516 6868 7580
rect 6932 7516 6933 7580
rect 6867 7515 6933 7516
rect 6683 5404 6749 5405
rect 6683 5340 6684 5404
rect 6748 5340 6749 5404
rect 6683 5339 6749 5340
rect 4843 3908 4909 3909
rect 4843 3844 4844 3908
rect 4908 3844 4909 3908
rect 4843 3843 4909 3844
rect 5763 3908 5829 3909
rect 5763 3844 5764 3908
rect 5828 3844 5829 3908
rect 5763 3843 5829 3844
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 6870 2821 6930 7515
rect 7054 4725 7114 10643
rect 7238 10437 7298 19075
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 10547 17780 10613 17781
rect 10547 17716 10548 17780
rect 10612 17716 10613 17780
rect 10547 17715 10613 17716
rect 8523 17508 8589 17509
rect 8523 17444 8524 17508
rect 8588 17444 8589 17508
rect 8523 17443 8589 17444
rect 9995 17508 10061 17509
rect 9995 17444 9996 17508
rect 10060 17444 10061 17508
rect 9995 17443 10061 17444
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 8339 12748 8405 12749
rect 8339 12684 8340 12748
rect 8404 12684 8405 12748
rect 8339 12683 8405 12684
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7419 11524 7485 11525
rect 7419 11460 7420 11524
rect 7484 11460 7485 11524
rect 7419 11459 7485 11460
rect 7235 10436 7301 10437
rect 7235 10372 7236 10436
rect 7300 10372 7301 10436
rect 7235 10371 7301 10372
rect 7235 9484 7301 9485
rect 7235 9420 7236 9484
rect 7300 9420 7301 9484
rect 7235 9419 7301 9420
rect 7238 5405 7298 9419
rect 7422 5677 7482 11459
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7603 10436 7669 10437
rect 7603 10372 7604 10436
rect 7668 10372 7669 10436
rect 7603 10371 7669 10372
rect 7419 5676 7485 5677
rect 7419 5612 7420 5676
rect 7484 5612 7485 5676
rect 7419 5611 7485 5612
rect 7235 5404 7301 5405
rect 7235 5340 7236 5404
rect 7300 5340 7301 5404
rect 7235 5339 7301 5340
rect 7051 4724 7117 4725
rect 7051 4660 7052 4724
rect 7116 4660 7117 4724
rect 7051 4659 7117 4660
rect 7606 4317 7666 10371
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 8342 7850 8402 12683
rect 8526 9757 8586 17443
rect 8707 16148 8773 16149
rect 8707 16084 8708 16148
rect 8772 16084 8773 16148
rect 8707 16083 8773 16084
rect 8710 10029 8770 16083
rect 9259 15876 9325 15877
rect 9259 15812 9260 15876
rect 9324 15812 9325 15876
rect 9259 15811 9325 15812
rect 8891 14244 8957 14245
rect 8891 14180 8892 14244
rect 8956 14180 8957 14244
rect 8891 14179 8957 14180
rect 8707 10028 8773 10029
rect 8707 9964 8708 10028
rect 8772 9964 8773 10028
rect 8707 9963 8773 9964
rect 8523 9756 8589 9757
rect 8523 9692 8524 9756
rect 8588 9692 8589 9756
rect 8523 9691 8589 9692
rect 8707 8124 8773 8125
rect 8707 8060 8708 8124
rect 8772 8060 8773 8124
rect 8707 8059 8773 8060
rect 8710 7850 8770 8059
rect 8342 7790 8770 7850
rect 8526 7445 8586 7790
rect 8523 7444 8589 7445
rect 8523 7380 8524 7444
rect 8588 7380 8589 7444
rect 8523 7379 8589 7380
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 8894 6357 8954 14179
rect 9075 13020 9141 13021
rect 9075 12956 9076 13020
rect 9140 12956 9141 13020
rect 9075 12955 9141 12956
rect 9078 12341 9138 12955
rect 9075 12340 9141 12341
rect 9075 12276 9076 12340
rect 9140 12276 9141 12340
rect 9075 12275 9141 12276
rect 9262 9482 9322 15811
rect 9811 13700 9877 13701
rect 9811 13636 9812 13700
rect 9876 13636 9877 13700
rect 9811 13635 9877 13636
rect 9443 12612 9509 12613
rect 9443 12548 9444 12612
rect 9508 12548 9509 12612
rect 9443 12547 9509 12548
rect 9078 9422 9322 9482
rect 9078 7989 9138 9422
rect 9259 9212 9325 9213
rect 9259 9148 9260 9212
rect 9324 9148 9325 9212
rect 9259 9147 9325 9148
rect 9075 7988 9141 7989
rect 9075 7924 9076 7988
rect 9140 7924 9141 7988
rect 9075 7923 9141 7924
rect 9262 7717 9322 9147
rect 9446 7853 9506 12547
rect 9814 12341 9874 13635
rect 9811 12340 9877 12341
rect 9811 12276 9812 12340
rect 9876 12276 9877 12340
rect 9811 12275 9877 12276
rect 9627 11524 9693 11525
rect 9627 11460 9628 11524
rect 9692 11460 9693 11524
rect 9627 11459 9693 11460
rect 9630 10981 9690 11459
rect 9627 10980 9693 10981
rect 9627 10916 9628 10980
rect 9692 10916 9693 10980
rect 9627 10915 9693 10916
rect 9814 10437 9874 12275
rect 9998 11661 10058 17443
rect 10179 14788 10245 14789
rect 10179 14724 10180 14788
rect 10244 14724 10245 14788
rect 10179 14723 10245 14724
rect 9995 11660 10061 11661
rect 9995 11596 9996 11660
rect 10060 11596 10061 11660
rect 9995 11595 10061 11596
rect 10182 10981 10242 14723
rect 10550 13973 10610 17715
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 12571 16828 12637 16829
rect 12571 16764 12572 16828
rect 12636 16764 12637 16828
rect 12571 16763 12637 16764
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11835 15332 11901 15333
rect 11835 15268 11836 15332
rect 11900 15268 11901 15332
rect 11835 15267 11901 15268
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 10547 13972 10613 13973
rect 10547 13908 10548 13972
rect 10612 13908 10613 13972
rect 10547 13907 10613 13908
rect 10363 12748 10429 12749
rect 10363 12684 10364 12748
rect 10428 12684 10429 12748
rect 10363 12683 10429 12684
rect 10366 12069 10426 12683
rect 10363 12068 10429 12069
rect 10363 12004 10364 12068
rect 10428 12004 10429 12068
rect 10363 12003 10429 12004
rect 10179 10980 10245 10981
rect 10179 10916 10180 10980
rect 10244 10916 10245 10980
rect 10179 10915 10245 10916
rect 9811 10436 9877 10437
rect 9811 10372 9812 10436
rect 9876 10372 9877 10436
rect 9811 10371 9877 10372
rect 10550 9690 10610 13907
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 10915 12884 10981 12885
rect 10915 12820 10916 12884
rect 10980 12820 10981 12884
rect 10915 12819 10981 12820
rect 10918 12069 10978 12819
rect 10915 12068 10981 12069
rect 10915 12004 10916 12068
rect 10980 12004 10981 12068
rect 10915 12003 10981 12004
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11838 10437 11898 15267
rect 12019 15196 12085 15197
rect 12019 15132 12020 15196
rect 12084 15132 12085 15196
rect 12019 15131 12085 15132
rect 11835 10436 11901 10437
rect 11835 10372 11836 10436
rect 11900 10372 11901 10436
rect 11835 10371 11901 10372
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 10550 9630 11162 9690
rect 9811 9620 9877 9621
rect 9811 9556 9812 9620
rect 9876 9556 9877 9620
rect 9811 9555 9877 9556
rect 9443 7852 9509 7853
rect 9443 7788 9444 7852
rect 9508 7788 9509 7852
rect 9443 7787 9509 7788
rect 9627 7852 9693 7853
rect 9627 7788 9628 7852
rect 9692 7788 9693 7852
rect 9627 7787 9693 7788
rect 9259 7716 9325 7717
rect 9259 7652 9260 7716
rect 9324 7652 9325 7716
rect 9259 7651 9325 7652
rect 9262 6930 9322 7651
rect 9630 7173 9690 7787
rect 9814 7173 9874 9555
rect 10179 9484 10245 9485
rect 10179 9420 10180 9484
rect 10244 9420 10245 9484
rect 10179 9419 10245 9420
rect 9627 7172 9693 7173
rect 9627 7108 9628 7172
rect 9692 7108 9693 7172
rect 9627 7107 9693 7108
rect 9811 7172 9877 7173
rect 9811 7108 9812 7172
rect 9876 7108 9877 7172
rect 9811 7107 9877 7108
rect 9262 6870 9690 6930
rect 9443 6628 9509 6629
rect 9443 6564 9444 6628
rect 9508 6564 9509 6628
rect 9443 6563 9509 6564
rect 8891 6356 8957 6357
rect 8891 6292 8892 6356
rect 8956 6292 8957 6356
rect 8891 6291 8957 6292
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 8523 5268 8589 5269
rect 8523 5204 8524 5268
rect 8588 5204 8589 5268
rect 8523 5203 8589 5204
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7603 4316 7669 4317
rect 7603 4252 7604 4316
rect 7668 4252 7669 4316
rect 7603 4251 7669 4252
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 6499 2820 6565 2821
rect 6499 2756 6500 2820
rect 6564 2756 6565 2820
rect 6499 2755 6565 2756
rect 6867 2820 6933 2821
rect 6867 2756 6868 2820
rect 6932 2756 6933 2820
rect 6867 2755 6933 2756
rect 6502 2685 6562 2755
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 6499 2684 6565 2685
rect 6499 2620 6500 2684
rect 6564 2620 6565 2684
rect 6499 2619 6565 2620
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 2128 8195 2688
rect 8526 2549 8586 5203
rect 9446 2821 9506 6563
rect 9630 3093 9690 6870
rect 9814 5541 9874 7107
rect 10182 6901 10242 9419
rect 10363 8804 10429 8805
rect 10363 8740 10364 8804
rect 10428 8740 10429 8804
rect 10363 8739 10429 8740
rect 10179 6900 10245 6901
rect 10179 6836 10180 6900
rect 10244 6836 10245 6900
rect 10179 6835 10245 6836
rect 10179 6764 10245 6765
rect 10179 6700 10180 6764
rect 10244 6700 10245 6764
rect 10179 6699 10245 6700
rect 10182 6221 10242 6699
rect 10366 6357 10426 8739
rect 10731 8668 10797 8669
rect 10731 8604 10732 8668
rect 10796 8604 10797 8668
rect 10731 8603 10797 8604
rect 10547 7716 10613 7717
rect 10547 7652 10548 7716
rect 10612 7652 10613 7716
rect 10547 7651 10613 7652
rect 10363 6356 10429 6357
rect 10363 6292 10364 6356
rect 10428 6292 10429 6356
rect 10363 6291 10429 6292
rect 9995 6220 10061 6221
rect 9995 6156 9996 6220
rect 10060 6156 10061 6220
rect 9995 6155 10061 6156
rect 10179 6220 10245 6221
rect 10179 6156 10180 6220
rect 10244 6156 10245 6220
rect 10179 6155 10245 6156
rect 9811 5540 9877 5541
rect 9811 5476 9812 5540
rect 9876 5476 9877 5540
rect 9811 5475 9877 5476
rect 9998 3501 10058 6155
rect 9995 3500 10061 3501
rect 9995 3436 9996 3500
rect 10060 3436 10061 3500
rect 9995 3435 10061 3436
rect 10182 3229 10242 6155
rect 10179 3228 10245 3229
rect 10179 3164 10180 3228
rect 10244 3164 10245 3228
rect 10179 3163 10245 3164
rect 9627 3092 9693 3093
rect 9627 3028 9628 3092
rect 9692 3028 9693 3092
rect 9627 3027 9693 3028
rect 9443 2820 9509 2821
rect 9443 2756 9444 2820
rect 9508 2756 9509 2820
rect 9443 2755 9509 2756
rect 10550 2549 10610 7651
rect 10734 5541 10794 8603
rect 10915 7716 10981 7717
rect 10915 7652 10916 7716
rect 10980 7652 10981 7716
rect 10915 7651 10981 7652
rect 10731 5540 10797 5541
rect 10731 5476 10732 5540
rect 10796 5476 10797 5540
rect 10731 5475 10797 5476
rect 10918 3093 10978 7651
rect 11102 5813 11162 9630
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11835 6900 11901 6901
rect 11835 6836 11836 6900
rect 11900 6836 11901 6900
rect 11835 6835 11901 6836
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11099 5812 11165 5813
rect 11099 5748 11100 5812
rect 11164 5748 11165 5812
rect 11099 5747 11165 5748
rect 11102 3773 11162 5747
rect 11340 5472 11660 6496
rect 11838 5813 11898 6835
rect 12022 5949 12082 15131
rect 12387 14108 12453 14109
rect 12387 14044 12388 14108
rect 12452 14044 12453 14108
rect 12387 14043 12453 14044
rect 12390 12341 12450 14043
rect 12387 12340 12453 12341
rect 12387 12276 12388 12340
rect 12452 12276 12453 12340
rect 12387 12275 12453 12276
rect 12203 9212 12269 9213
rect 12203 9148 12204 9212
rect 12268 9148 12269 9212
rect 12203 9147 12269 9148
rect 12206 7309 12266 9147
rect 12203 7308 12269 7309
rect 12203 7244 12204 7308
rect 12268 7244 12269 7308
rect 12203 7243 12269 7244
rect 12203 7172 12269 7173
rect 12203 7108 12204 7172
rect 12268 7108 12269 7172
rect 12203 7107 12269 7108
rect 12206 6221 12266 7107
rect 12203 6220 12269 6221
rect 12203 6156 12204 6220
rect 12268 6156 12269 6220
rect 12203 6155 12269 6156
rect 12390 5949 12450 12275
rect 12574 8805 12634 16763
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14595 13700 14661 13701
rect 14595 13636 14596 13700
rect 14660 13636 14661 13700
rect 14595 13635 14661 13636
rect 14227 13156 14293 13157
rect 14227 13092 14228 13156
rect 14292 13092 14293 13156
rect 14227 13091 14293 13092
rect 12755 12204 12821 12205
rect 12755 12140 12756 12204
rect 12820 12140 12821 12204
rect 12755 12139 12821 12140
rect 12571 8804 12637 8805
rect 12571 8740 12572 8804
rect 12636 8740 12637 8804
rect 12571 8739 12637 8740
rect 12019 5948 12085 5949
rect 12019 5884 12020 5948
rect 12084 5884 12085 5948
rect 12019 5883 12085 5884
rect 12387 5948 12453 5949
rect 12387 5884 12388 5948
rect 12452 5884 12453 5948
rect 12387 5883 12453 5884
rect 11835 5812 11901 5813
rect 11835 5748 11836 5812
rect 11900 5748 11901 5812
rect 11835 5747 11901 5748
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11838 4861 11898 5747
rect 11835 4860 11901 4861
rect 11835 4796 11836 4860
rect 11900 4796 11901 4860
rect 11835 4795 11901 4796
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11099 3772 11165 3773
rect 11099 3708 11100 3772
rect 11164 3708 11165 3772
rect 11099 3707 11165 3708
rect 11340 3296 11660 4320
rect 12022 3909 12082 5883
rect 12574 4725 12634 8739
rect 12571 4724 12637 4725
rect 12571 4660 12572 4724
rect 12636 4660 12637 4724
rect 12571 4659 12637 4660
rect 12019 3908 12085 3909
rect 12019 3844 12020 3908
rect 12084 3844 12085 3908
rect 12019 3843 12085 3844
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 10915 3092 10981 3093
rect 10915 3028 10916 3092
rect 10980 3028 10981 3092
rect 10915 3027 10981 3028
rect 8523 2548 8589 2549
rect 8523 2484 8524 2548
rect 8588 2484 8589 2548
rect 8523 2483 8589 2484
rect 10547 2548 10613 2549
rect 10547 2484 10548 2548
rect 10612 2484 10613 2548
rect 10547 2483 10613 2484
rect 11340 2208 11660 3232
rect 12758 2685 12818 12139
rect 13123 9212 13189 9213
rect 13123 9148 13124 9212
rect 13188 9148 13189 9212
rect 13123 9147 13189 9148
rect 12939 8668 13005 8669
rect 12939 8604 12940 8668
rect 13004 8604 13005 8668
rect 12939 8603 13005 8604
rect 12942 2957 13002 8603
rect 13126 4997 13186 9147
rect 14230 8261 14290 13091
rect 14227 8260 14293 8261
rect 14227 8196 14228 8260
rect 14292 8196 14293 8260
rect 14227 8195 14293 8196
rect 13307 7580 13373 7581
rect 13307 7516 13308 7580
rect 13372 7516 13373 7580
rect 13307 7515 13373 7516
rect 13123 4996 13189 4997
rect 13123 4932 13124 4996
rect 13188 4932 13189 4996
rect 13123 4931 13189 4932
rect 13310 3909 13370 7515
rect 13307 3908 13373 3909
rect 13307 3844 13308 3908
rect 13372 3844 13373 3908
rect 13307 3843 13373 3844
rect 12939 2956 13005 2957
rect 12939 2892 12940 2956
rect 13004 2892 13005 2956
rect 12939 2891 13005 2892
rect 14230 2821 14290 8195
rect 14411 8124 14477 8125
rect 14411 8060 14412 8124
rect 14476 8060 14477 8124
rect 14411 8059 14477 8060
rect 14414 4997 14474 8059
rect 14598 7581 14658 13635
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14595 7580 14661 7581
rect 14595 7516 14596 7580
rect 14660 7516 14661 7580
rect 14595 7515 14661 7516
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14411 4996 14477 4997
rect 14411 4932 14412 4996
rect 14476 4932 14477 4996
rect 14411 4931 14477 4932
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14227 2820 14293 2821
rect 14227 2756 14228 2820
rect 14292 2756 14293 2820
rect 14227 2755 14293 2756
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 12755 2684 12821 2685
rect 12755 2620 12756 2684
rect 12820 2620 12821 2684
rect 12755 2619 12821 2620
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 20483 9620 20549 9621
rect 20483 9556 20484 9620
rect 20548 9556 20549 9620
rect 20483 9555 20549 9556
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18827 6220 18893 6221
rect 18827 6156 18828 6220
rect 18892 6156 18893 6220
rect 18827 6155 18893 6156
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18830 2821 18890 6155
rect 20486 5813 20546 9555
rect 20483 5812 20549 5813
rect 20483 5748 20484 5812
rect 20548 5748 20549 5812
rect 20483 5747 20549 5748
rect 18827 2820 18893 2821
rect 18827 2756 18828 2820
rect 18892 2756 18893 2820
rect 18827 2755 18893 2756
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1624635492
transform 1 0 1840 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1624635492
transform 1 0 1932 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform 1 0 1656 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1624635492
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2116 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 2668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output122 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1624635492
transform 1 0 2668 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1624635492
transform 1 0 2208 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1624635492
transform 1 0 2208 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2852 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_20
timestamp 1624635492
transform 1 0 2944 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3864 0 1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1624635492
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1624635492
transform 1 0 3036 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1624635492
transform 1 0 4876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28
timestamp 1624635492
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_47
timestamp 1624635492
transform 1 0 5428 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48
timestamp 1624635492
transform 1 0 5520 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1624635492
transform -1 0 5520 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1624635492
transform 1 0 5612 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1624635492
transform -1 0 6348 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1624635492
transform -1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 8280 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1624635492
transform 1 0 8464 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1624635492
transform 1 0 7268 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1624635492
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  input66 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 8464 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10856 0 1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1624635492
transform 1 0 10028 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1624635492
transform -1 0 10764 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1624635492
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 13156 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1624635492
transform 1 0 11868 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1624635492
transform -1 0 11776 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1624635492
transform -1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1624635492
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1624635492
transform -1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 13984 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1624635492
transform -1 0 14536 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1624635492
transform -1 0 14444 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1624635492
transform 1 0 13156 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1624635492
transform -1 0 13064 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1624635492
transform -1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1624635492
transform -1 0 13800 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output163
timestamp 1624635492
transform -1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output175
timestamp 1624635492
transform -1 0 15272 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output174
timestamp 1624635492
transform -1 0 14904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1624635492
transform -1 0 15088 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1624635492
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output176
timestamp 1624635492
transform -1 0 15640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1624635492
transform -1 0 15640 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1624635492
transform -1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output180
timestamp 1624635492
transform -1 0 16008 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output177
timestamp 1624635492
transform -1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output181
timestamp 1624635492
transform -1 0 16376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output178
timestamp 1624635492
transform -1 0 16376 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_166
timestamp 1624635492
transform 1 0 16376 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output179
timestamp 1624635492
transform -1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 16928 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1624635492
transform -1 0 18584 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output164
timestamp 1624635492
transform -1 0 17572 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output165
timestamp 1624635492
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output182
timestamp 1624635492
transform -1 0 16836 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1624635492
transform -1 0 17756 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1624635492
transform 1 0 18584 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1624635492
transform -1 0 19228 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1624635492
transform -1 0 19504 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_207
timestamp 1624635492
transform 1 0 20148 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output171
timestamp 1624635492
transform -1 0 20148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output167
timestamp 1624635492
transform -1 0 20240 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output166
timestamp 1624635492
transform -1 0 19780 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1624635492
transform -1 0 19780 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output172
timestamp 1624635492
transform -1 0 20608 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output168
timestamp 1624635492
transform -1 0 20608 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1624635492
transform 1 0 20976 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1624635492
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output169
timestamp 1624635492
transform -1 0 20976 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output170
timestamp 1624635492
transform -1 0 21344 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output173
timestamp 1624635492
transform -1 0 20976 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output207
timestamp 1624635492
transform 1 0 21252 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2944 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1624635492
transform 1 0 2116 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1624635492
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1624635492
transform 1 0 1656 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 2116 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5704 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1624635492
transform 1 0 4140 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 8188 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1624635492
transform -1 0 6716 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 5888 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1624635492
transform 1 0 8188 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 10948 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 12420 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1624635492
transform -1 0 13248 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1624635492
transform 1 0 13248 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1624635492
transform -1 0 14260 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1624635492
transform -1 0 15732 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1624635492
transform -1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 17572 0 -1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15456 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1624635492
transform -1 0 17848 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1624635492
transform -1 0 18124 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1624635492
transform -1 0 19136 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1624635492
transform -1 0 18308 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1624635492
transform -1 0 19412 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1624635492
transform 1 0 19596 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_199
timestamp 1624635492
transform 1 0 19412 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1624635492
transform -1 0 20700 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output211
timestamp 1624635492
transform 1 0 21252 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output221
timestamp 1624635492
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 4140 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1624635492
transform -1 0 2668 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 1840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1624635492
transform 1 0 4140 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1624635492
transform -1 0 4692 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1624635492
transform -1 0 6348 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1624635492
transform -1 0 6716 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp 1624635492
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1624635492
transform 1 0 8280 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9476 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1624635492
transform -1 0 10580 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1624635492
transform -1 0 10856 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1624635492
transform -1 0 9476 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11960 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1624635492
transform -1 0 12788 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1624635492
transform -1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1624635492
transform -1 0 11224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1624635492
transform -1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1624635492
transform -1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14628 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1624635492
transform 1 0 12788 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 13892 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1624635492
transform -1 0 14076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1624635492
transform -1 0 14260 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_143
timestamp 1624635492
transform 1 0 14260 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1624635492
transform -1 0 16560 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1624635492
transform -1 0 16192 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14904 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1624635492
transform -1 0 15732 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_164
timestamp 1624635492
transform 1 0 16192 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1624635492
transform -1 0 16836 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 19136 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 17204 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1624635492
transform -1 0 17664 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1624635492
transform -1 0 17480 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_175
timestamp 1624635492
transform 1 0 17204 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1624635492
transform 1 0 19964 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1624635492
transform 1 0 19136 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 1624635492
transform 1 0 20240 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1624635492
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1624635492
transform -1 0 21344 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input105
timestamp 1624635492
transform -1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input106
timestamp 1624635492
transform -1 0 20792 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 2852 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2944 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1624635492
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1624635492
transform 1 0 4692 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 7084 0 -1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1624635492
transform -1 0 9016 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1624635492
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1624635492
transform 1 0 7084 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11132 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1624635492
transform -1 0 10304 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 9384 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_90
timestamp 1624635492
transform 1 0 9384 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1624635492
transform 1 0 11132 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12328 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1624635492
transform -1 0 12604 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_118
timestamp 1624635492
transform 1 0 11960 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_125
timestamp 1624635492
transform 1 0 12604 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 14168 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1624635492
transform -1 0 14536 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_142
timestamp 1624635492
transform 1 0 14168 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1624635492
transform -1 0 15456 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 15548 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 15088 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1624635492
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_156
timestamp 1624635492
transform 1 0 15456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1624635492
transform -1 0 18860 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1624635492
transform -1 0 18032 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1624635492
transform -1 0 17204 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1624635492
transform 1 0 19596 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 19504 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 19320 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1624635492
transform -1 0 19136 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_193
timestamp 1624635492
transform 1 0 18860 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1624635492
transform -1 0 21620 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input107
timestamp 1624635492
transform -1 0 21252 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input109
timestamp 1624635492
transform -1 0 20976 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 1624635492
transform -1 0 20700 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 2668 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1624635492
transform 1 0 1840 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1624635492
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1624635492
transform 1 0 4140 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1624635492
transform -1 0 7636 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1624635492
transform 1 0 5428 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input95
timestamp 1624635492
transform -1 0 5244 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 5428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1624635492
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_61
timestamp 1624635492
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1624635492
transform 1 0 7636 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624635492
transform -1 0 8648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1624635492
transform -1 0 8832 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 10672 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1624635492
transform -1 0 11500 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1624635492
transform -1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1624635492
transform -1 0 9200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1624635492
transform -1 0 13340 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1624635492
transform 1 0 11500 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 13340 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1624635492
transform -1 0 14996 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 14996 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 18032 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1624635492
transform -1 0 17756 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1624635492
transform -1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A1
timestamp 1624635492
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 16836 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_181
timestamp 1624635492
transform 1 0 17756 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1624635492
transform -1 0 20332 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1624635492
transform -1 0 21620 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 1624635492
transform -1 0 21252 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input112
timestamp 1624635492
transform -1 0 20976 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output217
timestamp 1624635492
transform 1 0 20424 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_209
timestamp 1624635492
transform 1 0 20332 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1624635492
transform 1 0 2852 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 1748 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 2024 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1624635492
transform -1 0 2852 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 3312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1624635492
transform 1 0 3312 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1624635492
transform 1 0 3312 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 4600 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input96
timestamp 1624635492
transform 1 0 4140 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4600 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 4140 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6348 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5428 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 1624635492
transform -1 0 5888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input98
timestamp 1624635492
transform -1 0 6164 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 6348 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_56
timestamp 1624635492
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1624635492
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1624635492
transform 1 0 8372 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1624635492
transform 1 0 7728 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1624635492
transform -1 0 8096 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input101
timestamp 1624635492
transform -1 0 7452 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 7636 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1624635492
transform -1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_71
timestamp 1624635492
transform 1 0 7636 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_78
timestamp 1624635492
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10856 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1624635492
transform -1 0 11224 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1624635492
transform -1 0 10396 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1624635492
transform -1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1624635492
transform -1 0 9292 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1624635492
transform -1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1624635492
transform -1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_89
timestamp 1624635492
transform 1 0 9292 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10856 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 12052 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0
timestamp 1624635492
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1624635492
transform 1 0 11684 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 12236 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12512 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1624635492
transform 1 0 13064 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14996 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_141
timestamp 1624635492
transform 1 0 14076 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1624635492
transform -1 0 16652 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16468 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A0
timestamp 1624635492
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1624635492
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_155
timestamp 1624635492
transform 1 0 15364 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1624635492
transform 1 0 16468 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1624635492
transform -1 0 17480 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1624635492
transform -1 0 16836 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_181
timestamp 1624635492
transform 1 0 17756 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_178
timestamp 1624635492
transform 1 0 17480 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1624635492
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1624635492
transform -1 0 18584 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 19504 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_190
timestamp 1624635492
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1624635492
transform -1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1624635492
transform -1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 19780 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 19964 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 20148 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1624635492
transform 1 0 20148 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 19228 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20700 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1624635492
transform -1 0 21620 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1624635492
transform -1 0 21620 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1624635492
transform -1 0 21252 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1624635492
transform -1 0 21252 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 20884 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_214
timestamp 1624635492
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1624635492
transform 1 0 2760 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1624635492
transform -1 0 2760 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5336 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6072 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 1624635492
transform -1 0 5612 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input100
timestamp 1624635492
transform -1 0 5888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 6072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6900 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1624635492
transform -1 0 7912 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1624635492
transform -1 0 8096 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1624635492
transform -1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1624635492
transform -1 0 8464 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1624635492
transform -1 0 8648 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1624635492
transform -1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1624635492
transform 1 0 9936 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1624635492
transform -1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 9292 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1
timestamp 1624635492
transform -1 0 9936 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1
timestamp 1624635492
transform 1 0 9476 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1624635492
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 13248 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1624635492
transform -1 0 11776 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1624635492
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1624635492
transform -1 0 14260 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 16100 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1624635492
transform -1 0 15916 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1624635492
transform -1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 14904 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_149
timestamp 1624635492
transform 1 0 14812 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1624635492
transform 1 0 16928 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18860 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1624635492
transform -1 0 17940 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_183
timestamp 1624635492
transform 1 0 17940 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1624635492
transform -1 0 20608 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1624635492
transform -1 0 19504 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 19780 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 19136 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_193
timestamp 1624635492
transform 1 0 18860 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1624635492
transform 1 0 20608 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 21620 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3312 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1624635492
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4140 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1624635492
transform 1 0 3312 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1624635492
transform 1 0 4968 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7636 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1624635492
transform -1 0 7452 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1624635492
transform -1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1624635492
transform 1 0 10304 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9108 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1
timestamp 1624635492
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1624635492
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1624635492
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1624635492
transform 1 0 13340 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1624635492
transform 1 0 14168 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A0
timestamp 1624635492
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1624635492
transform 1 0 14996 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1624635492
transform -1 0 16652 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1624635492
transform -1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1624635492
transform -1 0 17204 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1624635492
transform -1 0 18860 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1624635492
transform -1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A1
timestamp 1624635492
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1624635492
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1624635492
transform -1 0 19596 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624635492
transform -1 0 19228 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1624635492
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1624635492
transform 1 0 20424 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1624635492
transform -1 0 21620 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 1656 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 1656 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1624635492
transform 1 0 4692 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1624635492
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1624635492
transform 1 0 3128 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 7084 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_48
timestamp 1624635492
transform 1 0 5520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 8188 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7084 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 8188 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A1
timestamp 1624635492
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 12420 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1624635492
transform 1 0 12420 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1624635492
transform 1 0 13432 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1624635492
transform -1 0 16008 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1624635492
transform -1 0 17020 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 17940 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17112 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_173
timestamp 1624635492
transform 1 0 17020 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1624635492
transform -1 0 20516 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_199
timestamp 1624635492
transform 1 0 19412 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_201
timestamp 1624635492
transform 1 0 19596 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1624635492
transform 1 0 20516 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 21620 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_220
timestamp 1624635492
transform 1 0 21344 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2944 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1624635492
transform 1 0 2116 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1624635492
transform 1 0 1748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1624635492
transform 1 0 4692 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 4600 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_38
timestamp 1624635492
transform 1 0 4600 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1624635492
transform -1 0 6348 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1624635492
transform -1 0 8924 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7268 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8924 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1624635492
transform 1 0 9752 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11592 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 12512 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 15364 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 12972 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_128
timestamp 1624635492
transform 1 0 12880 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 15364 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1624635492
transform -1 0 17756 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1624635492
transform 1 0 17756 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1624635492
transform -1 0 19412 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1624635492
transform -1 0 20516 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A1
timestamp 1624635492
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_199
timestamp 1624635492
transform 1 0 19412 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1624635492
transform 1 0 20516 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1624635492
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1624635492
transform 1 0 2300 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1624635492
transform -1 0 2300 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1624635492
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1624635492
transform 1 0 3496 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1624635492
transform 1 0 3128 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1624635492
transform -1 0 5888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 5888 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1624635492
transform 1 0 7912 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1624635492
transform 1 0 8740 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1624635492
transform -1 0 10764 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1624635492
transform -1 0 11592 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11776 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11960 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1624635492
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1624635492
transform 1 0 13248 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 14628 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 17112 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 15640 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 15180 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1624635492
transform -1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1624635492
transform -1 0 17940 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A1
timestamp 1624635492
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_183
timestamp 1624635492
transform 1 0 17940 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 19596 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1624635492
transform 1 0 18676 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A0
timestamp 1624635492
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1624635492
transform 1 0 18584 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1624635492
transform -1 0 21620 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 21252 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1624635492
transform 1 0 2392 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1624635492
transform 1 0 2300 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1624635492
transform 1 0 1564 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1624635492
transform -1 0 2300 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 1564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1624635492
transform -1 0 3404 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1624635492
transform 1 0 3220 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1624635492
transform -1 0 4784 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4416 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 6256 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_47
timestamp 1624635492
transform 1 0 5428 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1624635492
transform 1 0 5520 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1624635492
transform 1 0 6256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 6716 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1624635492
transform -1 0 7544 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8556 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7544 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 8556 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 6900 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 10580 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 9108 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1624635492
transform -1 0 11408 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1624635492
transform -1 0 11408 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_86
timestamp 1624635492
transform 1 0 9016 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1624635492
transform 1 0 8924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 13892 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 13156 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1624635492
transform -1 0 12420 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1624635492
transform -1 0 11592 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1624635492
transform 1 0 14444 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1624635492
transform 1 0 13524 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1624635492
transform 1 0 14352 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1624635492
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_144
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1624635492
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16468 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1624635492
transform 1 0 16100 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_155
timestamp 1624635492
transform 1 0 15364 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_176
timestamp 1624635492
transform 1 0 17296 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1624635492
transform 1 0 17756 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1624635492
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 17848 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1624635492
transform -1 0 19044 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 18860 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform 1 0 19044 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 19596 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 19504 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1624635492
transform -1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1624635492
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1624635492
transform 1 0 19044 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1624635492
transform 1 0 20516 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1624635492
transform -1 0 21620 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1624635492
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 21252 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 2300 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1624635492
transform -1 0 2300 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1624635492
transform -1 0 4692 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1624635492
transform 1 0 4692 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_29
timestamp 1624635492
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1624635492
transform 1 0 5520 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1624635492
transform 1 0 7820 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1624635492
transform -1 0 9936 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9936 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_92
timestamp 1624635492
transform 1 0 9568 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 13616 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1624635492
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1624635492
transform 1 0 14076 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 13892 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 14076 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 16008 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1624635492
transform -1 0 16008 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_150
timestamp 1624635492
transform 1 0 14904 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1624635492
transform -1 0 18584 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20516 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1624635492
transform -1 0 20240 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1624635492
transform -1 0 19412 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20792 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1624635492
transform -1 0 21620 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1624635492
transform -1 0 21252 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_214
timestamp 1624635492
transform 1 0 20792 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 3220 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1624635492
transform 1 0 3220 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1624635492
transform 1 0 4692 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6624 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1624635492
transform -1 0 6624 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1624635492
transform -1 0 5796 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1624635492
transform 1 0 8096 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1624635492
transform 1 0 10580 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1624635492
transform -1 0 10580 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 9568 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1624635492
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 13248 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1624635492
transform -1 0 14168 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1624635492
transform -1 0 15180 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_132
timestamp 1624635492
transform 1 0 13248 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_142
timestamp 1624635492
transform 1 0 14168 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 16008 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1624635492
transform 1 0 15180 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1624635492
transform -1 0 19044 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 17572 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 17756 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_178
timestamp 1624635492
transform 1 0 17480 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_183
timestamp 1624635492
transform 1 0 17940 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1624635492
transform 1 0 19044 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1624635492
transform 1 0 19596 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1624635492
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1624635492
transform -1 0 21068 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1624635492
transform -1 0 21620 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 21252 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 20792 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1624635492
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1624635492
transform 1 0 2944 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform -1 0 2944 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1624635492
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1624635492
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1624635492
transform 1 0 3588 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1624635492
transform 1 0 4416 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_26
timestamp 1624635492
transform 1 0 3496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1624635492
transform 1 0 5244 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 7912 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1624635492
transform 1 0 5520 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1624635492
transform 1 0 8740 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1624635492
transform -1 0 8740 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1624635492
transform -1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1624635492
transform -1 0 13340 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1624635492
transform -1 0 13616 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 15180 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_136
timestamp 1624635492
transform 1 0 13616 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1624635492
transform -1 0 16836 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1624635492
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1624635492
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_153
timestamp 1624635492
transform 1 0 15180 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_156
timestamp 1624635492
transform 1 0 15456 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_161
timestamp 1624635492
transform 1 0 15916 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 16928 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1624635492
transform 1 0 18400 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1624635492
transform -1 0 20056 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1624635492
transform -1 0 20516 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 20240 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1624635492
transform -1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1624635492
transform -1 0 20792 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1624635492
transform -1 0 21620 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1624635492
transform 1 0 2760 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1624635492
transform -1 0 2668 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1624635492
transform 1 0 1748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_17
timestamp 1624635492
transform 1 0 2668 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1624635492
transform 1 0 3956 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1624635492
transform -1 0 5244 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 4416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 6992 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_47
timestamp 1624635492
transform 1 0 5428 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1624635492
transform 1 0 8188 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11776 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9108 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1624635492
transform -1 0 12604 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12788 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14720 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1624635492
transform 1 0 16192 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1624635492
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17480 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 17020 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_175
timestamp 1624635492
transform 1 0 17204 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20240 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624635492
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 19136 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_201 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 19596 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_208
timestamp 1624635492
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output143
timestamp 1624635492
transform 1 0 21252 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output154
timestamp 1624635492
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 20884 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_212
timestamp 1624635492
transform 1 0 20608 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output135
timestamp 1624635492
transform -1 0 2116 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output134
timestamp 1624635492
transform -1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output123
timestamp 1624635492
transform -1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1624635492
transform -1 0 2024 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2668 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1624635492
transform -1 0 3772 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2392 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1624635492
transform 1 0 2116 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2024 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 4416 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1624635492
transform -1 0 4416 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_26
timestamp 1624635492
transform 1 0 3496 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1624635492
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 5888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 5336 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1624635492
transform 1 0 5888 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_56
timestamp 1624635492
transform 1 0 6256 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6716 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9476 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 8188 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 7728 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_71
timestamp 1624635492
transform 1 0 7636 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1624635492
transform 1 0 9292 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1624635492
transform -1 0 10212 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_102
timestamp 1624635492
transform 1 0 10488 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1624635492
transform -1 0 10488 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 10580 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1624635492
transform -1 0 11592 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1624635492
transform 1 0 12052 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_130
timestamp 1624635492
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_134
timestamp 1624635492
transform 1 0 13432 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1624635492
transform 1 0 13432 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1624635492
transform 1 0 13156 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 14076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 14628 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1624635492
transform 1 0 14076 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15824 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1624635492
transform 1 0 14904 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1624635492
transform 1 0 15732 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1624635492
transform 1 0 15824 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_172
timestamp 1624635492
transform 1 0 16928 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_172
timestamp 1624635492
transform 1 0 16928 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_168
timestamp 1624635492
transform 1 0 16560 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 16928 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1624635492
transform -1 0 17848 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1624635492
transform -1 0 17848 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1624635492
transform 1 0 17848 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17848 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1624635492
transform 1 0 19320 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624635492
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 19228 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_207 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 20148 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_199
timestamp 1624635492
transform 1 0 19412 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_201 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 19596 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_213
timestamp 1624635492
transform 1 0 20700 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1624635492
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  Test_en_N_FTB01
timestamp 1624635492
transform -1 0 20608 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_217
timestamp 1624635492
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_217
timestamp 1624635492
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1624635492
transform -1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1624635492
transform -1 0 21068 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output156
timestamp 1624635492
transform 1 0 21252 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output155
timestamp 1624635492
transform 1 0 21252 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1624635492
transform 1 0 2116 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1624635492
transform 1 0 2392 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2668 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output136
timestamp 1624635492
transform -1 0 1748 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output137
timestamp 1624635492
transform -1 0 2116 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1624635492
transform -1 0 3128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 4968 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1624635492
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_24
timestamp 1624635492
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5520 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_42
timestamp 1624635492
transform 1 0 4968 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1624635492
transform -1 0 8096 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 8280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_78
timestamp 1624635492
transform 1 0 8280 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10212 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1624635492
transform -1 0 10212 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_86
timestamp 1624635492
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1624635492
transform -1 0 12512 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 12512 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 14996 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1624635492
transform -1 0 13524 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 15088 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_151
timestamp 1624635492
transform 1 0 14996 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1624635492
transform -1 0 16836 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1624635492
transform -1 0 18768 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1624635492
transform 1 0 16928 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1624635492
transform -1 0 19596 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_201
timestamp 1624635492
transform 1 0 19596 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1624635492
transform -1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output157
timestamp 1624635492
transform 1 0 21252 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1624635492
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_209
timestamp 1624635492
transform 1 0 20332 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1624635492
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1624635492
transform 1 0 2116 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1624635492
transform 1 0 2576 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output138
timestamp 1624635492
transform -1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output139
timestamp 1624635492
transform -1 0 2116 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A1
timestamp 1624635492
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A0
timestamp 1624635492
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1624635492
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1624635492
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_39
timestamp 1624635492
transform 1 0 4692 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1624635492
transform 1 0 5428 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 6716 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 6440 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A1
timestamp 1624635492
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_45
timestamp 1624635492
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7544 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 10580 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1624635492
transform 1 0 10580 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1624635492
transform -1 0 13340 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1624635492
transform 1 0 11408 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_123
timestamp 1624635492
transform 1 0 12420 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 15824 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 13340 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_136
timestamp 1624635492
transform 1 0 13616 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_142
timestamp 1624635492
transform 1 0 14168 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 17572 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_22_160
timestamp 1624635492
transform 1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 17572 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1624635492
transform 1 0 19044 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1624635492
transform 1 0 19596 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624635492
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_198
timestamp 1624635492
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1624635492
transform -1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output158
timestamp 1624635492
transform 1 0 21252 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output159
timestamp 1624635492
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1624635492
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1624635492
transform 1 0 1748 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1624635492
transform 1 0 2024 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1624635492
transform 1 0 2300 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1624635492
transform 1 0 2668 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output140
timestamp 1624635492
transform -1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_16
timestamp 1624635492
transform 1 0 2576 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1624635492
transform 1 0 3496 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 4876 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1624635492
transform 1 0 4048 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A0
timestamp 1624635492
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_31
timestamp 1624635492
transform 1 0 3956 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 6716 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_58
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1624635492
transform 1 0 7268 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1624635492
transform -1 0 9476 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 8648 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A0
timestamp 1624635492
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_63
timestamp 1624635492
transform 1 0 6900 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_78
timestamp 1624635492
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9476 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1624635492
transform 1 0 10304 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11684 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1624635492
transform 1 0 11500 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1624635492
transform -1 0 13984 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1624635492
transform 1 0 14812 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1624635492
transform -1 0 16468 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_148
timestamp 1624635492
transform 1 0 14720 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 17480 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1624635492
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_167
timestamp 1624635492
transform 1 0 16468 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_172
timestamp 1624635492
transform 1 0 16928 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20240 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20516 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_194
timestamp 1624635492
transform 1 0 18952 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_202
timestamp 1624635492
transform 1 0 19688 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1624635492
transform -1 0 21068 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output160
timestamp 1624635492
transform 1 0 21252 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1624635492
transform -1 0 20792 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_211
timestamp 1624635492
transform 1 0 20516 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_217
timestamp 1624635492
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3772 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output141
timestamp 1624635492
transform -1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output142
timestamp 1624635492
transform -1 0 2116 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1624635492
transform -1 0 2300 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1624635492
transform 1 0 4416 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1624635492
transform 1 0 4140 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_35
timestamp 1624635492
transform 1 0 4324 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 6072 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1624635492
transform -1 0 6900 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1624635492
transform 1 0 7728 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1624635492
transform -1 0 7728 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 1624635492
transform 1 0 8004 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_83
timestamp 1624635492
transform 1 0 8740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1624635492
transform -1 0 11408 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1624635492
transform -1 0 13064 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 11868 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_112
timestamp 1624635492
transform 1 0 11408 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1624635492
transform 1 0 13892 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1624635492
transform -1 0 13892 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1624635492
transform 1 0 14168 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1624635492
transform -1 0 15364 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1624635492
transform -1 0 16192 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_164 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 16192 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1624635492
transform -1 0 18676 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_24_176
timestamp 1624635492
transform 1 0 17296 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1624635492
transform -1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1624635492
transform -1 0 20240 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1624635492
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1624635492
transform 1 0 19780 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1624635492
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_191
timestamp 1624635492
transform 1 0 18676 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_199
timestamp 1624635492
transform 1 0 19412 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1624635492
transform -1 0 21068 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1624635492
transform -1 0 20792 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output161
timestamp 1624635492
transform 1 0 21252 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1624635492
transform -1 0 21252 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1624635492
transform 1 0 2392 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1624635492
transform -1 0 2392 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1624635492
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1624635492
transform 1 0 3220 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1624635492
transform 1 0 3496 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1624635492
transform 1 0 3772 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1624635492
transform -1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_40
timestamp 1624635492
transform 1 0 4784 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1624635492
transform -1 0 6072 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1624635492
transform -1 0 7360 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A0
timestamp 1624635492
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A1
timestamp 1624635492
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_56
timestamp 1624635492
transform 1 0 6256 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_58
timestamp 1624635492
transform 1 0 6440 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1624635492
transform -1 0 8188 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1624635492
transform -1 0 9016 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 11132 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_25_86
timestamp 1624635492
transform 1 0 9016 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_92
timestamp 1624635492
transform 1 0 9568 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 11868 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_109
timestamp 1624635492
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1624635492
transform 1 0 11500 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1624635492
transform -1 0 14168 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1624635492
transform 1 0 14168 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1624635492
transform 1 0 16100 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1624635492
transform 1 0 15272 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 16560 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_151
timestamp 1624635492
transform 1 0 14996 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1624635492
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_168
timestamp 1624635492
transform 1 0 16560 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1624635492
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1624635492
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1624635492
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1624635492
transform 1 0 20240 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1624635492
transform -1 0 20884 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output144
timestamp 1624635492
transform 1 0 21252 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output162
timestamp 1624635492
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 3220 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform 1 0 2668 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1624635492
transform -1 0 2668 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output124
timestamp 1624635492
transform -1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output125
timestamp 1624635492
transform -1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1624635492
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1624635492
transform 1 0 3220 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1624635492
transform 1 0 3496 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4048 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1624635492
transform 1 0 4140 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1624635492
transform 1 0 3864 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 5520 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 6072 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1624635492
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1624635492
transform -1 0 5152 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_44
timestamp 1624635492
transform 1 0 5152 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_54
timestamp 1624635492
transform 1 0 6072 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 8740 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 8832 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1624635492
transform 1 0 7912 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_26_64
timestamp 1624635492
transform 1 0 6992 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_89
timestamp 1624635492
transform 1 0 9292 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_99
timestamp 1624635492
transform 1 0 10212 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1624635492
transform -1 0 11316 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1624635492
transform -1 0 10672 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10672 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 12420 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12328 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13156 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1624635492
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 11868 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_111
timestamp 1624635492
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_117
timestamp 1624635492
transform 1 0 11868 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 13892 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14352 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1624635492
transform 1 0 13156 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A1
timestamp 1624635492
transform -1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_142
timestamp 1624635492
transform 1 0 14168 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 17480 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 15364 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_26_160
timestamp 1624635492
transform 1 0 15824 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1624635492
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1624635492
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1624635492
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1624635492
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_196
timestamp 1624635492
transform 1 0 19136 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_190
timestamp 1624635492
transform 1 0 18584 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_204
timestamp 1624635492
transform 1 0 19872 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_201
timestamp 1624635492
transform 1 0 19596 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_198
timestamp 1624635492
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1624635492
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1624635492
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20240 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_207
timestamp 1624635492
transform 1 0 20148 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_208
timestamp 1624635492
transform 1 0 20240 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1624635492
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_210
timestamp 1624635492
transform 1 0 20424 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1624635492
transform 1 0 20332 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  prog_clk_3_S_FTB01
timestamp 1624635492
transform 1 0 20516 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1624635492
transform -1 0 20792 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1624635492
transform -1 0 21252 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_S_FTB01_A
timestamp 1624635492
transform -1 0 21252 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1624635492
transform -1 0 21068 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1624635492
transform -1 0 21068 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output146
timestamp 1624635492
transform 1 0 21252 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output145
timestamp 1624635492
transform 1 0 21252 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2944 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1624635492
transform 1 0 2116 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624635492
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output126
timestamp 1624635492
transform -1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output127
timestamp 1624635492
transform -1 0 2116 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1624635492
transform 1 0 4876 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1624635492
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1624635492
transform 1 0 3864 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1624635492
transform -1 0 6900 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A0
timestamp 1624635492
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_50
timestamp 1624635492
transform 1 0 5704 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1624635492
transform 1 0 7820 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1624635492
transform 1 0 6992 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_63
timestamp 1624635492
transform 1 0 6900 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9936 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1624635492
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A1
timestamp 1624635492
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1624635492
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 9752 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_89
timestamp 1624635492
transform 1 0 9292 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1624635492
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1624635492
transform 1 0 10764 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1624635492
transform -1 0 12420 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_125
timestamp 1624635492
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1624635492
transform -1 0 13616 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 13892 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15180 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1624635492
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_139
timestamp 1624635492
transform 1 0 13892 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16008 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1624635492
transform 1 0 16008 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_171
timestamp 1624635492
transform 1 0 16836 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_183
timestamp 1624635492
transform 1 0 17940 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1624635492
transform -1 0 20424 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  clk_2_S_FTB01
timestamp 1624635492
transform 1 0 19872 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1624635492
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_E_FTB01_A
timestamp 1624635492
transform 1 0 19688 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1624635492
transform 1 0 19320 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_195
timestamp 1624635492
transform 1 0 19044 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1624635492
transform 1 0 19596 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1624635492
transform -1 0 20700 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 21252 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624635492
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output147
timestamp 1624635492
transform 1 0 21252 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1624635492
transform 1 0 2116 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1624635492
transform 1 0 2392 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2668 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624635492
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output128
timestamp 1624635492
transform -1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output129
timestamp 1624635492
transform -1 0 2116 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1624635492
transform -1 0 3128 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1624635492
transform 1 0 3956 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1624635492
transform 1 0 3128 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_29_40
timestamp 1624635492
transform 1 0 4784 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1624635492
transform 1 0 6440 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1624635492
transform -1 0 6348 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1624635492
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 5520 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1624635492
transform -1 0 9108 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1624635492
transform -1 0 8280 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_67
timestamp 1624635492
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 9476 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_87
timestamp 1624635492
transform 1 0 9108 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1624635492
transform 1 0 10948 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11684 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1624635492
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_110
timestamp 1624635492
transform 1 0 11224 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1624635492
transform -1 0 14720 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_131
timestamp 1624635492
transform 1 0 13156 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_143
timestamp 1624635492
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1624635492
transform -1 0 16652 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 16100 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_148
timestamp 1624635492
transform 1 0 14720 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_163
timestamp 1624635492
transform 1 0 16100 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1624635492
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1624635492
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1624635492
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_184
timestamp 1624635492
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_190
timestamp 1624635492
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1624635492
transform -1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1624635492
transform -1 0 19136 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_199
timestamp 1624635492
transform 1 0 19412 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_196
timestamp 1624635492
transform 1 0 19136 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1624635492
transform -1 0 19412 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1624635492
transform -1 0 19688 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1624635492
transform -1 0 19964 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_205
timestamp 1624635492
transform 1 0 19964 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_N_FTB01
timestamp 1624635492
transform -1 0 20332 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  clk_3_S_FTB01
timestamp 1624635492
transform 1 0 20608 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_E_FTB01
timestamp 1624635492
transform -1 0 20608 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624635492
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output148
timestamp 1624635492
transform 1 0 21252 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output149
timestamp 1624635492
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1624635492
transform 1 0 1748 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1624635492
transform 1 0 2024 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1624635492
transform 1 0 2300 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624635492
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output130
timestamp 1624635492
transform -1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1624635492
transform -1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1624635492
transform -1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1624635492
transform -1 0 3128 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4416 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1624635492
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1624635492
transform -1 0 3312 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1624635492
transform -1 0 3496 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1624635492
transform -1 0 3680 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1624635492
transform 1 0 3864 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1624635492
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1624635492
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_28
timestamp 1624635492
transform 1 0 3680 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1624635492
transform 1 0 6808 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 6808 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_45
timestamp 1624635492
transform 1 0 5244 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1624635492
transform -1 0 8096 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1624635492
transform 1 0 8096 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1624635492
transform -1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 10580 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1624635492
transform -1 0 10580 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1624635492
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1624635492
transform 1 0 8924 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_87
timestamp 1624635492
transform 1 0 9108 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_93
timestamp 1624635492
transform 1 0 9660 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1624635492
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1624635492
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_119
timestamp 1624635492
transform 1 0 12052 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_124
timestamp 1624635492
transform 1 0 12512 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1624635492
transform 1 0 14352 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1624635492
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1624635492
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_127
timestamp 1624635492
transform 1 0 12788 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_130
timestamp 1624635492
transform 1 0 13064 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_142
timestamp 1624635492
transform 1 0 14168 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1624635492
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_149
timestamp 1624635492
transform 1 0 14812 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_161
timestamp 1624635492
transform 1 0 15916 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1624635492
transform -1 0 18308 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1624635492
transform -1 0 18032 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1624635492
transform 1 0 17020 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1624635492
transform 1 0 17388 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1624635492
transform 1 0 17664 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_175
timestamp 1624635492
transform 1 0 17204 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_179
timestamp 1624635492
transform 1 0 17572 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_184
timestamp 1624635492
transform 1 0 18032 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_187
timestamp 1624635492
transform 1 0 18308 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_190
timestamp 1624635492
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1624635492
transform -1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  clk_3_W_FTB01
timestamp 1624635492
transform -1 0 18952 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input103
timestamp 1624635492
transform -1 0 19228 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input102
timestamp 1624635492
transform -1 0 19504 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_201
timestamp 1624635492
transform 1 0 19596 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1624635492
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_E_FTB01
timestamp 1624635492
transform 1 0 19688 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_E_FTB01
timestamp 1624635492
transform -1 0 20240 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_N_FTB01
timestamp 1624635492
transform 1 0 20240 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624635492
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output150
timestamp 1624635492
transform 1 0 21252 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output213
timestamp 1624635492
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output220
timestamp 1624635492
transform 1 0 20516 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1624635492
transform 1 0 1748 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624635492
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input116
timestamp 1624635492
transform 1 0 2024 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input117
timestamp 1624635492
transform 1 0 2300 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input120
timestamp 1624635492
transform 1 0 2852 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output131
timestamp 1624635492
transform -1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output218
timestamp 1624635492
transform -1 0 2852 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5612 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 4048 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1624635492
transform -1 0 3772 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1624635492
transform -1 0 3312 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1624635492
transform -1 0 3496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_26
timestamp 1624635492
transform 1 0 3496 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1624635492
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 1624635492
transform 1 0 5888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1624635492
transform -1 0 5796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1624635492
transform -1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1624635492
transform -1 0 6624 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1624635492
transform -1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1624635492
transform -1 0 6992 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_51
timestamp 1624635492
transform 1 0 5796 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8464 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8464 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1624635492
transform -1 0 9936 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 9568 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1624635492
transform 1 0 10396 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 10212 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_92
timestamp 1624635492
transform 1 0 9568 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_99
timestamp 1624635492
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1624635492
transform 1 0 12512 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1624635492
transform -1 0 12512 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11500 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1624635492
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1624635492
transform 1 0 11500 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1624635492
transform -1 0 13064 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1624635492
transform -1 0 13340 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1624635492
transform -1 0 13616 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1624635492
transform -1 0 13892 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1624635492
transform -1 0 14628 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1624635492
transform -1 0 14076 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1624635492
transform -1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_141
timestamp 1624635492
transform 1 0 14076 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1624635492
transform -1 0 15088 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1624635492
transform -1 0 15364 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1624635492
transform -1 0 15824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  prog_clk_1_W_FTB01
timestamp 1624635492
transform -1 0 16192 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1624635492
transform -1 0 14812 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1624635492
transform -1 0 15548 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1624635492
transform -1 0 16376 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_160
timestamp 1624635492
transform 1 0 15824 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_166
timestamp 1624635492
transform 1 0 16376 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_170
timestamp 1624635492
transform 1 0 16744 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1624635492
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1624635492
transform -1 0 16744 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_174
timestamp 1624635492
transform 1 0 17112 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1624635492
transform -1 0 17112 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1624635492
transform -1 0 17480 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_178
timestamp 1624635492
transform 1 0 17480 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1624635492
transform -1 0 17848 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1624635492
transform -1 0 18308 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1624635492
transform -1 0 18124 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  prog_clk_3_W_FTB01
timestamp 1624635492
transform -1 0 18676 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  clk_1_W_FTB01
timestamp 1624635492
transform -1 0 18952 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  prog_clk_0_FTB00
timestamp 1624635492
transform 1 0 18952 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_E_FTB01
timestamp 1624635492
transform 1 0 21344 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01
timestamp 1624635492
transform 1 0 20792 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624635492
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624635492
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 1624635492
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input114
timestamp 1624635492
transform 1 0 2392 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input115
timestamp 1624635492
transform 1 0 2668 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1624635492
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output132
timestamp 1624635492
transform -1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output222
timestamp 1624635492
transform -1 0 2116 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 5428 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1624635492
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 1624635492
transform 1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input119
timestamp 1624635492
transform 1 0 3220 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1624635492
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1624635492
transform -1 0 5704 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 5796 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_32_50
timestamp 1624635492
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1624635492
transform 1 0 7636 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1624635492
transform -1 0 8740 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1624635492
transform 1 0 7268 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1624635492
transform -1 0 8924 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1624635492
transform 1 0 8924 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1624635492
transform -1 0 9292 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1624635492
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_91
timestamp 1624635492
transform 1 0 9476 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1624635492
transform -1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1624635492
transform -1 0 9936 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_96
timestamp 1624635492
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1624635492
transform -1 0 10304 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1624635492
transform -1 0 10580 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 1624635492
transform -1 0 10856 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1624635492
transform -1 0 11684 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12420 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1624635492
transform -1 0 11040 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1624635492
transform -1 0 11224 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1624635492
transform -1 0 11408 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1624635492
transform -1 0 11868 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_117
timestamp 1624635492
transform 1 0 11868 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1624635492
transform 1 0 12420 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1624635492
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output202
timestamp 1624635492
transform -1 0 14720 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_135
timestamp 1624635492
transform 1 0 13524 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_148
timestamp 1624635492
transform 1 0 14720 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_160
timestamp 1624635492
transform 1 0 15824 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input92
timestamp 1624635492
transform 1 0 18124 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 1624635492
transform 1 0 17848 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input104
timestamp 1624635492
transform 1 0 17572 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output215
timestamp 1624635492
transform 1 0 17296 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output216
timestamp 1624635492
transform 1 0 17020 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_W_FTB01_A
timestamp 1624635492
transform 1 0 16836 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_N_FTB01_A
timestamp 1624635492
transform -1 0 16836 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_168
timestamp 1624635492
transform 1 0 16560 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_E_FTB01
timestamp 1624635492
transform -1 0 19504 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  clk_2_W_FTB01
timestamp 1624635492
transform -1 0 18676 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1624635492
transform -1 0 19228 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1624635492
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output210
timestamp 1624635492
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output219
timestamp 1624635492
transform 1 0 19596 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1624635492
transform -1 0 21252 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624635492
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output151
timestamp 1624635492
transform 1 0 21252 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output209
timestamp 1624635492
transform 1 0 20332 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624635492
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output133
timestamp 1624635492
transform -1 0 1748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output204
timestamp 1624635492
transform -1 0 2116 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output208
timestamp 1624635492
transform -1 0 2484 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output212
timestamp 1624635492
transform -1 0 2852 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output214
timestamp 1624635492
transform -1 0 3220 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1624635492
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1624635492
transform 1 0 3220 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1624635492
transform 1 0 3864 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1624635492
transform 1 0 4232 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1624635492
transform 1 0 4784 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1624635492
transform -1 0 3772 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1624635492
transform -1 0 4784 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1624635492
transform -1 0 7360 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1624635492
transform 1 0 6440 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1624635492
transform -1 0 5520 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1624635492
transform -1 0 5888 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1624635492
transform 1 0 6072 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1624635492
transform -1 0 6072 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1624635492
transform -1 0 7728 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1624635492
transform -1 0 8188 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1624635492
transform -1 0 8556 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1624635492
transform -1 0 8924 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_72
timestamp 1624635492
transform 1 0 7728 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1624635492
transform 1 0 9108 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input77
timestamp 1624635492
transform -1 0 10764 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1624635492
transform -1 0 9752 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1624635492
transform -1 0 10120 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1624635492
transform -1 0 10488 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1624635492
transform -1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1624635492
transform -1 0 9384 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1624635492
transform 1 0 11776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output183
timestamp 1624635492
transform -1 0 11224 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output194
timestamp 1624635492
transform -1 0 11592 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output195
timestamp 1624635492
transform -1 0 12236 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output196
timestamp 1624635492
transform -1 0 12604 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output197
timestamp 1624635492
transform -1 0 12972 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_105
timestamp 1624635492
transform 1 0 10764 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1624635492
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1624635492
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output198
timestamp 1624635492
transform -1 0 13340 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output199
timestamp 1624635492
transform -1 0 13708 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output200
timestamp 1624635492
transform -1 0 14076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output201
timestamp 1624635492
transform -1 0 14444 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output184
timestamp 1624635492
transform -1 0 15088 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output185
timestamp 1624635492
transform -1 0 15456 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output186
timestamp 1624635492
transform -1 0 15824 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output187
timestamp 1624635492
transform -1 0 16192 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output188
timestamp 1624635492
transform -1 0 16652 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_146
timestamp 1624635492
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_164
timestamp 1624635492
transform 1 0 16192 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1624635492
transform 1 0 17112 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1624635492
transform -1 0 18584 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output189
timestamp 1624635492
transform -1 0 17020 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output190
timestamp 1624635492
transform -1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output191
timestamp 1624635492
transform -1 0 17940 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output192
timestamp 1624635492
transform -1 0 18308 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1624635492
transform 1 0 17020 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_N_FTB01
timestamp 1624635492
transform -1 0 20148 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1624635492
transform 1 0 19780 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output121
timestamp 1624635492
transform -1 0 18952 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output193
timestamp 1624635492
transform -1 0 19320 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output205
timestamp 1624635492
transform 1 0 20148 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output206
timestamp 1624635492
transform 1 0 19412 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_198
timestamp 1624635492
transform 1 0 19320 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624635492
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output152
timestamp 1624635492
transform 1 0 21252 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output153
timestamp 1624635492
transform 1 0 20884 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output203
timestamp 1624635492
transform 1 0 20516 0 1 20128
box -38 -48 406 592
<< labels >>
rlabel metal2 s 18602 22200 18658 23000 6 Test_en_N_out
port 0 nsew signal tristate
rlabel metal2 s 21086 0 21142 800 6 Test_en_S_in
port 1 nsew signal input
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 2 nsew signal input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 3 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 4 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 bottom_left_grid_pin_45_
port 5 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 bottom_left_grid_pin_46_
port 6 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 bottom_left_grid_pin_47_
port 7 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 bottom_left_grid_pin_48_
port 8 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 bottom_left_grid_pin_49_
port 9 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 ccff_head
port 10 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 ccff_tail
port 11 nsew signal tristate
rlabel metal3 s 0 3544 800 3664 6 chanx_left_in[0]
port 12 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[10]
port 13 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 chanx_left_in[11]
port 14 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[12]
port 15 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[13]
port 16 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[14]
port 17 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 chanx_left_in[15]
port 18 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[16]
port 19 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[17]
port 20 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 chanx_left_in[18]
port 21 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[19]
port 22 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 chanx_left_in[1]
port 23 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[2]
port 24 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[3]
port 25 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[4]
port 26 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 chanx_left_in[5]
port 27 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 chanx_left_in[6]
port 28 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 chanx_left_in[7]
port 29 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[8]
port 30 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 chanx_left_in[9]
port 31 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 chanx_left_out[0]
port 32 nsew signal tristate
rlabel metal3 s 0 16192 800 16312 6 chanx_left_out[10]
port 33 nsew signal tristate
rlabel metal3 s 0 16736 800 16856 6 chanx_left_out[11]
port 34 nsew signal tristate
rlabel metal3 s 0 17144 800 17264 6 chanx_left_out[12]
port 35 nsew signal tristate
rlabel metal3 s 0 17552 800 17672 6 chanx_left_out[13]
port 36 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[14]
port 37 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[15]
port 38 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[16]
port 39 nsew signal tristate
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[17]
port 40 nsew signal tristate
rlabel metal3 s 0 19592 800 19712 6 chanx_left_out[18]
port 41 nsew signal tristate
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[19]
port 42 nsew signal tristate
rlabel metal3 s 0 12384 800 12504 6 chanx_left_out[1]
port 43 nsew signal tristate
rlabel metal3 s 0 12792 800 12912 6 chanx_left_out[2]
port 44 nsew signal tristate
rlabel metal3 s 0 13336 800 13456 6 chanx_left_out[3]
port 45 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[4]
port 46 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[5]
port 47 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[6]
port 48 nsew signal tristate
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[7]
port 49 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 chanx_left_out[8]
port 50 nsew signal tristate
rlabel metal3 s 0 15784 800 15904 6 chanx_left_out[9]
port 51 nsew signal tristate
rlabel metal3 s 22200 3544 23000 3664 6 chanx_right_in[0]
port 52 nsew signal input
rlabel metal3 s 22200 7760 23000 7880 6 chanx_right_in[10]
port 53 nsew signal input
rlabel metal3 s 22200 8168 23000 8288 6 chanx_right_in[11]
port 54 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[12]
port 55 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[13]
port 56 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[14]
port 57 nsew signal input
rlabel metal3 s 22200 9800 23000 9920 6 chanx_right_in[15]
port 58 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[16]
port 59 nsew signal input
rlabel metal3 s 22200 10752 23000 10872 6 chanx_right_in[17]
port 60 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[18]
port 61 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[19]
port 62 nsew signal input
rlabel metal3 s 22200 3952 23000 4072 6 chanx_right_in[1]
port 63 nsew signal input
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[2]
port 64 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[3]
port 65 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[4]
port 66 nsew signal input
rlabel metal3 s 22200 5584 23000 5704 6 chanx_right_in[5]
port 67 nsew signal input
rlabel metal3 s 22200 5992 23000 6112 6 chanx_right_in[6]
port 68 nsew signal input
rlabel metal3 s 22200 6400 23000 6520 6 chanx_right_in[7]
port 69 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[8]
port 70 nsew signal input
rlabel metal3 s 22200 7352 23000 7472 6 chanx_right_in[9]
port 71 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_out[0]
port 72 nsew signal tristate
rlabel metal3 s 22200 16192 23000 16312 6 chanx_right_out[10]
port 73 nsew signal tristate
rlabel metal3 s 22200 16736 23000 16856 6 chanx_right_out[11]
port 74 nsew signal tristate
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[12]
port 75 nsew signal tristate
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[13]
port 76 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[14]
port 77 nsew signal tristate
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[15]
port 78 nsew signal tristate
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[16]
port 79 nsew signal tristate
rlabel metal3 s 22200 19184 23000 19304 6 chanx_right_out[17]
port 80 nsew signal tristate
rlabel metal3 s 22200 19592 23000 19712 6 chanx_right_out[18]
port 81 nsew signal tristate
rlabel metal3 s 22200 20136 23000 20256 6 chanx_right_out[19]
port 82 nsew signal tristate
rlabel metal3 s 22200 12384 23000 12504 6 chanx_right_out[1]
port 83 nsew signal tristate
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_out[2]
port 84 nsew signal tristate
rlabel metal3 s 22200 13336 23000 13456 6 chanx_right_out[3]
port 85 nsew signal tristate
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[4]
port 86 nsew signal tristate
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[5]
port 87 nsew signal tristate
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[6]
port 88 nsew signal tristate
rlabel metal3 s 22200 14968 23000 15088 6 chanx_right_out[7]
port 89 nsew signal tristate
rlabel metal3 s 22200 15376 23000 15496 6 chanx_right_out[8]
port 90 nsew signal tristate
rlabel metal3 s 22200 15784 23000 15904 6 chanx_right_out[9]
port 91 nsew signal tristate
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_in[0]
port 92 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 chany_bottom_in[10]
port 93 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[11]
port 94 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[12]
port 95 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[13]
port 96 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 chany_bottom_in[14]
port 97 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 chany_bottom_in[15]
port 98 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[16]
port 99 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[17]
port 100 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[18]
port 101 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 chany_bottom_in[19]
port 102 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_in[1]
port 103 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_in[2]
port 104 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_in[3]
port 105 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_in[4]
port 106 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[5]
port 107 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_in[6]
port 108 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[7]
port 109 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[8]
port 110 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[9]
port 111 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_out[0]
port 112 nsew signal tristate
rlabel metal2 s 16854 0 16910 800 6 chany_bottom_out[10]
port 113 nsew signal tristate
rlabel metal2 s 17314 0 17370 800 6 chany_bottom_out[11]
port 114 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[12]
port 115 nsew signal tristate
rlabel metal2 s 18142 0 18198 800 6 chany_bottom_out[13]
port 116 nsew signal tristate
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[14]
port 117 nsew signal tristate
rlabel metal2 s 18970 0 19026 800 6 chany_bottom_out[15]
port 118 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 chany_bottom_out[16]
port 119 nsew signal tristate
rlabel metal2 s 19798 0 19854 800 6 chany_bottom_out[17]
port 120 nsew signal tristate
rlabel metal2 s 20258 0 20314 800 6 chany_bottom_out[18]
port 121 nsew signal tristate
rlabel metal2 s 20626 0 20682 800 6 chany_bottom_out[19]
port 122 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_out[1]
port 123 nsew signal tristate
rlabel metal2 s 13542 0 13598 800 6 chany_bottom_out[2]
port 124 nsew signal tristate
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_out[3]
port 125 nsew signal tristate
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_out[4]
port 126 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 chany_bottom_out[5]
port 127 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_out[6]
port 128 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_out[7]
port 129 nsew signal tristate
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_out[8]
port 130 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[9]
port 131 nsew signal tristate
rlabel metal2 s 3238 22200 3294 23000 6 chany_top_in[0]
port 132 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[10]
port 133 nsew signal input
rlabel metal2 s 7470 22200 7526 23000 6 chany_top_in[11]
port 134 nsew signal input
rlabel metal2 s 7838 22200 7894 23000 6 chany_top_in[12]
port 135 nsew signal input
rlabel metal2 s 8206 22200 8262 23000 6 chany_top_in[13]
port 136 nsew signal input
rlabel metal2 s 8574 22200 8630 23000 6 chany_top_in[14]
port 137 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[15]
port 138 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[16]
port 139 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[17]
port 140 nsew signal input
rlabel metal2 s 10138 22200 10194 23000 6 chany_top_in[18]
port 141 nsew signal input
rlabel metal2 s 10506 22200 10562 23000 6 chany_top_in[19]
port 142 nsew signal input
rlabel metal2 s 3606 22200 3662 23000 6 chany_top_in[1]
port 143 nsew signal input
rlabel metal2 s 3974 22200 4030 23000 6 chany_top_in[2]
port 144 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[3]
port 145 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[4]
port 146 nsew signal input
rlabel metal2 s 5170 22200 5226 23000 6 chany_top_in[5]
port 147 nsew signal input
rlabel metal2 s 5538 22200 5594 23000 6 chany_top_in[6]
port 148 nsew signal input
rlabel metal2 s 5906 22200 5962 23000 6 chany_top_in[7]
port 149 nsew signal input
rlabel metal2 s 6274 22200 6330 23000 6 chany_top_in[8]
port 150 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[9]
port 151 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_out[0]
port 152 nsew signal tristate
rlabel metal2 s 14738 22200 14794 23000 6 chany_top_out[10]
port 153 nsew signal tristate
rlabel metal2 s 15106 22200 15162 23000 6 chany_top_out[11]
port 154 nsew signal tristate
rlabel metal2 s 15474 22200 15530 23000 6 chany_top_out[12]
port 155 nsew signal tristate
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[13]
port 156 nsew signal tristate
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[14]
port 157 nsew signal tristate
rlabel metal2 s 16670 22200 16726 23000 6 chany_top_out[15]
port 158 nsew signal tristate
rlabel metal2 s 17038 22200 17094 23000 6 chany_top_out[16]
port 159 nsew signal tristate
rlabel metal2 s 17406 22200 17462 23000 6 chany_top_out[17]
port 160 nsew signal tristate
rlabel metal2 s 17774 22200 17830 23000 6 chany_top_out[18]
port 161 nsew signal tristate
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[19]
port 162 nsew signal tristate
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_out[1]
port 163 nsew signal tristate
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_out[2]
port 164 nsew signal tristate
rlabel metal2 s 12070 22200 12126 23000 6 chany_top_out[3]
port 165 nsew signal tristate
rlabel metal2 s 12438 22200 12494 23000 6 chany_top_out[4]
port 166 nsew signal tristate
rlabel metal2 s 12806 22200 12862 23000 6 chany_top_out[5]
port 167 nsew signal tristate
rlabel metal2 s 13174 22200 13230 23000 6 chany_top_out[6]
port 168 nsew signal tristate
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[7]
port 169 nsew signal tristate
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[8]
port 170 nsew signal tristate
rlabel metal2 s 14370 22200 14426 23000 6 chany_top_out[9]
port 171 nsew signal tristate
rlabel metal3 s 22200 20544 23000 20664 6 clk_1_E_out
port 172 nsew signal tristate
rlabel metal2 s 18970 22200 19026 23000 6 clk_1_N_in
port 173 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 clk_1_W_out
port 174 nsew signal tristate
rlabel metal3 s 22200 20952 23000 21072 6 clk_2_E_out
port 175 nsew signal tristate
rlabel metal2 s 19338 22200 19394 23000 6 clk_2_N_in
port 176 nsew signal input
rlabel metal2 s 21638 22200 21694 23000 6 clk_2_N_out
port 177 nsew signal tristate
rlabel metal2 s 21454 0 21510 800 6 clk_2_S_out
port 178 nsew signal tristate
rlabel metal3 s 0 20952 800 21072 6 clk_2_W_out
port 179 nsew signal tristate
rlabel metal3 s 22200 21360 23000 21480 6 clk_3_E_out
port 180 nsew signal tristate
rlabel metal2 s 19706 22200 19762 23000 6 clk_3_N_in
port 181 nsew signal input
rlabel metal2 s 22006 22200 22062 23000 6 clk_3_N_out
port 182 nsew signal tristate
rlabel metal2 s 21914 0 21970 800 6 clk_3_S_out
port 183 nsew signal tristate
rlabel metal3 s 0 21360 800 21480 6 clk_3_W_out
port 184 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 185 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 186 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 187 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 left_bottom_grid_pin_37_
port 188 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 left_bottom_grid_pin_38_
port 189 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 left_bottom_grid_pin_39_
port 190 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 left_bottom_grid_pin_40_
port 191 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 left_bottom_grid_pin_41_
port 192 nsew signal input
rlabel metal2 s 20074 22200 20130 23000 6 prog_clk_0_N_in
port 193 nsew signal input
rlabel metal3 s 22200 21768 23000 21888 6 prog_clk_1_E_out
port 194 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 prog_clk_1_N_in
port 195 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 prog_clk_1_W_out
port 196 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 prog_clk_2_E_out
port 197 nsew signal tristate
rlabel metal2 s 20902 22200 20958 23000 6 prog_clk_2_N_in
port 198 nsew signal input
rlabel metal2 s 22374 22200 22430 23000 6 prog_clk_2_N_out
port 199 nsew signal tristate
rlabel metal2 s 22282 0 22338 800 6 prog_clk_2_S_out
port 200 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 prog_clk_2_W_out
port 201 nsew signal tristate
rlabel metal3 s 22200 22584 23000 22704 6 prog_clk_3_E_out
port 202 nsew signal tristate
rlabel metal2 s 21270 22200 21326 23000 6 prog_clk_3_N_in
port 203 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 prog_clk_3_N_out
port 204 nsew signal tristate
rlabel metal2 s 22742 0 22798 800 6 prog_clk_3_S_out
port 205 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 prog_clk_3_W_out
port 206 nsew signal tristate
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 207 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 208 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 209 nsew signal input
rlabel metal3 s 22200 1368 23000 1488 6 right_bottom_grid_pin_37_
port 210 nsew signal input
rlabel metal3 s 22200 1776 23000 1896 6 right_bottom_grid_pin_38_
port 211 nsew signal input
rlabel metal3 s 22200 2184 23000 2304 6 right_bottom_grid_pin_39_
port 212 nsew signal input
rlabel metal3 s 22200 2592 23000 2712 6 right_bottom_grid_pin_40_
port 213 nsew signal input
rlabel metal3 s 22200 3000 23000 3120 6 right_bottom_grid_pin_41_
port 214 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 215 nsew signal input
rlabel metal2 s 570 22200 626 23000 6 top_left_grid_pin_43_
port 216 nsew signal input
rlabel metal2 s 938 22200 994 23000 6 top_left_grid_pin_44_
port 217 nsew signal input
rlabel metal2 s 1306 22200 1362 23000 6 top_left_grid_pin_45_
port 218 nsew signal input
rlabel metal2 s 1674 22200 1730 23000 6 top_left_grid_pin_46_
port 219 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_47_
port 220 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_48_
port 221 nsew signal input
rlabel metal2 s 2870 22200 2926 23000 6 top_left_grid_pin_49_
port 222 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 223 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 224 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 225 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 226 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 227 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
