* NGSPICE file created from tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_1 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_2 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

.subckt tile VGND VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_ bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ ccff_head_1 ccff_head_2 ccff_tail ccff_tail_0 chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23] chanx_left_in[24]
+ chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28] chanx_left_in[29]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23] chanx_left_out[24]
+ chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28] chanx_left_out[29]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in_0[0] chanx_right_in_0[10]
+ chanx_right_in_0[11] chanx_right_in_0[12] chanx_right_in_0[13] chanx_right_in_0[14]
+ chanx_right_in_0[15] chanx_right_in_0[16] chanx_right_in_0[17] chanx_right_in_0[18]
+ chanx_right_in_0[19] chanx_right_in_0[1] chanx_right_in_0[20] chanx_right_in_0[21]
+ chanx_right_in_0[22] chanx_right_in_0[23] chanx_right_in_0[24] chanx_right_in_0[25]
+ chanx_right_in_0[26] chanx_right_in_0[27] chanx_right_in_0[28] chanx_right_in_0[29]
+ chanx_right_in_0[2] chanx_right_in_0[3] chanx_right_in_0[4] chanx_right_in_0[5]
+ chanx_right_in_0[6] chanx_right_in_0[7] chanx_right_in_0[8] chanx_right_in_0[9]
+ chanx_right_out_0[0] chanx_right_out_0[10] chanx_right_out_0[11] chanx_right_out_0[12]
+ chanx_right_out_0[13] chanx_right_out_0[14] chanx_right_out_0[15] chanx_right_out_0[16]
+ chanx_right_out_0[17] chanx_right_out_0[18] chanx_right_out_0[19] chanx_right_out_0[1]
+ chanx_right_out_0[20] chanx_right_out_0[21] chanx_right_out_0[22] chanx_right_out_0[23]
+ chanx_right_out_0[24] chanx_right_out_0[25] chanx_right_out_0[26] chanx_right_out_0[27]
+ chanx_right_out_0[28] chanx_right_out_0[29] chanx_right_out_0[2] chanx_right_out_0[3]
+ chanx_right_out_0[4] chanx_right_out_0[5] chanx_right_out_0[6] chanx_right_out_0[7]
+ chanx_right_out_0[8] chanx_right_out_0[9] chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21] chany_bottom_in[22]
+ chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25] chany_bottom_in[26]
+ chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21] chany_bottom_out[22]
+ chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25] chany_bottom_out[26]
+ chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in_0[0] chany_top_in_0[10]
+ chany_top_in_0[11] chany_top_in_0[12] chany_top_in_0[13] chany_top_in_0[14] chany_top_in_0[15]
+ chany_top_in_0[16] chany_top_in_0[17] chany_top_in_0[18] chany_top_in_0[19] chany_top_in_0[1]
+ chany_top_in_0[20] chany_top_in_0[21] chany_top_in_0[22] chany_top_in_0[23] chany_top_in_0[24]
+ chany_top_in_0[25] chany_top_in_0[26] chany_top_in_0[27] chany_top_in_0[28] chany_top_in_0[29]
+ chany_top_in_0[2] chany_top_in_0[3] chany_top_in_0[4] chany_top_in_0[5] chany_top_in_0[6]
+ chany_top_in_0[7] chany_top_in_0[8] chany_top_in_0[9] chany_top_out_0[0] chany_top_out_0[10]
+ chany_top_out_0[11] chany_top_out_0[12] chany_top_out_0[13] chany_top_out_0[14]
+ chany_top_out_0[15] chany_top_out_0[16] chany_top_out_0[17] chany_top_out_0[18]
+ chany_top_out_0[19] chany_top_out_0[1] chany_top_out_0[20] chany_top_out_0[21] chany_top_out_0[22]
+ chany_top_out_0[23] chany_top_out_0[24] chany_top_out_0[25] chany_top_out_0[26]
+ chany_top_out_0[27] chany_top_out_0[28] chany_top_out_0[29] chany_top_out_0[2] chany_top_out_0[3]
+ chany_top_out_0[4] chany_top_out_0[5] chany_top_out_0[6] chany_top_out_0[7] chany_top_out_0[8]
+ chany_top_out_0[9] clk0 prog_clk prog_reset_bottom_in prog_reset_bottom_out prog_reset_left_in
+ prog_reset_right_out prog_reset_top_in prog_reset_top_out reset_bottom_in reset_bottom_out
+ reset_left_out reset_right_in reset_top_in reset_top_out right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ right_width_0_height_0_subtile_0__pin_O_10_
+ right_width_0_height_0_subtile_0__pin_O_11_ right_width_0_height_0_subtile_0__pin_O_12_
+ right_width_0_height_0_subtile_0__pin_O_13_ right_width_0_height_0_subtile_0__pin_O_14_
+ right_width_0_height_0_subtile_0__pin_O_15_ right_width_0_height_0_subtile_0__pin_O_8_
+ right_width_0_height_0_subtile_0__pin_O_9_ sc_in sc_out test_enable_bottom_in test_enable_bottom_out
+ test_enable_left_out test_enable_right_in test_enable_top_in test_enable_top_out
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
+ top_width_0_height_0_subtile_0__pin_O_0_ top_width_0_height_0_subtile_0__pin_O_1_
+ top_width_0_height_0_subtile_0__pin_O_2_ top_width_0_height_0_subtile_0__pin_O_3_
+ top_width_0_height_0_subtile_0__pin_O_4_ top_width_0_height_0_subtile_0__pin_O_5_
+ top_width_0_height_0_subtile_0__pin_O_6_ top_width_0_height_0_subtile_0__pin_O_7_
+ top_width_0_height_0_subtile_0__pin_cin_0_ top_width_0_height_0_subtile_0__pin_reg_in_0_
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_1__S sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_37.mux_l1_in_1_ net68 net38 sb_1__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_35_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_53_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_53_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input127_A reset_right_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_3_ net321 net116 cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_3__379 VGND VGND VPWR VPWR net379 sb_1__1_.mux_bottom_track_21.mux_l2_in_3__379/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_363_ net81 VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input92_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_294_ net11 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_10.mux_l4_in_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_right_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l2_in_0_ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_3_ sb_1__1_.mux_bottom_track_29.out net69 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_2_ net14 net35 cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_0_ net122 net108 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_4__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_41_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_37_prog_clk
+ sb_1__1_.mem_bottom_track_13.ccff_tail net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_3.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_2_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_346_ net92 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output296_A net296 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_277_ sb_1__1_.mux_left_track_1.out VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ net150 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_23_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_3__A0 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_0.mux_l2_in_3_ net409 net4 sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_64_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_28.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_20_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput253 net253 VGND VGND VPWR VPWR chany_top_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput242 net242 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
Xoutput220 net220 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
Xoutput231 net231 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xoutput264 net264 VGND VGND VPWR VPWR chany_top_out_0[27] sky130_fd_sc_hd__buf_12
Xoutput286 net286 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_15_
+ sky130_fd_sc_hd__buf_12
Xoutput275 net275 VGND VGND VPWR VPWR prog_reset_bottom_out sky130_fd_sc_hd__buf_12
Xoutput297 net297 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_4_ sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_10.mux_l3_in_1_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l1_in_1_ net65 net134 sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_input55_A chanx_right_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_3.mux_l1_in_1_ net48 net93 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in net138 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__351
+ VGND VGND VPWR VPWR net351 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__351/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_46_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l2_in_3__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_1__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__330
+ VGND VGND VPWR VPWR net330 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__330/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_2__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_329_ net107 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_39_prog_clk sb_1__1_.mem_bottom_track_5.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_3.mux_l4_in_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_14.mux_l3_in_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_10.mux_l2_in_2__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_8_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_21.mux_l2_in_2__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_7.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA__312__A net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_4__S sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_ net149 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_10.mux_l2_in_2_ net13 sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_right_track_10.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_3_ net326 sb_1__1_.mux_bottom_track_53.out cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_4__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_2__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_0.mux_l4_in_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input18_A chanx_left_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__341
+ VGND VGND VPWR VPWR net341 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__341/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_45_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_4__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_2__A0 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_3.mux_l3_in_1_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_6_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_1__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk sb_1__1_.mem_right_track_28.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_1_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_89_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_2.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_top_track_28.mux_l2_in_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput120 chany_top_in_0[7] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
Xinput142 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND VGND VPWR
+ VPWR net142 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput131 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND VGND VPWR
+ VPWR net131 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_3__A1 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_12_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_10.mux_l1_in_3_ net75 net136 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_2__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_4_ net94 net92 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l2_in_3__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l2_in_1__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_37.mux_l1_in_0_ net98 net110 sb_1__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_4__A0 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_0.mux_l3_in_1_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_top_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_22_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_22_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_2_ net85 sb_1__1_.mux_bottom_track_37.out cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_45_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_362_ sb_1__1_.mux_top_track_10.out VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_293_ sb_1__1_.mux_right_track_28.out VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input85_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_top_track_12.mux_l1_in_1__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l4_in_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_36_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_2_ net107 net76 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_1_ net4 cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__320__A net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.out sky130_fd_sc_hd__clkbuf_2
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_41_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_28.mux_l1_in_1_ net44 net61 sb_1__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_1.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net368 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_345_ sb_1__1_.mux_top_track_44.out VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_2
X_276_ sb_1__1_.mux_left_track_3.out VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_3__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_0.mux_l2_in_2_ net21 net24 sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_28.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput210 net210 VGND VGND VPWR VPWR chanx_right_out_0[5] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput243 net243 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
Xoutput221 net221 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
Xoutput232 net232 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
Xoutput265 net265 VGND VGND VPWR VPWR chany_top_out_0[28] sky130_fd_sc_hd__buf_12
Xoutput254 net254 VGND VGND VPWR VPWR chany_top_out_0[18] sky130_fd_sc_hd__buf_12
XFILLER_87_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput276 net276 VGND VGND VPWR VPWR prog_reset_right_out sky130_fd_sc_hd__buf_12
Xoutput298 net298 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_5_ sky130_fd_sc_hd__buf_12
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput287 net287 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_8_ sky130_fd_sc_hd__buf_12
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_10.mux_l3_in_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l1_in_0_ net117 net95 sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l3_in_1_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net347 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_13.mux_l1_in_2_ net41 net10 cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input48_A chanx_right_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.out sky130_fd_sc_hd__buf_4
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_3.mux_l1_in_0_ net122 net108 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_1__A0 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_328_ net106 VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_2
X_259_ sb_1__1_.mux_left_track_37.out VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_41_prog_clk sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_56_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__353
+ VGND VGND VPWR VPWR net353 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__353/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_53.mux_l1_in_2__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input102_A chany_top_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_0.mux_l1_in_3_ net64 net81 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_3__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_0__A0 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_right_track_10.mux_l2_in_1_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_65_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_2_ net86 cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_3__305 VGND VGND VPWR VPWR net305 cbx_1__1_.mux_top_ipin_3.mux_l2_in_3__305/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_80_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_47_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_2__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_2__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_3.mux_l3_in_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_34_prog_clk sb_1__1_.mem_right_track_20.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net361 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__mux2_2
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_89_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_2__A0 net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_20.mux_l1_in_1__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput110 chany_top_in_0[25] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput121 chany_top_in_0[8] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput143 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND VGND VPWR
+ VPWR net143 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput132 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND VGND VPWR
+ VPWR net132 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input30_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_0.mux_l2_in_2__A0 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_42_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_10.mux_l1_in_2_ net134 net132 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_3_ sb_1__1_.mux_bottom_track_29.out net69 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__318__A net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_1.mux_l2_in_3__387 VGND VGND VPWR VPWR net387 sb_1__1_.mux_left_track_1.mux_l2_in_3__387/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_0.mux_l3_in_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_top_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_1_ net65 cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_361_ sb_1__1_.mux_top_track_12.out VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_21.mux_l2_in_3_ net390 net300 sb_1__1_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_292_ net9 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input78_A chany_bottom_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_0__A0 sb_1__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk sb_1__1_.mem_left_track_11.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_37_prog_clk
+ sb_1__1_.mem_bottom_track_13.mem_out\[2\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_32_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_28.mux_l1_in_0_ net39 net141 sb_1__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_41_prog_clk net429 net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input132_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_344_ net90 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_1__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_275_ sb_1__1_.mux_left_track_5.out VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk
+ sb_1__1_.mem_bottom_track_45.mem_out\[1\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_45.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l2_in_3__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_0.mux_l2_in_1_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk sb_1__1_.mem_top_track_28.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_20_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__365
+ VGND VGND VPWR VPWR net365 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__365/LO
+ sky130_fd_sc_hd__conb_1
Xoutput200 net200 VGND VGND VPWR VPWR chanx_right_out_0[23] sky130_fd_sc_hd__buf_12
Xcby_1__1_.mux_right_ipin_3.mux_l1_in_2_ net106 net75 cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xoutput211 net211 VGND VGND VPWR VPWR chanx_right_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput233 net233 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
Xoutput244 net244 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
Xoutput222 net222 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
Xoutput277 net277 VGND VGND VPWR VPWR prog_reset_top_out sky130_fd_sc_hd__buf_12
Xoutput266 net266 VGND VGND VPWR VPWR chany_top_out_0[29] sky130_fd_sc_hd__buf_12
Xoutput255 net255 VGND VGND VPWR VPWR chany_top_out_0[19] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput299 net299 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_6_ sky130_fd_sc_hd__buf_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput288 net288 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_9_ sky130_fd_sc_hd__buf_12
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net138 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_top_track_28.mux_l2_in_3__414 VGND VGND VPWR VPWR net414 sb_1__1_.mux_top_track_28.mux_l2_in_3__414/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net304 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_4__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_2.mux_l2_in_3_ net401 net32 sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l3_in_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_13.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_327_ sb_1__1_.mux_bottom_track_21.out VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_0__A0 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_258_ net35 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_41_prog_clk sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_6_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_3__A0 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_21.mux_l4_in_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA__326__A net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_53.mux_l1_in_2__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_4.mux_l1_in_0__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_0.mux_l1_in_2_ net34 net51 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_3_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input60_A chanx_right_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_left_track_13.mux_l2_in_3__389 VGND VGND VPWR VPWR net389 sb_1__1_.mux_left_track_13.mux_l2_in_3__389/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_93_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_3__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_3__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_0__A1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l2_in_3__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.out sky130_fd_sc_hd__buf_4
Xsb_1__1_.mux_right_track_10.mux_l2_in_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_1_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_16_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l2_in_2__A0 net296 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_32_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_2__A0 net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_21.mux_l3_in_1_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_56_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_2.mux_l4_in_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_right_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_18_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_2__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput111 chany_top_in_0[26] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_4
Xinput100 chany_top_in_0[16] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
Xinput144 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND VGND VPWR
+ VPWR net144 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput122 chany_top_in_0[9] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_4
Xinput133 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND VGND VPWR
+ VPWR net133 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input23_A chanx_left_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_48_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_0.mux_l2_in_2__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_10.mux_l1_in_1_ net130 net118 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_2_ net107 net76 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_79_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net357 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_1__A0 sb_1__1_.mux_left_track_11.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__334__A sb_1__1_.mux_bottom_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_360_ net78 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_21.mux_l2_in_2_ net294 net85 sb_1__1_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_291_ net8 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_31_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_31_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_3_ net305 net56 cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_16_prog_clk sb_1__1_.mem_left_track_11.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_76_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk
+ sb_1__1_.mem_bottom_track_13.mem_out\[1\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_2.mux_l3_in_1_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_right_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_83_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__329__A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.out sky130_fd_sc_hd__buf_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_33_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_3__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input125_A prog_reset_top_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_343_ net89 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_2
X_274_ sb_1__1_.mux_left_track_7.out VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input90_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_12.mux_l2_in_3_ net411 net26 sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk
+ sb_1__1_.mem_bottom_track_45.mem_out\[0\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_45.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_0.mux_l2_in_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_20.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_3.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xoutput201 net201 VGND VGND VPWR VPWR chanx_right_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput212 net212 VGND VGND VPWR VPWR chanx_right_out_0[7] sky130_fd_sc_hd__buf_12
Xoutput223 net223 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
Xoutput234 net234 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
Xoutput256 net256 VGND VGND VPWR VPWR chany_top_out_0[1] sky130_fd_sc_hd__buf_12
Xoutput267 net267 VGND VGND VPWR VPWR chany_top_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput245 net245 VGND VGND VPWR VPWR chany_top_out_0[0] sky130_fd_sc_hd__buf_12
Xoutput289 net289 VGND VGND VPWR VPWR sc_out sky130_fd_sc_hd__buf_12
Xoutput278 net278 VGND VGND VPWR VPWR reset_bottom_out sky130_fd_sc_hd__buf_12
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_2.mux_l2_in_2_ net18 net91 sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_78_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net365 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_29_prog_clk sb_1__1_.mem_right_track_2.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_326_ net103 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
XANTENNA_output294_A net294 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_0__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_257_ net34 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_3.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_3__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_3.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA__342__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__373
+ VGND VGND VPWR VPWR net373 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__373/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_68_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_0.mux_l1_in_1_ net53 net145 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA__252__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input53_A chanx_right_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_61_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_3__420 VGND VGND VPWR VPWR net420 cbx_1__1_.mux_top_ipin_0.mux_l2_in_3__420/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_91_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_309_ net115 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l2_in_2__A0 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_0__S sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_80_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_2.mux_l1_in_3_ net92 net78 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l1_in_1__A0 sb_1__1_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_12.mux_l4_in_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_3_ net310 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_56_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_left_track_1.mux_l2_in_2__A1 net293 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_2__A1 net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_3__381 VGND VGND VPWR VPWR net381 sb_1__1_.mux_bottom_track_3.mux_l2_in_3__381/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_left_track_21.mux_l3_in_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_53.mux_l2_in_1__396 VGND VGND VPWR VPWR net396 sb_1__1_.mux_left_track_53.mux_l2_in_1__396/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__1_.mux_top_ipin_3.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_3_ net380 net14 sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_0__A0 net141 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xinput101 chany_top_in_0[17] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput145 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND VGND VPWR
+ VPWR net145 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput112 chany_top_in_0[27] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
Xinput134 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND VGND VPWR
+ VPWR net134 sky130_fd_sc_hd__clkbuf_2
Xinput123 prog_reset_bottom_in VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input16_A chanx_left_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net343 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__mux2_4
XFILLER_8_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_10.mux_l1_in_0_ net103 net110 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_79_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_12.mux_l3_in_1_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_1_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_4_ net34 net32 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__350__A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_290_ net7 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_3__426 VGND VGND VPWR VPWR net426 cbx_1__1_.mux_top_ipin_14.mux_l2_in_3__426/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_21.mux_l2_in_1_ net71 sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_2_ net25 sb_1__1_.mux_left_track_37.out cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l1_in_1__A0 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_0__A0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__260__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_11.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_49_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_37_prog_clk
+ sb_1__1_.mem_bottom_track_13.mem_out\[0\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_2.mux_l3_in_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_right_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_2__A0 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_8.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_0.mux_l2_in_3__409 VGND VGND VPWR VPWR net409 sb_1__1_.mux_top_track_0.mux_l2_in_3__409/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_3__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_2__S sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input118_A chany_top_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_0.mux_l2_in_3__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_342_ net88 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
X_273_ net51 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input83_A chany_bottom_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_12.mux_l2_in_2_ net10 net12 sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk
+ sb_1__1_.mem_bottom_track_37.ccff_tail net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mux_left_track_29.mux_l1_in_1__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_29.mux_l4_in_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_bottom_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_3.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_5_prog_clk cby_1__1_.mem_right_ipin_1.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput235 net235 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
Xoutput224 net224 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
Xoutput213 net213 VGND VGND VPWR VPWR chanx_right_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput202 net202 VGND VGND VPWR VPWR chanx_right_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput257 net257 VGND VGND VPWR VPWR chany_top_out_0[20] sky130_fd_sc_hd__buf_12
Xoutput246 net246 VGND VGND VPWR VPWR chany_top_out_0[10] sky130_fd_sc_hd__buf_12
Xoutput268 net268 VGND VGND VPWR VPWR chany_top_out_0[3] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_3__S sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput279 net279 VGND VGND VPWR VPWR reset_left_out sky130_fd_sc_hd__buf_12
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_21.mux_l1_in_2_ net75 net55 sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_82_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_1__A0 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_2.mux_l2_in_1_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_51_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_2.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_8.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
X_325_ net102 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output287_A net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_256_ net62 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_2__S sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_3__325 VGND VGND VPWR VPWR net325 cby_1__1_.mux_right_ipin_7.mux_l2_in_3__325/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__374
+ VGND VGND VPWR VPWR net374 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__374/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_0.mux_l1_in_0_ net142 net147 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net304 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_29.mux_l3_in_1_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_bottom_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input46_A chanx_right_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_11.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_3__428 VGND VGND VPWR VPWR net428 cbx_1__1_.mux_top_ipin_2.mux_l2_in_3__428/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_75_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_308_ net104 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l2_in_2__A1 sb_1__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_2.mux_l1_in_2_ net136 net133 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_25_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_2_ net26 cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_0__A0 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_25_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input100_A chany_top_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_3.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_86_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l2_in_2__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__366
+ VGND VGND VPWR VPWR net366 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__366/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_3__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__348__A net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_2_ net31 net9 sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_80_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_1__A0 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput102 chany_top_in_0[18] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_4
XFILLER_88_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input148_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput113 chany_top_in_0[28] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput135 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND VGND VPWR
+ VPWR net135 sky130_fd_sc_hd__clkbuf_2
Xinput124 prog_reset_left_in VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput146 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND VGND VPWR
+ VPWR net146 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_2__A0 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__258__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_12.mux_l3_in_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_3_ sb_1__1_.mux_left_track_29.out net9 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_50_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_3__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_58_prog_clk cby_1__1_.mem_right_ipin_4.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_21.mux_l2_in_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_41_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_left_track_37.mux_l1_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_1_ net5 cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l1_in_1__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_0__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_16_prog_clk sb_1__1_.mem_left_track_11.ccff_head
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net372 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_40_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_40_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_40_prog_clk
+ sb_1__1_.mem_bottom_track_11.ccff_tail net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_2__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_0_prog_clk cbx_1__1_.mem_top_ipin_12.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_5.mux_l2_in_1__A0 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_41_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_58_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_341_ sb_1__1_.mux_top_track_52.out VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_272_ sb_1__1_.mux_left_track_11.out VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_12.mux_l2_in_1_ net86 sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input76_A chany_bottom_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_29.mux_l1_in_1__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_14.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__369
+ VGND VGND VPWR VPWR net369 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__369/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_32_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput214 net214 VGND VGND VPWR VPWR chanx_right_out_0[9] sky130_fd_sc_hd__buf_12
Xoutput225 net225 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
Xoutput203 net203 VGND VGND VPWR VPWR chanx_right_out_0[26] sky130_fd_sc_hd__buf_12
Xoutput247 net247 VGND VGND VPWR VPWR chany_top_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput258 net258 VGND VGND VPWR VPWR chany_top_out_0[21] sky130_fd_sc_hd__buf_12
Xoutput236 net236 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
Xoutput269 net269 VGND VGND VPWR VPWR chany_top_out_0[4] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_left_track_21.mux_l1_in_1_ net41 net115 sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_67_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_3.mux_l1_in_2_ net46 net15 cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_82_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net338 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA__356__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_8_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_2.mux_l2_in_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_2_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_2.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input130_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_8.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__266__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_324_ net101 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
X_255_ sb_1__1_.mux_left_track_45.out VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_3_ net314 net115 cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_12.mux_l1_in_2_ net72 net56 sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_29.mux_l3_in_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_2.mux_l2_in_3__A1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_2__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input39_A chanx_right_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_11.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_86_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_307_ sb_1__1_.mux_right_track_0.out VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_1__A0 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_2.mux_l1_in_1_ net130 net122 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_25_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_4.mux_l2_in_2__A0 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_0__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk cby_1__1_.mem_right_ipin_7.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l2_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_2__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_4_ sb_1__1_.mux_bottom_track_45.out net90 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__335
+ VGND VGND VPWR VPWR net335 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__335/LO
+ sky130_fd_sc_hd__conb_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_4__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_15.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_left_track_45.mux_l1_in_1__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_1_ net281 net44 sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_1__A1 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput125 prog_reset_top_in VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
Xinput114 chany_top_in_0[29] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput103 chany_top_in_0[19] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_4
Xinput136 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND VGND VPWR
+ VPWR net136 sky130_fd_sc_hd__clkbuf_2
Xinput147 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND VGND VPWR
+ VPWR net147 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_2__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__274__A sb_1__1_.mux_left_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.mux_l4_in_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_94_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_2_ net47 net16 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_31_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_58_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__359__A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_37.mux_l1_in_1__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in net138 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_sb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l2_in_1__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__269__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input21_A chanx_left_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_55_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_3_ net319 net122 cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_1__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l2_in_2__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_340_ net86 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_271_ sb_1__1_.mux_left_track_13.out VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_10.mux_l3_in_1_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_1.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_12.mux_l2_in_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_input69_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net304 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_14.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xoutput226 net226 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
Xoutput215 net215 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
Xoutput204 net204 VGND VGND VPWR VPWR chanx_right_out_0[27] sky130_fd_sc_hd__buf_12
Xoutput259 net259 VGND VGND VPWR VPWR chany_top_out_0[22] sky130_fd_sc_hd__buf_12
Xoutput248 net248 VGND VGND VPWR VPWR chany_top_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput237 net237 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
XFILLER_87_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_21.mux_l1_in_0_ net101 net105 sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_2__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_3.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_11_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__372__A net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l2_in_3__A1 net300 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_19_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_0.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input123_A prog_reset_bottom_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_323_ sb_1__1_.mux_bottom_track_29.out VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_2
X_254_ net60 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__282__A net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_3_ net426 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_89_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_1__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_45.mux_l3_in_0_ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_2_ net74 cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__333
+ VGND VGND VPWR VPWR net333 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__333/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_68_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_12.mux_l1_in_1_ net40 net42 sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_2__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcby_1__1_.mux_right_ipin_15.mux_l4_in_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.ccff_tail VGND
+ VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_74_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__277__A sb_1__1_.mux_left_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l2_in_1__A0 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_306_ sb_1__1_.mux_right_track_2.out VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__347
+ VGND VGND VPWR VPWR net347 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__347/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_40_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_53.mux_l1_in_1__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_1__A1 net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_2.mux_l1_in_0_ net108 net114 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_12.mux_l2_in_3__411 VGND VGND VPWR VPWR net411 sb_1__1_.mux_top_track_12.mux_l2_in_3__411/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_4.mux_l2_in_2__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_4_ net34 net32 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_1__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_3__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_34_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_45.mux_l2_in_1_ net394 sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_45.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input51_A chanx_right_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_2__S sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_2__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_3_ net98 net67 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_21_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__355
+ VGND VGND VPWR VPWR net355 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__355/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_45.mux_l1_in_1__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_15.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_53_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_60_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_14.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_15.mux_l3_in_1_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA__380__A net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput104 chany_top_in_0[1] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_4
Xinput115 chany_top_in_0[2] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_4
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput126 reset_bottom_in VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_12
Xinput137 sc_in VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
Xinput148 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND VGND VPWR
+ VPWR net148 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input99_A chany_top_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__290__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_4.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_1__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.out sky130_fd_sc_hd__clkbuf_2
XFILLER_62_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_37.mux_l2_in_1__382 VGND VGND VPWR VPWR net382 sb_1__1_.mux_bottom_track_37.mux_l2_in_1__382/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_6.mux_l2_in_2__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_45.mux_l1_in_2_ net297 net91 sb_1__1_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_53_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__375__A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input14_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_29.mux_l1_in_1_ net39 net52 sb_1__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_67_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_14.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_2_ net91 net99 cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ sb_1__1_.mem_bottom_track_37.mem_out\[1\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_37.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ net149 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_0__A0 sb_1__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net354 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__mux2_4
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input6_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l2_in_2__A0 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_270_ net48 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_10.mux_l3_in_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_22_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l2_in_3__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_13_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_0.ccff_tail
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xoutput216 net216 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xoutput205 net205 VGND VGND VPWR VPWR chanx_right_out_0[28] sky130_fd_sc_hd__buf_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput249 net249 VGND VGND VPWR VPWR chany_top_out_0[13] sky130_fd_sc_hd__buf_12
Xoutput227 net227 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
Xoutput238 net238 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_2__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_3.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_95_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_3_ net322 net115 cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_59_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_59_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__359
+ VGND VGND VPWR VPWR net359 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__359/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input116_A chany_top_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_322_ net99 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_253_ net59 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input81_A chany_bottom_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_2_ net26 cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_1__A1 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_1_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_12.mux_l1_in_0_ net145 net147 sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_2__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__383__A net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_3__A0 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_10.ccff_tail
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_1__S sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net374 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_305_ sb_1__1_.mux_right_track_4.out VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_11_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_7.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_69_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_53.mux_l1_in_1__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_4_ sb_1__1_.mux_bottom_track_45.out net90 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_4_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_top_track_36.mux_l3_in_0_ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l2_in_1__A0 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_50_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_3_ sb_1__1_.mux_left_track_29.out net9 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_43_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_1__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__370
+ VGND VGND VPWR VPWR net370 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__370/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_left_track_45.mux_l2_in_0_ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_4__A0 sb_1__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_1__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input44_A chanx_right_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__288__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_4.mux_l4_in_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_2_ sb_1__1_.mux_bottom_track_21.out net73 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_51_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net328 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l2_in_2__A0 net297 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_15.mux_l3_in_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_0__A0 sb_1__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput105 chany_top_in_0[20] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput116 chany_top_in_0[3] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_4
Xinput127 reset_right_in VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
Xinput149 top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput138 test_enable_bottom_in VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_12
XFILLER_29_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_3__A1 net282 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_79_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_36.mux_l2_in_1_ net415 sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.out sky130_fd_sc_hd__buf_4
XFILLER_79_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_1__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net138 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_3_ net327 net119 cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_89_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_3.ccff_tail
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_2__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_45.mux_l1_in_1_ net67 net37 sb_1__1_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_4__A0 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input146_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_4.mux_l3_in_1_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__348
+ VGND VGND VPWR VPWR net348 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__348/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_29.mux_l1_in_0_ net104 net99 sb_1__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_11.ccff_tail
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_1_ net68 cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_14.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_94_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ sb_1__1_.mem_bottom_track_37.mem_out\[0\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_37.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_3__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l2_in_2__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_36.mux_l1_in_2_ net8 net20 sb_1__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_top_track_6.mux_l2_in_3_ net419 net29 sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_4__S sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net126 net137 net138 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk cby_1__1_.mem_right_ipin_13.ccff_tail
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_1_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XANTENNA__296__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l2_in_1__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput217 net217 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
Xoutput206 net206 VGND VGND VPWR VPWR chanx_right_out_0[29] sky130_fd_sc_hd__buf_12
Xoutput239 net239 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
Xoutput228 net228 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
XFILLER_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_2_ net74 cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_3__A1 net295 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_28_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input109_A chany_top_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_321_ net98 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_252_ net58 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_9.mux_l4_in_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_22_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input74_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_15.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.out sky130_fd_sc_hd__buf_4
XFILLER_77_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_40_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_6.mux_l1_in_4_ net16 net89 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_2__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_3__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_11.mux_l2_in_3__388 VGND VGND VPWR VPWR net388 sb_1__1_.mux_left_track_11.mux_l2_in_3__388/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_304_ sb_1__1_.mux_right_track_6.out VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_7_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_3_ net98 net67 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_3__318 VGND VGND VPWR VPWR net318 cby_1__1_.mux_right_ipin_14.mux_l2_in_3__318/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_45_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_6.mux_l4_in_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_6.ccff_tail
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_9.mux_l3_in_1_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_2_ net47 net16 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_4__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input37_A chanx_right_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_43_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_14.ccff_tail
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l2_in_3__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput106 chany_top_in_0[21] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_4
Xinput117 chany_top_in_0[4] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput139 test_enable_right_in VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
Xinput128 reset_top_in VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_28.mux_l2_in_1__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_36.mux_l2_in_0_ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA__299__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_6.mux_l3_in_1_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_0.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_28.mux_l2_in_3_ net403 net14 sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_2_ net88 net99 cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l2_in_3__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_2__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_45.mux_l1_in_0_ net97 net112 sb_1__1_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_42_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_3__424 VGND VGND VPWR VPWR net424 cbx_1__1_.mux_top_ipin_12.mux_l2_in_3__424/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_4__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_3__312 VGND VGND VPWR VPWR net312 cby_1__1_.mux_right_ipin_0.mux_l2_in_3__312/LO
+ sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_4.mux_l3_in_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input139_A test_enable_right_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_94_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ sb_1__1_.mem_bottom_track_29.ccff_tail net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_90_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_2__S cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_0__A0 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_3_ net378 net26 sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_36.mux_l1_in_1_ net68 net57 sb_1__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk cbx_1__1_.mem_top_ipin_0.ccff_tail
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_top_track_6.mux_l2_in_2_ net31 sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_top_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l2_in_2__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_30_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net336 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__mux2_2
Xoutput207 net207 VGND VGND VPWR VPWR chanx_right_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput229 net229 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
Xoutput218 net218 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
XFILLER_4_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_6.mux_l2_in_3__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net363 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_1_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l1_in_2__A0 net281 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_right_track_28.mux_l4_in_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_right_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_320_ net97 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_12.mux_l1_in_2__A0 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_251_ sb_1__1_.mux_left_track_53.out VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_36.mux_l1_in_2__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_15.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input67_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l2_in_3__A1 sb_1__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_6.mux_l1_in_3_ net76 net59 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_3__323 VGND VGND VPWR VPWR net323 cby_1__1_.mux_right_ipin_5.mux_l2_in_3__323/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input121_A chany_top_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_303_ net21 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_2__A0 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_4__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_bottom_track_13.mux_l4_in_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_2_ sb_1__1_.mux_bottom_track_21.out net73 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_80_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_21.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_12.mux_l2_in_1__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_28.mux_l3_in_1_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_right_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_9.mux_l3_in_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_56_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l2_in_2__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_12_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_4__A0 net296 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_53.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net346 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.out sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xinput107 chany_top_in_0[22] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_4
Xinput118 chany_top_in_0[5] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_4
Xinput129 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND VGND VPWR
+ VPWR net129 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_1__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_56_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_28.mux_l2_in_1__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_13.mux_l3_in_1_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_3.ccff_tail
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_4_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_6.mux_l3_in_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_0.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_28.mux_l2_in_2_ net9 net74 sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_43_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_1_ net68 cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_20_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input97_A chany_top_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__337
+ VGND VGND VPWR VPWR net337 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__337/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_75_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_3__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_0__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_2_ net10 net12 sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_85_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_3__A0 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l1_in_1__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l1_in_2__A0 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_2__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_36.mux_l1_in_0_ net38 net142 sb_1__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_6.mux_l2_in_1_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l2_in_2__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input12_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_9.mux_l1_in_2_ net106 net75 cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_60_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xoutput208 net208 VGND VGND VPWR VPWR chanx_right_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput219 net219 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l2_in_2__A0 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_36.mux_l2_in_1__415 VGND VGND VPWR VPWR net415 sb_1__1_.mux_top_track_36.mux_l2_in_1__415/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_6.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l1_in_2__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_3_ net306 net55 cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_2__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_12.mux_l1_in_2__A1 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_250_ net56 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_top_track_36.mux_l1_in_2__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_15.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_37_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_37_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l2_in_2__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_1__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_379_ net138 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_3_ net384 net30 sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_68_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_20.mux_l2_in_3__402 VGND VGND VPWR VPWR net402 sb_1__1_.mux_right_track_20.mux_l2_in_3__402/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_6.mux_l1_in_2_ net46 net49 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__360
+ VGND VGND VPWR VPWR net360 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__360/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input114_A chany_top_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_302_ sb_1__1_.mux_right_track_10.out VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_2__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_4__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_6.ccff_tail
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_92_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_21.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__356
+ VGND VGND VPWR VPWR net356 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__356/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_81_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk sb_1__1_.mem_left_track_5.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_4_ sb_1__1_.mux_left_track_45.out net30 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_21.mux_l2_in_1__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_28.mux_l3_in_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_29_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_3__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_52_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_52_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output283_A net283 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_4__A1 net294 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_53.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_53.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l2_in_3__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput108 chany_top_in_0[23] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput119 chany_top_in_0[6] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_4
XANTENNA_sb_1__1_.mux_right_track_10.mux_l2_in_3__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_56_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_10_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_13.mux_l3_in_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__329
+ VGND VGND VPWR VPWR net329 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__329/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_79_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_5.mux_l4_in_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_input42_A chanx_right_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_27_prog_clk sb_1__1_.mem_top_track_0.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_2__A0 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_28.mux_l2_in_1_ net69 net82 sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_43_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_1__A0 net282 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_2__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_3_ net311 net59 cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_19_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput90 chany_bottom_in[7] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_4
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ sb_1__1_.mem_bottom_track_29.mem_out\[2\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_11.mux_l2_in_3__A1 net300 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_4.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_40_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_0__A0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_1_ net285 sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_3__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l1_in_1__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_20.mux_l1_in_2__A1 net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_2__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_5.mux_l3_in_1_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_6.mux_l2_in_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input144_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__340
+ VGND VGND VPWR VPWR net340 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__340/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_9.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_25_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_20.mux_l2_in_3_ net413 net25 sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xoutput209 net209 VGND VGND VPWR VPWR chanx_right_out_0[4] sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l2_in_2__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
XFILLER_63_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_7_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_6.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_2_ net14 cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_2__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_89_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_9.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_378_ net152 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_1__1_.mux_bottom_track_13.mux_l1_in_2_ net287 net56 sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_2_ net17 net20 sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_6.mux_l1_in_1_ net145 net143 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_38_prog_clk sb_1__1_.mem_bottom_track_1.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_36_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input107_A chany_top_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_301_ sb_1__1_.mux_right_track_12.out VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input72_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_37_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk sb_1__1_.mem_left_track_21.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_3__311 VGND VGND VPWR VPWR net311 cbx_1__1_.mux_top_ipin_9.mux_l2_in_3__311/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_5.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_3_ net38 net7 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in net138 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_68_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_20.mux_l4_in_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net344 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_9.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_1__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_1__A0 net283 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_5.mux_l2_in_3_ net395 net298 sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_21_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_21_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_45.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net364 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xinput109 chany_top_in_0[24] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input35_A chanx_right_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_28_prog_clk net2
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_2__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_28.mux_l2_in_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_1__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_2__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_20.mux_l3_in_1_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__363
+ VGND VGND VPWR VPWR net363 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__363/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_38_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_2_ net28 net39 cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_93_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_3__A0 net283 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net335 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__352
+ VGND VGND VPWR VPWR net352 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__352/LO
+ sky130_fd_sc_hd__conb_1
Xinput80 chany_bottom_in[25] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_4
Xinput91 chany_bottom_in[8] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ sb_1__1_.mem_bottom_track_29.mem_out\[1\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_4.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_0__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_3__308 VGND VGND VPWR VPWR net308 cbx_1__1_.mux_top_ipin_6.mux_l2_in_3__308/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__310__A net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_2__S sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_5.mux_l3_in_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_5.mux_l4_in_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_right_track_28.mux_l1_in_1_ net131 net104 sb_1__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_94_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input137_A sc_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_9.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_45_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_20.mux_l2_in_2_ net11 net15 sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l2_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_27_prog_clk sb_1__1_.mem_top_track_6.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net373 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__mux2_2
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_3__A0 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_46_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_377_ net126 VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_13.mux_l1_in_1_ net42 net49 sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_0__A0 net143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_1_ net284 sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_5.mux_l3_in_1_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_95_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_6.mux_l1_in_0_ net141 net147 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_37_prog_clk sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_91_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_300_ net18 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input65_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_13.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_73_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_2__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_10.mux_l2_in_3__410 VGND VGND VPWR VPWR net410 sb_1__1_.mux_top_track_10.mux_l2_in_3__410/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_5.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_2_ sb_1__1_.mux_left_track_21.out net13 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_2__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput1 ccff_head_1 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l2_in_2__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_9.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_86_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_5.mux_l1_in_2_ net281 net60 sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_1__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_5.mux_l2_in_2_ net295 net90 sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_51_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_61_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_61_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__364
+ VGND VGND VPWR VPWR net364 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__364/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_3_ net315 sb_1__1_.mux_bottom_track_53.out
+ cby_1__1_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_4__A0 sb_1__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__313__A net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_1__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_42_prog_clk sb_1__1_.mem_bottom_track_7.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput190 net190 VGND VGND VPWR VPWR chanx_right_out_0[14] sky130_fd_sc_hd__buf_12
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input28_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_20.mux_l3_in_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_1_ net8 cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__308__A net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_3__A1 net281 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput70 chany_bottom_in[16] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
Xinput81 chany_bottom_in[26] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_4
XANTENNA_cby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk
+ sb_1__1_.mem_bottom_track_29.mem_out\[0\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput92 chany_bottom_in[9] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_4
XFILLER_1_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_3_ net422 net55 cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_48_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_2__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_28.mux_l1_in_0_ net99 net100 sb_1__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_11.mux_l4_in_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_43_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input95_A chany_top_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_0__A0 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_20.mux_l2_in_1_ net85 sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_9.mux_l1_in_2_ net46 net15 cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_68_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_4.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mux_left_track_21.mux_l2_in_3__390 VGND VGND VPWR VPWR net390 sb_1__1_.mux_left_track_21.mux_l2_in_3__390/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_31_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__321__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_73_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_4__A0 sb_1__1_.mux_left_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_10.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_3__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_4_ sb_1__1_.mux_left_track_45.out net30 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input10_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_15_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_15_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
X_376_ net126 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net333 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_13.mux_l1_in_0_ net116 net102 sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_output299_A net299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_2__A0 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_5.mux_l3_in_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_39_prog_clk sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__316__A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_11.mux_l3_in_1_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input2_A ccff_head_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_20.mux_l1_in_2_ net71 net55 sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_53.mux_l1_in_1__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_37.mux_l3_in_0_ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input58_A chanx_right_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net138 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_2__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_3.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_359_ net77 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_3__316 VGND VGND VPWR VPWR net316 cby_1__1_.mux_right_ipin_12.mux_l2_in_3__316/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_2__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ net152 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xinput2 ccff_head_2 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.out sky130_fd_sc_hd__buf_4
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_3_ net427 net62 cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_input112_A chany_top_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_5.mux_l1_in_1_ net36 net47 sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_5.mux_l2_in_1_ net77 sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.out sky130_fd_sc_hd__buf_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_30_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_2_ net86 net97 cby_1__1_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_4__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__342
+ VGND VGND VPWR VPWR net342 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__342/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_84_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_37.mux_l2_in_1_ net382 sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in net138 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_42_prog_clk sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xoutput191 net191 VGND VGND VPWR VPWR chanx_right_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput180 net180 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output281_A net281 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_3__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__324__A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput82 chany_bottom_in[27] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
Xinput71 chany_bottom_in[17] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_4
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ sb_1__1_.mem_bottom_track_21.ccff_tail net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput60 chanx_right_in_0[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
Xinput93 chany_top_in_0[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlymetal6s2s_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net353 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_3_ net312 net119 cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_3__422 VGND VGND VPWR VPWR net422 cbx_1__1_.mux_top_ipin_10.mux_l2_in_3__422/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_84_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_5.mux_l1_in_2_ net83 net60 sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input40_A chanx_right_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l2_in_3__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_2_ net14 cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_37.mux_l1_in_2_ net27 net8 sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_15.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X net154 VGND VGND VPWR VPWR
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_59_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_44.mux_l2_in_1__406 VGND VGND VPWR VPWR net406 sb_1__1_.mux_right_track_44.mux_l2_in_1__406/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__319__A sb_1__1_.mux_bottom_track_37.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_33_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_89_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_2__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_0.mux_l2_in_2__A0 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_0__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_20.mux_l2_in_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_input88_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_9.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_3__378 VGND VGND VPWR VPWR net378 sb_1__1_.mux_bottom_track_13.mux_l2_in_3__378/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_12.mux_l2_in_3_ net400 net26 sb_1__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_3__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_4_ sb_1__1_.mux_bottom_track_37.out net65 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_10.mux_l2_in_3__399 VGND VGND VPWR VPWR net399 sb_1__1_.mux_right_track_10.mux_l2_in_3__399/LO
+ sky130_fd_sc_hd__conb_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_10.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l1_in_2__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_3_ net38 net7 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input142_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_375_ net126 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
XFILLER_70_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_55_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__1_.mux_top_ipin_15.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_5_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_0.mux_l4_in_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_2__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_53.mux_l3_in_0_ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.ccff_head VGND
+ VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_41_prog_clk sb_1__1_.mem_bottom_track_1.ccff_head
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net355 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__mux2_4
XFILLER_91_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__332__A sb_1__1_.mux_bottom_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_13.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.mux_l3_in_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_86_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_20.mux_l1_in_1_ net36 net41 sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_3__321 VGND VGND VPWR VPWR net321 cby_1__1_.mux_right_ipin_3.mux_l2_in_3__321/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_67_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_358_ net76 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l2_in_1__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_289_ sb_1__1_.mux_right_track_36.out VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_3_ net323 net104 cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_83_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput3 chanx_left_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_45.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_0_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_12.mux_l4_in_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_86_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_2_ net31 net39 cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A chany_top_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_0.mux_l3_in_1_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_5.mux_l1_in_0_ net120 net107 sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_5.mux_l2_in_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_1__A1 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_53.mux_l2_in_1_ net396 sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_53.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input70_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_1_ net66 cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_10.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_27_prog_clk sb_1__1_.mem_top_track_10.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_2__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_37.mux_l2_in_0_ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_37_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_42_prog_clk sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xoutput170 net170 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
Xoutput192 net192 VGND VGND VPWR VPWR chanx_right_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput181 net181 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_2.mux_l2_in_3_ net412 net3 sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_12_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_3__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_49_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_12.mux_l3_in_1_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xinput50 chanx_right_in_0[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput72 chany_bottom_in[18] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_4
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_2__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput61 chanx_right_in_0[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput94 chany_top_in_0[10] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_4
Xinput83 chany_bottom_in[28] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
XANTENNA__340__A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_2_ net88 cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_5.mux_l1_in_1_ net47 net117 sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_53.mux_l1_in_2_ net298 net87 sb_1__1_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_4__A0 sb_1__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_right_track_28.mux_l1_in_0__A0 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_5.mux_l4_in_0_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA__250__A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.mux_l1_in_2_ net103 net72 cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input33_A chanx_right_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_75_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_1__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_37.mux_l1_in_1_ net282 net38 sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_5_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_33_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__335__A sb_1__1_.mux_bottom_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_0.mux_l2_in_2__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_9.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_4_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_29.mux_l1_in_0__A0 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_right_track_12.mux_l2_in_2_ net12 net86 sb_1__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_75_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_right_track_0.mux_l2_in_3__398 VGND VGND VPWR VPWR net398 sb_1__1_.mux_right_track_0.mux_l2_in_3__398/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net304 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_3__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_3_ net102 net71 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_11.mux_l2_in_3_ net388 net300 sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_2.mux_l4_in_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_10.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l1_in_2__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_5.mux_l3_in_1_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_2_ sb_1__1_.mux_left_track_21.out net13 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_4__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input135_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_374_ net126 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_15.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_24_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_53.mux_l2_in_1__385 VGND VGND VPWR VPWR net385 sb_1__1_.mux_bottom_track_53.mux_l2_in_1__385/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_13.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_2__A0 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_20.mux_l1_in_0_ net146 net148 sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_top_track_2.mux_l2_in_2__A0 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.mux_l1_in_4_ net296 net294 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_2.mux_l3_in_1_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_top_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_60_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_357_ sb_1__1_.mux_top_track_20.out VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_288_ net5 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
XANTENNA_load_slew303_A net304 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_2_ net63 net94 cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xinput4 chanx_left_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
Xsb_1__1_.mux_top_track_44.mux_l3_in_0_ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net369 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l2_in_3__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_24_prog_clk sb_1__1_.mem_left_track_45.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_45.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__343__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_4__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_1_ net8 cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_0__S sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_0.mux_l3_in_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_42_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_11.mux_l4_in_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA__253__A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_53.mux_l2_in_0_ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input63_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_39_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net138 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_61_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_4.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_27_prog_clk sb_1__1_.mem_top_track_10.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_2__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l2_in_3__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_1__S sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__338__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_0__A0 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_42_prog_clk sb_1__1_.mem_bottom_track_5.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__331
+ VGND VGND VPWR VPWR net331 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__331/LO
+ sky130_fd_sc_hd__conb_1
Xoutput160 net160 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
Xoutput171 net171 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
Xoutput193 net193 VGND VGND VPWR VPWR chanx_right_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput182 net182 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_top_track_2.mux_l2_in_2_ net32 net18 sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_1__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__248__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_7.mux_l2_in_3__397 VGND VGND VPWR VPWR net397 sb_1__1_.mux_left_track_7.mux_l2_in_3__397/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_2__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_44.mux_l2_in_1_ net417 sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_44.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_0__S sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_12.mux_l3_in_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput40 chanx_right_in_0[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput51 chanx_right_in_0[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_4
Xinput73 chany_bottom_in[19] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_4
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_2__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput62 chanx_right_in_0[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xcbx_1__1_.mux_top_ipin_15.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xinput95 chany_top_in_0[11] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
Xinput84 chany_bottom_in[29] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_4
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_1_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net371 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_5.mux_l1_in_0_ net120 net107 sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_11.mux_l3_in_1_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_53.mux_l1_in_1_ net65 net35 sb_1__1_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_4__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_58_prog_clk cby_1__1_.mem_right_ipin_0.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_37.mux_l1_in_0__A0 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_input26_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_1__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_49_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_49_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_3__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_37.mux_l1_in_0_ net53 net98 sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_32_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_top_track_2.mux_l1_in_3_ net92 net78 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA__351__A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_0__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l2_in_1__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_44.mux_l1_in_2_ net7 net22 sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_25_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__261__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_12.mux_l2_in_1_ net72 sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_3__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net304 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_2__A0 net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__334
+ VGND VGND VPWR VPWR net334 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__334/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_left_track_11.mux_l2_in_2_ net298 sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_left_track_11.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_10.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l2_in_3__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_10.ccff_head
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__346__A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_5.mux_l3_in_0_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l2_in_2__A0 net297 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_3__S sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input128_A reset_top_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_4.mux_l1_in_2__A0 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__256__A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_373_ net126 VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input93_A chany_top_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_13.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_2__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_12.mux_l1_in_2_ net79 net135 sb_1__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_40_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_2.mux_l2_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_1__A0 net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net337 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__mux2_4
XFILLER_18_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.mux_l1_in_3_ net88 net73 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_60_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_2.mux_l3_in_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_top_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_41_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_356_ net73 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_2
XANTENNA_output297_A net297 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_287_ net4 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_1_ net92 cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 chanx_left_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_0__A0 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_37.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_32_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_4.mux_l2_in_1__A0 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_4__A1 net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_3__376 VGND VGND VPWR VPWR net376 sb_1__1_.mux_bottom_track_1.mux_l2_in_3__376/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__338
+ VGND VGND VPWR VPWR net338 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__338/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_0_prog_clk cby_1__1_.mem_right_ipin_3.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input56_A chanx_right_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_1__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_339_ net85 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_4.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_31_prog_clk sb_1__1_.mem_top_track_10.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_45.mux_l1_in_0__A0 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_0__A1 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__354__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_11.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput161 net161 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput194 net194 VGND VGND VPWR VPWR chanx_right_out_0[18] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_top_track_2.mux_l2_in_1_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_1__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input110_A chany_top_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__264__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_5.mux_l1_in_2_ net103 net72 cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_44.mux_l2_in_0_ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_44.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l2_in_3__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_45.mux_l2_in_1__394 VGND VGND VPWR VPWR net394 sb_1__1_.mux_left_track_45.mux_l2_in_1__394/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_right_track_4.mux_l2_in_3_ net405 net30 sb_1__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput30 chanx_left_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_4
Xinput52 chanx_right_in_0[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 chanx_right_in_0[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
Xinput63 chany_bottom_in[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
Xcbx_1__1_.mux_top_ipin_15.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xinput96 chany_top_in_0[12] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 chany_bottom_in[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_4
Xinput74 chany_bottom_in[1] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_4
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_13.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_11.mux_l3_in_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_53.mux_l1_in_0_ net95 net113 sb_1__1_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_57_prog_clk cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_3_ net420 net59 cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_52_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_11.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_87_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_input19_A chanx_left_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__259__A sb_1__1_.mux_left_track_37.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__346
+ VGND VGND VPWR VPWR net346 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__346/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_73_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_3__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_18_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_3__306 VGND VGND VPWR VPWR net306 cbx_1__1_.mux_top_ipin_4.mux_l2_in_3__306/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_32_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_3_ net376 net4 sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_2.mux_l1_in_2_ net62 net48 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_3_ net379 net25 sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_44.mux_l1_in_1_ net67 net33 sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_80_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_12.mux_l2_in_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l2_in_2__A0 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_2__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_11.mux_l2_in_1_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_4_ sb_1__1_.mux_left_track_37.out net5 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__350
+ VGND VGND VPWR VPWR net350 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__350/LO
+ sky130_fd_sc_hd__conb_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.out sky130_fd_sc_hd__clkbuf_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l2_in_2__A1 net294 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_4.mux_l1_in_2__A1 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_372_ net302 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_right_track_4.mux_l4_in_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input86_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__272__A sb_1__1_.mux_left_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_6.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_79_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_0__A0 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_0.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_33_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_33_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_11.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_86_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_12.mux_l1_in_1_ net129 net116 sb_1__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_14.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input140_A test_enable_top_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_1.mux_l4_in_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.mux_l1_in_2_ net80 net58 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_355_ net72 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_286_ net32 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_21.mux_l4_in_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_0_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_53.mux_l1_in_0__A0 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 chanx_left_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_0__A1 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_3_ net307 net44 cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_4.mux_l3_in_1_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_0__A0 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net366 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__mux2_2
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_0.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_2_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_0__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input49_A chanx_right_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ net74 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_269_ net47 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_10.ccff_head
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_4.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_1.mux_l3_in_1_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_bottom_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__370__A net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput151 net151 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_
+ sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_top_track_2.mux_l2_in_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xoutput173 net173 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
Xoutput162 net162 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
Xoutput195 net195 VGND VGND VPWR VPWR chanx_right_out_0[19] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.out sky130_fd_sc_hd__buf_4
Xoutput184 net184 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
XFILLER_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_2.mux_l2_in_3__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__358
+ VGND VGND VPWR VPWR net358 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__358/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input103_A chany_top_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_21.mux_l3_in_1_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_43_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_5.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__280__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_2__A0 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_0__A0 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_20_prog_clk cbx_1__1_.mem_top_ipin_0.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_19_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_4.mux_l2_in_2_ net17 net90 sb_1__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xinput31 chanx_left_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
Xinput20 chanx_left_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xinput53 chanx_right_in_0[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput42 chanx_right_in_0[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xcbx_1__1_.mux_top_ipin_15.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xinput64 chany_bottom_in[10] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_4
Xinput97 chany_top_in_0[13] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_2
XFILLER_6_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput75 chany_bottom_in[20] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
Xinput86 chany_bottom_in[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_4
XANTENNA_cby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_57_prog_clk cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_37_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_2_ net28 cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net350 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_6.mux_l2_in_3__419 VGND VGND VPWR VPWR net419 sb_1__1_.mux_top_track_6.mux_l2_in_3__419/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__345
+ VGND VGND VPWR VPWR net345 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__345/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_5.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_58_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_58_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk cby_1__1_.mem_right_ipin_9.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_32_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_2_ net21 net23 sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_2.mux_l1_in_1_ net52 net146 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_2_ net6 net11 sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_2__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_44.mux_l1_in_0_ net37 net143 sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_48_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input31_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_0__S sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l2_in_2__A1 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.mux_l2_in_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_3_ net42 net11 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_5.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_3_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_3_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l1_in_1__A0 sb_1__1_.mux_left_track_11.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_2__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_371_ net302 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input79_A chany_bottom_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_0__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_3_ net285 net282 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l2_in_3_ net387 net299 sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_12.mux_l1_in_0_ net102 net109 sb_1__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_10_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__373__A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_2__A0 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_56_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input133_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.mux_l1_in_1_ net43 net118 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_354_ net71 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__283__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_285_ sb_1__1_.mux_right_track_44.out VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_3__314 VGND VGND VPWR VPWR net314 cby_1__1_.mux_right_ipin_10.mux_l2_in_3__314/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput7 chanx_left_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_4
XFILLER_76_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_3.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_51_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_2_ net3 net34 cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xoutput300 net300 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_7_ sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_right_track_36.mux_l3_in_0_ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_4.mux_l3_in_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_59_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__368__A net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_0__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_0.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_3__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_52.mux_l2_in_1__418 VGND VGND VPWR VPWR net418 sb_1__1_.mux_top_track_52.mux_l2_in_1__418/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_76_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__278__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_0_prog_clk net432 net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_337_ sb_1__1_.mux_bottom_track_1.out VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_2
X_268_ net46 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l2_in_2__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_2.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_load_slew301_A net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l2_in_2__A0 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_1.mux_l3_in_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_bottom_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_left_track_1.mux_l4_in_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput152 net152 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ sky130_fd_sc_hd__buf_12
Xoutput174 net174 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chanx_right_out_0[0] sky130_fd_sc_hd__buf_12
Xoutput196 net196 VGND VGND VPWR VPWR chanx_right_out_0[1] sky130_fd_sc_hd__buf_12
XFILLER_87_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xsb_1__1_.mux_bottom_track_21.mux_l3_in_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_30_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_5.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_11_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_2__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input61_A chanx_right_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_3__S sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_36.mux_l2_in_1_ net404 sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_4.mux_l2_in_1_ net66 sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xinput10 chanx_left_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
Xinput21 chanx_left_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
Xinput54 chanx_right_in_0[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 chanx_right_in_0[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
Xinput32 chanx_left_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
Xinput98 chany_top_in_0[14] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_4
Xinput87 chany_bottom_in[4] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
Xinput76 chany_bottom_in[21] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_4
Xinput65 chany_bottom_in[11] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_4
XANTENNA_sb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_59_prog_clk net1
+ net123 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_1__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_38_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__381__A net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_3__421 VGND VGND VPWR VPWR net421 cbx_1__1_.mux_top_ipin_1.mux_l2_in_3__421/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_3__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__291__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_9.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_27_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_33_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_1_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l3_in_1_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_left_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_2.mux_l1_in_0_ net143 net148 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_1_ net286 sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_2__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net138 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__sdfrtp_2
XANTENNA__376__A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_3__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_36.mux_l1_in_2_ net8 net68 sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_68_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_4.mux_l1_in_2_ net77 net134 sb_1__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input24_A chanx_left_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__286__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_10.ccff_head
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l2_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_6.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_5.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_2__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_370_ net303 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_2_ net287 net57 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_28.mux_l2_in_3__403 VGND VGND VPWR VPWR net403 sb_1__1_.mux_right_track_28.mux_l2_in_3__403/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_left_track_1.mux_l2_in_2_ net296 net293 sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_68_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l1_in_2__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_21.mux_l1_in_2_ net288 net55 sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in net138 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_3__427 VGND VGND VPWR VPWR net427 cbx_1__1_.mux_top_ipin_15.mux_l2_in_3__427/LO
+ sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_42_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_42_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_5__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_2__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_56_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_24_prog_clk sb_1__1_.mem_left_track_37.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_11.mux_l1_in_0_ net96 net103 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input126_A reset_bottom_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_353_ sb_1__1_.mux_top_track_28.out VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input91_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_284_ net30 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_28.mux_l1_in_1__A0 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 chanx_left_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_4
Xsb_1__1_.mux_right_track_6.mux_l2_in_3__408 VGND VGND VPWR VPWR net408 sb_1__1_.mux_right_track_6.mux_l2_in_3__408/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_64_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_1_ net32 cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_2.ccff_tail
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_left_track_1.mux_l1_in_3_ net63 net64 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l2_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_3__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_2__S sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__294__A net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_336_ sb_1__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_2
XANTENNA_output295_A net295 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_267_ sb_1__1_.mux_left_track_21.out VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net339 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_28_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net348 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__mux2_4
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l2_in_2__A1 sb_1__1_.mux_left_track_37.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_10.ccff_tail
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput175 net175 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
Xoutput186 net186 VGND VGND VPWR VPWR chanx_right_out_0[10] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
XFILLER_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput197 net197 VGND VGND VPWR VPWR chanx_right_out_0[20] sky130_fd_sc_hd__buf_12
XFILLER_75_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__379__A net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input54_A chanx_right_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_5.mux_l1_in_2_ net43 net12 cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_93_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_36.mux_l2_in_0_ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_4.mux_l2_in_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_319_ sb_1__1_.mux_bottom_track_37.out VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
Xinput11 chanx_left_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_4
Xinput22 chanx_left_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
Xinput33 chanx_right_in_0[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput44 chanx_right_in_0[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xinput55 chanx_right_in_0[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xinput66 chany_bottom_in[12] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
Xinput77 chany_bottom_in[22] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_4
Xinput88 chany_bottom_in[5] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_4
Xinput99 chany_top_in_0[15] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_2
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_3__326 VGND VGND VPWR VPWR net326 cby_1__1_.mux_right_ipin_8.mux_l2_in_3__326/LO
+ sky130_fd_sc_hd__conb_1
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_43_prog_clk cby_1__1_.mem_right_ipin_12.ccff_tail
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_52_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_9.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_3__A1 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_3_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_3_ net316 net119 cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_41_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l3_in_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_left_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__367
+ VGND VGND VPWR VPWR net367 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__367/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_right_track_36.mux_l1_in_1_ net83 net132 sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_88_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_4.mux_l1_in_1_ net131 net120 sb_1__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l2_in_1__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_3__377 VGND VGND VPWR VPWR net377 sb_1__1_.mux_bottom_track_11.mux_l2_in_3__377/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input17_A chanx_left_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_94_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_4_ sb_1__1_.mux_bottom_track_37.out net65 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_3_ net423 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_36.mux_l1_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_5.ccff_tail
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_1_ net34 net51 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_79_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_1.mux_l2_in_1_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net334 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l1_in_2__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_21.mux_l1_in_1_ net41 net50 sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l2_in_2__A1 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_11_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_12.mux_l4_in_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_13.ccff_tail
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_23_prog_clk sb_1__1_.mem_left_track_37.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_37.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input119_A chany_top_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_3__A0 net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_352_ net69 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_283_ net29 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input84_A chany_bottom_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_1__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_3__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput9 chanx_left_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XFILLER_64_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_18_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_32_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_0__S cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_57_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_1.mux_l1_in_2_ net81 net34 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_335_ sb_1__1_.mux_bottom_track_5.out VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_266_ net43 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
XANTENNA_output288_A net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_3__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_12.mux_l3_in_1_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_60_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l2_in_2__A0 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xoutput176 net176 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xoutput165 net165 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
Xoutput187 net187 VGND VGND VPWR VPWR chanx_right_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput198 net198 VGND VGND VPWR VPWR chanx_right_out_0[21] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__1_.mux_right_track_10.mux_l2_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_34_prog_clk sb_1__1_.mem_right_track_20.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_5.mux_l2_in_3__395 VGND VGND VPWR VPWR net395 sb_1__1_.mux_left_track_5.mux_l2_in_3__395/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input47_A chanx_right_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_5.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_93_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_8_prog_clk cbx_1__1_.ccff_head
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_318_ net95 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
Xinput12 chanx_left_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_4
Xinput45 chanx_right_in_0[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput34 chanx_right_in_0[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_4
Xinput23 chanx_left_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
X_249_ net55 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput78 chany_bottom_in[23] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_4
Xinput89 chany_bottom_in[6] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_4
Xinput67 chany_bottom_in[13] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_4
Xinput56 chanx_right_in_0[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_2__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_9.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_75_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input101_A chany_top_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_52.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_8.ccff_tail
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_2_ net88 cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_41_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_36_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_36_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l1_in_0__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_1__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_36.mux_l1_in_0_ net96 net98 sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net123 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input149_A top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_4.mux_l1_in_0_ net107 net113 sb_1__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_48_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l2_in_1__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_3_ net313 net118 cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_50_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_3__S cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_2.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l1_in_1__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_4__A0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__328
+ VGND VGND VPWR VPWR net328 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__328/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_1__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_12.mux_l1_in_1__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_3_ net102 net71 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_2_ net26 net37 cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_21_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_top_track_36.mux_l1_in_1__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net138 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_0_ net94 net111 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l2_in_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l2_in_3__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_21.mux_l1_in_0_ net115 net101 sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_51_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk sb_1__1_.mem_left_track_29.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_351_ net68 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_3__A1 net283 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_282_ net28 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mux_bottom_track_45.mux_l3_in_0_ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_1__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_3__A1 net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input77_A chany_bottom_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_2.ccff_tail
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_3_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_1.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_1.mux_l1_in_1_ net51 net94 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_23_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input131_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_1.mux_l4_in_0_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_92_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ sb_1__1_.mux_bottom_track_7.out VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_265_ net42 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_3__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_12.mux_l3_in_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l2_in_2__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xoutput155 net155 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
Xoutput166 net166 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
Xoutput177 net177 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR chanx_right_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR chanx_right_out_0[22] sky130_fd_sc_hd__buf_12
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_45.mux_l2_in_1_ net383 sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_45.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk sb_1__1_.mem_right_track_20.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_5.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_93_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net330 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__mux2_4
XFILLER_61_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_317_ net94 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_3_ net324 net119 cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xinput13 chanx_left_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
Xinput46 chanx_right_in_0[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
Xinput35 chanx_right_in_0[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
Xinput24 chanx_left_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
X_248_ net44 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
Xinput79 chany_bottom_in[24] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
Xinput68 chany_bottom_in[14] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_4
Xinput57 chanx_right_in_0[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_0__A0 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_1__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net375 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ net153 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcby_1__1_.mux_right_ipin_1.mux_l3_in_1_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_6_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_top_track_4.mux_l2_in_3__416 VGND VGND VPWR VPWR net416 sb_1__1_.mux_top_track_4.mux_l2_in_3__416/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_28_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk sb_1__1_.mem_right_track_52.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_1_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_78_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_45.mux_l1_in_2_ net3 net7 sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__368
+ VGND VGND VPWR VPWR net368 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__368/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_2__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l1_in_0__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l1_in_1__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_1__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_4_ sb_1__1_.mux_bottom_track_37.out net65 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_29.mux_l2_in_3__391 VGND VGND VPWR VPWR net391 sb_1__1_.mux_left_track_29.mux_l2_in_3__391/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_31_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_37_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__1_.mux_right_track_20.mux_l2_in_3_ net402 net25 sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_94_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_2_ net87 net98 cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_5.ccff_tail
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_2.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_20.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_6.mux_l4_in_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_4__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_1__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_1_ net6 cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A chanx_left_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net352 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l2_in_3__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_20_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_52.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_0__A0 sb_1__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_350_ net67 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_281_ sb_1__1_.mux_right_track_52.out VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_76_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.out sky130_fd_sc_hd__clkbuf_2
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l2_in_3__A1 sb_1__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_6.mux_l3_in_1_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_1.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_11.mux_l1_in_2_ net43 net12 cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_55_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_1.mux_l1_in_0_ net111 net114 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_20.mux_l4_in_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_76_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input124_A prog_reset_left_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_333_ net111 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_2__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_264_ net41 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput167 net167 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
Xoutput189 net189 VGND VGND VPWR VPWR chanx_right_out_0[13] sky130_fd_sc_hd__buf_12
Xoutput178 net178 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
XFILLER_87_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_45.mux_l2_in_0_ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_55_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk sb_1__1_.mem_right_track_20.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_2_ net88 cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_316_ net122 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output293_A net293 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 chanx_right_in_0[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput25 chanx_left_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
Xinput14 chanx_left_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_4
Xinput47 chanx_right_in_0[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
Xinput69 chany_bottom_in[15] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_4
Xinput58 chanx_right_in_0[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_4
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_4__A0 sb_1__1_.mux_left_track_37.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_0__A1 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_1__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_20.mux_l3_in_1_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_2__A0 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_8.ccff_tail
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_1.mux_l3_in_0_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_44.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk sb_1__1_.mem_left_track_7.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_51_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_27_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input52_A chanx_right_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_3_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l2_in_3__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_45.mux_l1_in_1_ net283 net37 sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_45_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__300__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_3_ net102 net71 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_20.mux_l2_in_2_ net11 net85 sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xhold3 cby_1__1_.mem_right_ipin_1.ccff_tail VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_1_ net67 cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_2.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_20.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_21_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__332
+ VGND VGND VPWR VPWR net332 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__332/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_3_2__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input15_A chanx_left_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_21_prog_clk sb_1__1_.mem_left_track_29.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_8_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_60_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__349
+ VGND VGND VPWR VPWR net349 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__349/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__375
+ VGND VGND VPWR VPWR net375 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__375/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input7_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_52.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_53.mux_l1_in_0__A0 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_280_ net26 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_1.mux_l1_in_2_ net108 net77 cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_1_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_4.mux_l2_in_3__405 VGND VGND VPWR VPWR net405 sb_1__1_.mux_right_track_4.mux_l2_in_3__405/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_1__A0 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_0.mux_l2_in_3_ net398 net4 sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_6.mux_l3_in_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_1.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__1_.mux_top_ipin_11.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_67_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_52.mux_l3_in_0_ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_0.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_0__S sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_12.mux_l2_in_3__400 VGND VGND VPWR VPWR net400 sb_1__1_.mux_right_track_12.mux_l2_in_3__400/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_28.mux_l2_in_3__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input117_A chany_top_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_332_ sb_1__1_.mux_bottom_track_11.out VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_0__A1 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_263_ sb_1__1_.mux_left_track_29.out VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input82_A chany_bottom_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_3__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput168 net168 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
XANTENNA__303__A net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput157 net157 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
XFILLER_87_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput179 net179 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
XFILLER_83_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_0__A0 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_12.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_11_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_3.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_74_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_1_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_315_ sb_1__1_.mux_bottom_track_45.out VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_56_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput37 chanx_right_in_0[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_4
XANTENNA_output286_A net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput26 chanx_left_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_4
Xinput15 chanx_left_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
Xinput48 chanx_right_in_0[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__372
+ VGND VGND VPWR VPWR net372 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__372/LO
+ sky130_fd_sc_hd__conb_1
Xinput59 chanx_right_in_0[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_52.mux_l2_in_1_ net418 sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_52.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_20.mux_l3_in_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_33_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_2__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_16_prog_clk sb_1__1_.mem_left_track_7.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_3__319 VGND VGND VPWR VPWR net319 cby_1__1_.mux_right_ipin_15.mux_l2_in_3__319/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_right_track_0.mux_l4_in_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input45_A chanx_right_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_7__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_bottom_track_45.mux_l1_in_0_ net54 net97 sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_1__A0 sb_1__1_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_14_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_88_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_52.mux_l1_in_2_ net5 net23 sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_20.mux_l2_in_1_ net71 sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold4 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_39_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_0_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_62_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_2__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_3_ net421 net58 cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_0.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__311__A sb_1__1_.mux_bottom_track_53.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_3__S sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_3__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_20.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_0.mux_l3_in_1_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_right_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_53_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_2__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net356 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input147_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net370 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk sb_1__1_.mem_left_track_29.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_3__425 VGND VGND VPWR VPWR net425 cbx_1__1_.mux_top_ipin_13.mux_l2_in_3__425/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_94_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_3__313 VGND VGND VPWR VPWR net313 cby_1__1_.mux_right_ipin_1.mux_l2_in_3__313/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l2_in_3__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_right_track_12.mux_l2_in_3__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_10.mux_l2_in_3_ net410 net28 sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_58_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_44.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_53.mux_l1_in_0__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_20.mux_l1_in_2_ net80 net136 sb_1__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_1.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_29.mux_l2_in_3_ net391 net295 sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net341 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_0.mux_l2_in_2_ net21 net87 sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_11.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk sb_1__1_.mem_bottom_track_53.ccff_tail
+ net304 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_3__A1 net299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_331_ sb_1__1_.mux_bottom_track_13.out VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_46_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_262_ net39 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_1.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_input75_A chany_bottom_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_0__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_10.mux_l1_in_4_ net13 net88 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_39_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_3__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput158 net158 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput169 net169 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
XFILLER_68_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_3__392 VGND VGND VPWR VPWR net392 sb_1__1_.mux_left_track_3.mux_l2_in_3__392/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_2_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk cby_1__1_.ccff_tail net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_0.mux_l1_in_3_ net64 net81 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
X_314_ net120 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l2_in_2__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput27 chanx_left_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput16 chanx_left_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_4
Xinput49 chanx_right_in_0[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_6__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput38 chanx_right_in_0[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
XANTENNA_sb_1__1_.mux_top_track_12.mux_l1_in_2__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_10.mux_l4_in_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_52.mux_l2_in_0_ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_3_ net308 net59 cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_2__A0 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_3__324 VGND VGND VPWR VPWR net324 cby_1__1_.mux_right_ipin_6.mux_l2_in_3__324/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_92_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_29.mux_l4_in_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_left_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA__314__A net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net367 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__mux2_4
XFILLER_57_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_1.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_7.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_24_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_2.mux_l2_in_3__412 VGND VGND VPWR VPWR net412 sb_1__1_.mux_top_track_2.mux_l2_in_3__412/LO
+ sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_3_ net386 net29 sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in net138 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_78_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input38_A chanx_right_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_4__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_54_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_54_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__309__A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_1__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_10.mux_l3_in_1_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_52.mux_l1_in_1_ net65 net35 sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_4_ sb_1__1_.mux_left_track_37.out net5 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_12_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_20.mux_l2_in_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_39_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_29.mux_l3_in_1_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_left_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_2__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_3__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_2_ net27 net38 cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_12.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_0.mux_l3_in_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_right_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_4_ net19 net285 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_53_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_6.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_3__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_1__1_.mem_left_track_29.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_1__A1 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_21.mux_l2_in_3__A1 net300 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_7.mux_l4_in_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_10.mux_l2_in_2_ net6 sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_top_track_10.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__322__A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_41_prog_clk
+ sb_1__1_.mem_bottom_track_11.mem_out\[2\] net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_36_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_20.mux_l1_in_1_ net130 net115 sb_1__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_1.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_1_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_29.mux_l2_in_2_ net74 net69 sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_49_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dfrtp_1
XANTENNA_input20_A chanx_left_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_0.mux_l2_in_1_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_6.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__317__A net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_9_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_20.mux_l1_in_2__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_330_ net108 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ net38 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_5__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input68_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_12.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_1_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_7.mux_l3_in_1_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_10.mux_l1_in_3_ net73 net58 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_60_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput159 net159 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l2_in_2__A0 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_86_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input122_A chany_top_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_0.mux_l1_in_2_ net135 net132 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_313_ net119 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput28 chanx_left_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_4
Xinput17 chanx_left_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_4
Xinput39 chanx_right_in_0[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XANTENNA_sb_1__1_.mux_top_track_12.mux_l1_in_2__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_44.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_2_ net28 cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_2__A1 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__361
+ VGND VGND VPWR VPWR net361 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__361/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_1__A0 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__330__A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_1.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_5.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_3__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_2_ net16 sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_bottom_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net345 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_4__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_23_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__325__A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_10.mux_l3_in_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_52.mux_l1_in_0_ net54 net144 sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_3_ net42 net11 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input50_A chanx_right_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_29.mux_l3_in_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_61_prog_clk net430 net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_2__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_1_ net7 cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_26_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_3_ net283 net281 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_7.mux_l2_in_3_ net397 net299 sb_1__1_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_10.mux_l2_in_3__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_21.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input98_A chany_top_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_4__A0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_10.mux_l2_in_1_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_1__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_40_prog_clk
+ sb_1__1_.mem_bottom_track_11.mem_out\[1\] net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_20.mux_l1_in_0_ net101 net105 sb_1__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_4__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_29.mux_l2_in_1_ net70 net44 sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_49_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input13_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_1.mux_l1_in_2_ net48 net17 cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_0.mux_l2_in_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_2.mux_l2_in_3__401 VGND VGND VPWR VPWR net401 sb_1__1_.mux_right_track_2.mux_l2_in_3__401/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net359 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l1_in_4_ net295 net293 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_6.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__333__A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_44.mux_l3_in_0_ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_20.mux_l1_in_2__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ net37 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_12.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_66_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_7.mux_l3_in_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l4_in_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_45_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_10.mux_l1_in_2_ net43 net45 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_48_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_48_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l2_in_2__A1 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_0.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA__328__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk sb_1__1_.mem_bottom_track_1.ccff_tail
+ net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_0__A0 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input115_A chany_top_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_0.mux_l1_in_1_ net129 net93 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_312_ net118 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input80_A chany_bottom_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_left_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_4
Xinput29 chanx_left_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_44.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_44.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_44.mux_l2_in_1_ net406 sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_44.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l2_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_4__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net138 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_68_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_3__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_1_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l3_in_1_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_0__A1 net141 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_2__A0 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net349 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__mux2_4
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_16_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_55_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_12_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_12.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__354
+ VGND VGND VPWR VPWR net354 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__354/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_right_track_44.mux_l1_in_2_ net7 net67 sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input43_A chanx_right_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_2__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_1__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_2_ net287 net59 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l2_in_2_ net297 sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_left_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__336__A sb_1__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_right_track_36.mux_l2_in_1__404 VGND VGND VPWR VPWR net404 sb_1__1_.mux_right_track_36.mux_l2_in_1__404/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_4.mux_l1_in_1__A0 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_3_ net317 net115 cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_52_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_44.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_4__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_10.mux_l2_in_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_41_prog_clk
+ sb_1__1_.mem_bottom_track_11.mem_out\[0\] net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_3__309 VGND VGND VPWR VPWR net309 cbx_1__1_.mux_top_ipin_7.mux_l2_in_3__309/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_left_track_29.mux_l2_in_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_39_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input145_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_1.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_3__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_7.mux_l1_in_3_ net89 net76 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_67_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_3_ net424 net59 cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_58_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_3__A1 net282 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l2_in_3__A1 sb_1__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_12.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_0.mux_l2_in_3__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_10.mux_l1_in_1_ net146 net144 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_82_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_17_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_17_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_13.mux_l4_in_0_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_0.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_2__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_29.mux_l1_in_1_ net39 net104 sb_1__1_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__344__A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_2.mux_l2_in_2__A0 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_1__S sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_0__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input108_A chany_top_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_0.mux_l1_in_0_ net94 net111 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_311_ sb_1__1_.mux_bottom_track_53.out VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput19 chanx_left_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_4
XANTENNA__254__A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_36.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_input73_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_69_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_44.mux_l2_in_0_ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_44.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_80_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_4_ sb_1__1_.mux_left_track_37.out net5 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_2__S sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_2__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__339__A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_4__A0 sb_1__1_.mux_left_track_37.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l3_in_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__249__A net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_2__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_12.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_13.mux_l3_in_1_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_1__S sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_32_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_12.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_6.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_44.mux_l1_in_1_ net84 net133 sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input36_A chanx_right_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l2_in_1__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_1__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_0__A0 sb_1__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_1_ net40 net46 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l2_in_1_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__352__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_4.mux_l1_in_1__A1 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_12.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_2_ net74 net95 cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_44.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_44.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__262__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_2.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.out sky130_fd_sc_hd__buf_4
XFILLER_47_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_42_prog_clk
+ sb_1__1_.mem_bottom_track_11.ccff_head net303 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__347__A net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_4__S sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l2_in_3__A1 net299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input138_A test_enable_bottom_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_1.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_10.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA__257__A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_3__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_3_ net320 sb_1__1_.mux_bottom_track_53.out cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_7.mux_l1_in_2_ net82 net59 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_82_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_45.mux_l2_in_1__383 VGND VGND VPWR VPWR net383 sb_1__1_.mux_bottom_track_45.mux_l2_in_1__383/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_4__A0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_2_ net28 cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_43_prog_clk cby_1__1_.mem_right_ipin_12.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_10.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_66_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_10.mux_l1_in_0_ net142 net148 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_72_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l2_in_1__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_27_prog_clk sb_1__1_.mem_right_track_0.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_57_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_57_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_29.mux_l1_in_0_ net99 net109 sb_1__1_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_7__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__362
+ VGND VGND VPWR VPWR net362 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__362/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__360__A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_2.mux_l2_in_2__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_310_ net116 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_4_ net94 net92 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_42_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input66_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_1__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__270__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_3_ net42 net11 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_2__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__355__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_2.mux_l4_in_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_3__317 VGND VGND VPWR VPWR net317 cby_1__1_.mux_right_ipin_13.mux_l2_in_3__317/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_59_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input120_A chany_top_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__265__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_2_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_13.mux_l3_in_0_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_5.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_1__A0 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_2__A0 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_27_prog_clk sb_1__1_.mem_top_track_12.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_6.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net331 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__mux2_4
Xsb_1__1_.mux_right_track_44.mux_l1_in_0_ net121 net97 sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_3_ net325 sb_1__1_.mux_bottom_track_45.out cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xoutput290 net290 VGND VGND VPWR VPWR test_enable_bottom_out sky130_fd_sc_hd__buf_12
XFILLER_59_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input29_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__343
+ VGND VGND VPWR VPWR net343 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__343/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_0_prog_clk cbx_1__1_.mem_top_ipin_13.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_20.mux_l2_in_3__413 VGND VGND VPWR VPWR net413 sb_1__1_.mux_top_track_20.mux_l2_in_3__413/LO
+ sky130_fd_sc_hd__conb_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew301 net123 VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__buf_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_2.mux_l3_in_1_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_0_ net119 net106 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l2_in_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_1__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_1_ net64 cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_12.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_36.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk cby_1__1_.mem_right_ipin_15.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR cby_1__1_.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_79_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_3__423 VGND VGND VPWR VPWR net423 cbx_1__1_.mux_top_ipin_11.mux_l2_in_3__423/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l2_in_3__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_4.mux_l2_in_3_ net416 net27 sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__363__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_1__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_44_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input96_A chany_top_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__273__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_53.mux_l3_in_0_ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_53.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__357
+ VGND VGND VPWR VPWR net357 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__357/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_2_ net86 cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_25_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_7.mux_l1_in_1_ net46 net119 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_67_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_7.mux_l4_in_0_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_4__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_13.mux_l1_in_2_ net101 net70 cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_86_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__358__A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_2__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_1__A1 net143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input150_A top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_77_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__268__A net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input11_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_25_prog_clk sb_1__1_.mem_right_track_0.ccff_head
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_63_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_8.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_26_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_26_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l2_in_1__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_86_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input3_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_53.mux_l2_in_1_ net385 sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_53.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_3_ sb_1__1_.mux_bottom_track_29.out net69 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_left_track_37.mux_l1_in_2__A0 net296 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_13.mux_l2_in_3_ net389 net299 sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_4.mux_l4_in_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_1__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input59_A chanx_right_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l2_in_3__A1 sb_1__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_7.mux_l3_in_1_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_3__322 VGND VGND VPWR VPWR net322 cby_1__1_.mux_right_ipin_4.mux_l2_in_3__322/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_369_ net301 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_5.mux_l2_in_2__A0 net295 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__371__A net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_2__A0 net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input113_A chany_top_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_53.mux_l1_in_2_ net5 net24 sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_1__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_4.mux_l3_in_1_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_24_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_41_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_2__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_6.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_27_prog_clk sb_1__1_.mem_top_track_10.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xoutput280 net280 VGND VGND VPWR VPWR reset_top_out sky130_fd_sc_hd__buf_12
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_2_ net90 net101 cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xoutput291 net291 VGND VGND VPWR VPWR test_enable_left_out sky130_fd_sc_hd__buf_12
XFILLER_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__276__A sb_1__1_.mux_left_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output282_A net282 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew302 net304 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_16
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_2.mux_l3_in_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_13.mux_l4_in_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_2.mem_out\[2\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net360 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__mux2_4
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_1__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_0_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_56_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_39_prog_clk cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_15.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_15_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input41_A chanx_right_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_85_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_1__S sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_3_ net377 net28 sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_90_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_54_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_4.mux_l2_in_2_ net30 net17 sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l2_in_1__A0 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_2__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__336
+ VGND VGND VPWR VPWR net336 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__336/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_1__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_2__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input89_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_1_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l1_in_0_ net121 net106 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_28.mux_l1_in_0__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_13.mux_l3_in_1_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l2_in_3__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_3__386 VGND VGND VPWR VPWR net386 sb_1__1_.mux_bottom_track_7.mux_l2_in_3__386/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_63_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_13.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in net138 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_left_track_45.mux_l1_in_2__A0 net297 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_2__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__374__A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_4_ net15 net286 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net362 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input143_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__284__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_36.mem_out\[1\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_36_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_86_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__369__A net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_11.mux_l4_in_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_53.mux_l2_in_0_ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_2_ net107 net76 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_54_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_13.mux_l2_in_2_ net293 net86 sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_37.mux_l1_in_2__A1 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l2_in_2__A0 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__279__A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_7.mux_l3_in_0_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_33_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_368_ net123 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_299_ net17 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_left_track_5.mux_l2_in_2__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_2__A1 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l2_in_3__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_5.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input106_A chany_top_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input71_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_4__S sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_11.mux_l3_in_1_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_53.mux_l1_in_1_ net284 net33 sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_88_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_37.mux_l2_in_1__393 VGND VGND VPWR VPWR net393 sb_1__1_.mux_left_track_37.mux_l2_in_1__393/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_4.mux_l3_in_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_64_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__382__A net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_2__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_4.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_10_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_10_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_1_ net70 cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xoutput270 net270 VGND VGND VPWR VPWR chany_top_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput292 net292 VGND VGND VPWR VPWR test_enable_top_out sky130_fd_sc_hd__buf_12
XFILLER_58_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput281 net281 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_10_
+ sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_0__S sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_30_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_90_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__292__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_2__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xload_slew303 net304 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__buf_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l1_in_0__A0 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__377__A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_12.mux_l1_in_0__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_36.mux_l1_in_0__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_4_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_3__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk net431
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_input34_A chanx_right_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_2_ net13 sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_bottom_track_11.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__287__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_0_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_4.mux_l2_in_1_ net90 sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_2__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.out sky130_fd_sc_hd__clkbuf_2
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_7.mux_l1_in_2_ net108 net77 cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_4.mux_l2_in_3__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_10.ccff_head
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_25_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_2__A0 net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_6.mux_l2_in_3_ net408 net29 sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_80_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_4__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_2__A0 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_28.mux_l1_in_0__A1 net141 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_13.mux_l3_in_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_3_ net428 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_48_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_13.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_45.mux_l1_in_2__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_11.ccff_tail
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_3_ net284 net282 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input136_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_3_ net381 net32 sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_8.mem_out\[2\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_82_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_4.mux_l1_in_2_ net77 net60 sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_53_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_2__A0 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk sb_1__1_.mem_right_track_36.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_51_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_6.mux_l1_in_4_ net89 net70 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_35_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_13.mux_l2_in_1_ net72 sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_4_ net34 net32 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_89_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l2_in_2__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_3__S sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__295__A net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
X_367_ sb_1__1_.mux_top_track_0.out VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_298_ net16 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_load_slew304_A net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_6.mux_l4_in_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_right_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_2.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_3__310 VGND VGND VPWR VPWR net310 cbx_1__1_.mux_top_ipin_8.mux_l2_in_3__310/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_74_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_34_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input64_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_4.ccff_tail
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_11.mux_l3_in_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_53.mux_l1_in_0_ net35 net95 sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_3.mux_l4_in_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_83_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_13.mux_l1_in_2_ net79 net56 sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_1__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l1_in_0__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_0__A0 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_50_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_0_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xoutput271 net271 VGND VGND VPWR VPWR chany_top_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput260 net260 VGND VGND VPWR VPWR chany_top_out_0[23] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput293 net293 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_0_ sky130_fd_sc_hd__buf_12
XFILLER_58_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput282 net282 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_11_
+ sky130_fd_sc_hd__buf_12
XFILLER_43_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_3_ net309 sb_1__1_.mux_left_track_45.out cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_12.ccff_tail
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_11_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_2__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_6.mux_l3_in_1_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xload_slew304 net123 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__buf_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_36.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_2.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_69_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l1_in_0__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_0__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_4__A0 net295 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk cby_1__1_.mem_right_ipin_14.ccff_tail
+ net304 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input27_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_1_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l2_in_2__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_3.mux_l3_in_1_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_bottom_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_4.mux_l2_in_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net351 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_left_track_53.mux_l1_in_2__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net342 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__mux2_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l2_in_2__A0 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_7.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_3__307 VGND VGND VPWR VPWR net307 cbx_1__1_.mux_top_ipin_5.mux_l2_in_3__307/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.out sky130_fd_sc_hd__buf_4
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_6.mux_l2_in_2_ net16 sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_right_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_4__A1 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_0__A1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_2__A1 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__298__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net126 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net138 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_2_ net26 cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output300_A net300 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_1 cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_ VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_7.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_2_ net288 net58 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_2_ net18 net22 sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_input129_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_72_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_4.mux_l1_in_1_ net47 net50 sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_383_ net138 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_1
XFILLER_82_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_4__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input94_A chany_top_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_5_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_5_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_2__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_28.ccff_tail
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_63_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_7.ccff_tail
+ net301 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_0_clk0_A clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_1__S cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_6.mux_l1_in_3_ net76 net135 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_6.mux_l2_in_3__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_24_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_13.mux_l2_in_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_50_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_3_ sb_1__1_.mux_left_track_29.out net9 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_18_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_366_ sb_1__1_.mux_top_track_2.out VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_297_ sb_1__1_.mux_right_track_20.out VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mux_top_track_44.mux_l2_in_1__417 VGND VGND VPWR VPWR net417 sb_1__1_.mux_top_track_44.mux_l2_in_1__417/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__1_.mux_top_ipin_7.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_3_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_3_ net286 net283 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_3_ net392 net300 sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_input1_A ccff_head_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l2_in_3__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net340 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_52_prog_clk
+ sb_1__1_.mem_bottom_track_21.mem_out\[2\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__371
+ VGND VGND VPWR VPWR net371 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__371/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input57_A chanx_right_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l2_in_2__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_349_ sb_1__1_.mux_top_track_36.out VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_13.mux_l1_in_1_ net42 net116 sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_68_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_0__A1 net143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput261 net261 VGND VGND VPWR VPWR chany_top_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput250 net250 VGND VGND VPWR VPWR chany_top_out_0[14] sky130_fd_sc_hd__buf_12
XFILLER_79_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput294 net294 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_1_ sky130_fd_sc_hd__buf_12
Xoutput272 net272 VGND VGND VPWR VPWR chany_top_out_0[7] sky130_fd_sc_hd__buf_12
Xoutput283 net283 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_12_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input111_A chany_top_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_2_ net30 net41 cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk
+ sb_1__1_.mem_bottom_track_53.mem_out\[1\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_53.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_right_track_6.mux_l3_in_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_36.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_2.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk cbx_1__1_.mem_top_ipin_1.ccff_tail
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_84_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_3__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_4__A1 net293 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_3.mux_l3_in_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_bottom_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l4_in_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_11_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l2_in_2__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_4__S cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_7.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_29_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_29_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_6.mux_l2_in_1_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_25_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_2 cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l2_in_3__A1 net299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_14_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_1_ net43 net45 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_53_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_1_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l3_in_1_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_left_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_72_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_top_track_28.mux_l2_in_2__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_top_track_4.mux_l1_in_0_ net144 net141 sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_382_ net138 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_1__A0 sb_1__1_.mux_left_track_11.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input87_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_4.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_28.mux_l2_in_3_ net414 net14 sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_95_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput150 top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR net150
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_50_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_6.mux_l1_in_2_ net133 net131 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_44_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_44_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_2_ net47 net16 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input141_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_3__380 VGND VGND VPWR VPWR net380 sb_1__1_.mux_bottom_track_29.mux_l2_in_3__380/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_365_ sb_1__1_.mux_top_track_4.out VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_1
X_296_ net13 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_7.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_3__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_2_ net288 net61 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_2_ net297 net294 sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_59_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_4.ccff_tail
+ net301 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_3__315 VGND VGND VPWR VPWR net315 cby_1__1_.mux_right_ipin_11.mux_l2_in_3__315/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_41_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk
+ sb_1__1_.mem_bottom_track_21.mem_out\[1\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_3.mem_out\[2\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_348_ net65 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l2_in_2__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_279_ net25 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_13.mux_l1_in_0_ net100 net102 sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput262 net262 VGND VGND VPWR VPWR chany_top_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput251 net251 VGND VGND VPWR VPWR chany_top_out_0[15] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_top_track_28.mux_l4_in_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_top_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xoutput240 net240 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
Xoutput295 net295 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_2_ sky130_fd_sc_hd__buf_12
Xoutput273 net273 VGND VGND VPWR VPWR chany_top_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput284 net284 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_13_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_1_ net10 cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input104_A chany_top_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk
+ sb_1__1_.mem_bottom_track_53.mem_out\[0\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_53.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_28.ccff_tail
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_37.mux_l3_in_0_ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_3.mux_l1_in_3_ net92 net78 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_1__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l2_in_2__A0 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_28.mux_l3_in_1_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_top_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_12.mux_l2_in_2__A0 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_7.mux_l1_in_2_ net48 net17 cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_43_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_6.mux_l2_in_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l2_in_3__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_37.mux_l2_in_1_ net393 sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input32_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net303 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_3 sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l3_in_0_ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_0_ net118 net103 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_28.mem_out\[2\]
+ net303 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_3_ net318 sb_1__1_.mux_bottom_track_53.out
+ cby_1__1_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_2__A0 net293 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l3_in_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_left_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_45_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_7.ccff_tail
+ net304 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_28.mux_l2_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_381_ net138 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_82_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_4.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_28.mux_l2_in_2_ net9 net19 sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput140 test_enable_top_in VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_6.mux_l1_in_1_ net129 net119 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net332 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_37.mux_l1_in_2_ net296 net66 sb_1__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_35_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_13_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input134_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.out sky130_fd_sc_hd__buf_4
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_364_ sb_1__1_.mux_top_track_6.out VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_295_ net12 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l2_in_1__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__344
+ VGND VGND VPWR VPWR net344 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__344/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_3__320 VGND VGND VPWR VPWR net320 cby_1__1_.mux_right_ipin_2.mux_l2_in_3__320/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_52.mux_l2_in_1_ net407 sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_52.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_4_ net94 net92 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_3_ net425 net55 cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_44_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_1__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_1_ net62 net48 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_1_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_59_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net358 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_41_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk
+ sb_1__1_.mem_bottom_track_21.mem_out\[0\] net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_3.mem_out\[1\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l2_in_3__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
X_347_ net64 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_278_ net14 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_14.mux_l4_in_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_load_slew302_A net304 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput252 net252 VGND VGND VPWR VPWR chany_top_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput230 net230 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xoutput241 net241 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
Xoutput263 net263 VGND VGND VPWR VPWR chany_top_out_0[26] sky130_fd_sc_hd__buf_12
Xoutput274 net274 VGND VGND VPWR VPWR chany_top_out_0[9] sky130_fd_sc_hd__buf_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput285 net285 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_14_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput296 net296 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_3_ sky130_fd_sc_hd__buf_12
XFILLER_59_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ sb_1__1_.mem_bottom_track_45.ccff_tail net304 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_55_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net329 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l1_in_2_ net5 net63 sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input62_A chanx_right_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net303 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_3.mux_l1_in_2_ net84 net62 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_1__A0 net281 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_2__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_33_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_3__327 VGND VGND VPWR VPWR net327 cby_1__1_.mux_right_ipin_9.mux_l2_in_3__327/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_62_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_14.mux_l3_in_1_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_0__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l2_in_2__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_28.mux_l3_in_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_21.mux_l2_in_2__A0 net294 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_12.mux_l2_in_2__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_7.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_38_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_10.mux_l2_in_3_ net399 net28 sb_1__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_37.mux_l2_in_0_ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_4_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input25_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_3__384 VGND VGND VPWR VPWR net384 sb_1__1_.mux_bottom_track_5.mux_l2_in_3__384/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_4 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net304 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_2__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_9_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net301 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net303 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__339
+ VGND VGND VPWR VPWR net339 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__339/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk sb_1__1_.mem_right_track_28.mem_out\[1\]
+ net304 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_13.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_2_ net86 cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_2__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_380_ net138 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_4.mem_out\[0\]
+ net302 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mux_top_track_28.mux_l2_in_1_ net74 net69 sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xinput141 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND VGND VPWR
+ VPWR net141 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput130 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND VGND VPWR
+ VPWR net130 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net302 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_52.mux_l2_in_1__407 VGND VGND VPWR VPWR net407 sb_1__1_.mux_right_track_52.mux_l2_in_1__407/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net302 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_10.mux_l1_in_4_ net88 net73 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_6.mux_l1_in_0_ net106 net112 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_59_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net301 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

