magic
tech sky130A
magscale 1 2
timestamp 1656243173
<< obsli1 >>
rect 1104 2159 10856 11441
<< obsm1 >>
rect 750 2128 11118 11472
<< metal2 >>
rect 754 0 810 800
rect 2226 0 2282 800
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6642 0 6698 800
rect 8114 0 8170 800
rect 9586 0 9642 800
rect 11058 0 11114 800
<< obsm2 >>
rect 756 856 11112 11461
rect 866 800 2170 856
rect 2338 800 3642 856
rect 3810 800 5114 856
rect 5282 800 6586 856
rect 6754 800 8058 856
rect 8226 800 9530 856
rect 9698 800 11002 856
<< obsm3 >>
rect 2170 2143 9830 11457
<< metal4 >>
rect 2168 2128 2488 11472
rect 3392 2128 3712 11472
rect 4616 2128 4936 11472
rect 5840 2128 6160 11472
rect 7064 2128 7384 11472
rect 8288 2128 8608 11472
rect 9512 2128 9832 11472
<< labels >>
rlabel metal4 s 3392 2128 3712 11472 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 5840 2128 6160 11472 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8288 2128 8608 11472 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2168 2128 2488 11472 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4616 2128 4936 11472 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7064 2128 7384 11472 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 9512 2128 9832 11472 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 754 0 810 800 6 x[0]
port 3 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 x[1]
port 4 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 x[2]
port 5 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 x[3]
port 6 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 x[4]
port 7 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 x[5]
port 8 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 x[6]
port 9 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 x[7]
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 12000 14000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 113718
string GDS_FILE /home/marwan/clear_signoff_final/openlane/tie_array/runs/tie_array/results/signoff/tie_array.magic.gds
string GDS_START 23752
<< end >>

