* NGSPICE file created from sb_1__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

.subckt sb_1__0_ SC_IN_TOP SC_OUT_TOP Test_en_N_out Test_en_S_in VGND VPWR ccff_head
+ ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11]
+ chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16]
+ chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2]
+ chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7]
+ chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11]
+ chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16]
+ chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] chany_top_out[9] clk_3_N_out clk_3_S_in left_bottom_grid_pin_11_
+ left_bottom_grid_pin_13_ left_bottom_grid_pin_15_ left_bottom_grid_pin_17_ left_bottom_grid_pin_1_
+ left_bottom_grid_pin_3_ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_
+ prog_clk_0_N_in prog_clk_3_N_out prog_clk_3_S_in right_bottom_grid_pin_11_ right_bottom_grid_pin_13_
+ right_bottom_grid_pin_15_ right_bottom_grid_pin_17_ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_
+ right_bottom_grid_pin_5_ right_bottom_grid_pin_7_ right_bottom_grid_pin_9_ top_left_grid_pin_42_
+ top_left_grid_pin_43_ top_left_grid_pin_44_ top_left_grid_pin_45_ top_left_grid_pin_46_
+ top_left_grid_pin_47_ top_left_grid_pin_48_ top_left_grid_pin_49_
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 top_left_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_062_ chanx_right_in[4] VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_10.mux_l3_in_0_ mux_top_track_10.mux_l2_in_1_/X mux_top_track_10.mux_l2_in_0_/X
+ mux_top_track_10.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_10.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l1_in_2__A1 left_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_114_ chanx_left_in[7] VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
X_045_ VGND VGND VPWR VPWR _045_/HI _045_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_10.mux_l2_in_1_ _032_/HI chanx_left_in[9] mux_top_track_10.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_10.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_028_ VGND VGND VPWR VPWR _028_/HI _028_/LO sky130_fd_sc_hd__conb_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 right_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_1__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_6.mux_l1_in_2__S mux_top_track_6.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l2_in_2__A0 left_bottom_grid_pin_9_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l2_in_3__A1 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_10.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_10.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_061_ _061_/A VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _061_/A sky130_fd_sc_hd__buf_4
X_113_ chanx_left_in[11] VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_044_ VGND VGND VPWR VPWR _044_/HI _044_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_10.mux_l2_in_0_ chanx_right_in[19] mux_top_track_10.mux_l1_in_0_/X
+ mux_top_track_10.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_10.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_8.mux_l2_in_3_ _030_/HI chanx_left_in[16] mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _069_/A sky130_fd_sc_hd__buf_4
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_3_ _031_/HI chanx_left_in[2] mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_33.mux_l1_in_1__S mux_left_track_33.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_9.mux_l2_in_2__A1 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_10.mux_l2_in_0__A0 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_3__A0 right_bottom_grid_pin_9_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_10.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_060_ chanx_right_in[2] VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_13 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_112_ chanx_left_in[15] VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
X_043_ VGND VGND VPWR VPWR _043_/HI _043_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__056__A SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_8.mux_l2_in_2_ chanx_left_in[6] right_bottom_grid_pin_17_ mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_2_ chanx_left_in[0] chanx_right_in[2] mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 top_left_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_22.mux_l2_in_0_ mux_top_track_22.mux_l1_in_1_/X mux_top_track_22.mux_l1_in_0_/X
+ mux_top_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_22.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_10.mux_l1_in_0_ chanx_right_in[9] top_left_grid_pin_43_ mux_top_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__064__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_3__A1 right_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_2.mux_l1_in_2__S mux_top_track_2.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xprog_clk_0_FTB00 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
Xmux_top_track_22.mux_l1_in_1_ _039_/HI chanx_left_in[17] mux_top_track_22.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_22.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_12 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_8.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_10.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l2_in_2__A0 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_111_ chanx_left_in[19] VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_042_ VGND VGND VPWR VPWR _042_/HI _042_/LO sky130_fd_sc_hd__conb_1
XANTENNA__072__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xprog_clk_3_N_FTB01 prog_clk_3_S_in VGND VGND VPWR VPWR prog_clk_3_N_out sky130_fd_sc_hd__buf_4
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__067__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ chanx_right_in[1] top_left_grid_pin_48_ mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_1_ right_bottom_grid_pin_9_ right_bottom_grid_pin_1_
+ mux_right_track_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_2.mux_l1_in_1__A1 top_left_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_22.sky130_fd_sc_hd__buf_4_0_ mux_top_track_22.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _108_/A sky130_fd_sc_hd__buf_4
XFILLER_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__080__A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0__A0 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_22.mux_l1_in_0_ chanx_right_in[17] top_left_grid_pin_49_ mux_top_track_22.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_22.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA__075__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _105_/A sky130_fd_sc_hd__buf_4
XFILLER_23_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l2_in_2__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_110_ top_left_grid_pin_43_ VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
X_041_ VGND VGND VPWR VPWR _041_/HI _041_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_14.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _097_/A sky130_fd_sc_hd__buf_4
XANTENNA__083__A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l2_in_0_ top_left_grid_pin_46_ mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l2_in_0_ chany_top_in[16] mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 right_bottom_grid_pin_9_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_22.mux_l1_in_0__A0 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_6__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_14.mux_l1_in_0__A1 top_left_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__091__A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0__A0 top_left_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_2.mux_l2_in_0__S mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_040_ VGND VGND VPWR VPWR _040_/HI _040_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_38.sky130_fd_sc_hd__buf_4_0_ mux_top_track_38.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _116_/A sky130_fd_sc_hd__buf_4
XANTENNA__086__A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l1_in_2__A0 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__094__A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A0 right_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_6__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_22.mux_l1_in_0__A1 top_left_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_8.mux_l1_in_0_ chany_top_in[9] chany_top_in[2] mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_44_ top_left_grid_pin_42_ mux_top_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_6.mux_l1_in_0__A1 top_left_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_099_ _099_/A VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _093_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_24.mux_l1_in_1__A0 right_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_4.mux_l1_in_6_ chanx_left_in[14] chanx_left_in[5] mux_right_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_3.mux_l2_in_1__A0 left_bottom_grid_pin_3_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_left_track_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_3_ _048_/HI left_bottom_grid_pin_15_ mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_098_ _098_/A VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.mux_l1_in_1__A0 right_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_Test_en_N_FTB01_A Test_en_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_4.mux_l1_in_1__S mux_top_track_4.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_5_ right_bottom_grid_pin_17_ right_bottom_grid_pin_15_
+ mux_right_track_4.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_5_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _059_/A sky130_fd_sc_hd__buf_4
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l2_in_3__A1 left_bottom_grid_pin_17_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_2_ left_bottom_grid_pin_11_ left_bottom_grid_pin_7_ mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_2__S mux_left_track_5.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_3_ _029_/HI mux_right_track_4.mux_l1_in_6_/X mux_right_track_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_097_ _097_/A VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_32.mux_l1_in_1__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_17.mux_l1_in_1__A0 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_4_ right_bottom_grid_pin_13_ right_bottom_grid_pin_11_
+ mux_right_track_4.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_4_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_5__S mux_left_track_5.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_3.mux_l2_in_1_ left_bottom_grid_pin_3_ chanx_right_in[13] mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_9.mux_l2_in_3__S mux_left_track_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_3__A1 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_3__A0 left_bottom_grid_pin_5_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_track_4.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_096_ chanx_left_in[18] VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_2_ mux_right_track_4.mux_l1_in_5_/X mux_right_track_4.mux_l1_in_4_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_3_ _053_/HI chanx_left_in[17] mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
X_079_ _079_/A VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_17.mux_l1_in_0__S mux_left_track_17.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_20.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_20.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l1_in_1_ _035_/HI chanx_left_in[13] mux_top_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_3_ right_bottom_grid_pin_9_ right_bottom_grid_pin_7_
+ mux_right_track_4.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_32.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l2_in_0_ chanx_right_in[4] mux_left_track_3.mux_l1_in_0_/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_3__A1 left_bottom_grid_pin_3_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_1__A0 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.mux_l2_in_1_ mux_right_track_16.mux_l1_in_3_/X mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__111__A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_095_ chanx_left_in[17] VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 right_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_3__S mux_left_track_17.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_4.mux_l1_in_2__S mux_right_track_4.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_12.sky130_fd_sc_hd__buf_4_0_ mux_top_track_12.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _103_/A sky130_fd_sc_hd__buf_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_16.mux_l1_in_2_ chanx_left_in[8] right_bottom_grid_pin_11_ mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_078_ _078_/A VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_2_ right_bottom_grid_pin_5_ right_bottom_grid_pin_3_
+ mux_right_track_4.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_20.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l1_in_0_ chanx_right_in[13] top_left_grid_pin_46_ mux_top_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l2_in_2__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_6.mux_l1_in_3_ _043_/HI chanx_left_in[6] mux_top_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_6.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA__114__A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_33.mux_l1_in_1__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_4.mux_l1_in_5__S mux_right_track_4.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[6] mux_left_track_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_094_ chanx_left_in[16] VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
Xmux_top_track_6.mux_l3_in_0_ mux_top_track_6.mux_l2_in_1_/X mux_top_track_6.mux_l2_in_0_/X
+ mux_top_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l2_in_3__S mux_right_track_8.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ _077_/A VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l1_in_1_ right_bottom_grid_pin_3_ chany_top_in[17] mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_6.mux_l2_in_1_ mux_top_track_6.mux_l1_in_3_/X mux_top_track_6.mux_l1_in_2_/X
+ mux_top_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_1_ chany_top_in[15] mux_right_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l2_in_2__A1 right_bottom_grid_pin_17_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l1_in_2_ chanx_right_in[11] chanx_right_in[6] mux_top_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_6.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_6__A0 left_bottom_grid_pin_17_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_6_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_6.mux_l1_in_0__S mux_top_track_6.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_093_ _093_/A VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_076_ chanx_right_in[18] VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_6.mux_l2_in_0_ mux_top_track_6.mux_l1_in_1_/X mux_top_track_6.mux_l1_in_0_/X
+ mux_top_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l1_in_0_ chany_top_in[10] chany_top_in[3] mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_0_ chany_top_in[8] chany_top_in[1] mux_right_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_10.mux_l1_in_0__A0 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__buf_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_059_ _059_/A VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
XFILLER_32_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_6.sky130_fd_sc_hd__buf_4_0_ mux_top_track_6.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _100_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_0.mux_l2_in_2__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_6.mux_l1_in_1_ top_left_grid_pin_49_ top_left_grid_pin_47_ mux_top_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_6.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_6.mux_l1_in_3__S mux_top_track_6.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_6__A1 left_bottom_grid_pin_15_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 right_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_092_ chanx_left_in[14] VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
XFILLER_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_075_ chanx_right_in[17] VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _085_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_10.mux_l1_in_0__A1 top_left_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ _058_/A VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 top_left_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_6.mux_l1_in_0_ top_left_grid_pin_45_ top_left_grid_pin_43_ mux_top_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_33.mux_l1_in_2__S mux_left_track_33.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 right_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _057_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_091_ chanx_left_in[13] VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_3__A1 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_2.mux_l1_in_0__S mux_top_track_2.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_074_ chanx_right_in[16] VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__062__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_12.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_12.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_057_ _057_/A VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 top_left_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_109_ _109_/A VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_9.mux_l2_in_3_ _051_/HI left_bottom_grid_pin_17_ mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA__070__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_0.mux_l2_in_3_ _052_/HI chanx_left_in[12] mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_2.mux_l1_in_3__S mux_top_track_2.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l2_in_1__A1 top_left_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_090_ chanx_left_in[12] VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_073_ _073_/A VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_10.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_12.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_056_ SC_IN_TOP VGND VGND VPWR VPWR SC_OUT_TOP sky130_fd_sc_hd__buf_2
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__068__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_5__A0 right_bottom_grid_pin_17_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_108_ _108_/A VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
X_039_ VGND VGND VPWR VPWR _039_/HI _039_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_17.mux_l1_in_3_ _046_/HI left_bottom_grid_pin_11_ mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_18.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l2_in_2_ left_bottom_grid_pin_9_ left_bottom_grid_pin_1_ mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_0.mux_l2_in_2_ chanx_left_in[2] right_bottom_grid_pin_17_ mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_12.mux_l2_in_0_ mux_top_track_12.mux_l1_in_1_/X mux_top_track_12.mux_l1_in_0_/X
+ mux_top_track_12.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_12.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__buf_4
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_12.mux_l1_in_1__A1 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__076__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_12.mux_l1_in_1_ _033_/HI chanx_left_in[10] mux_top_track_12.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_12.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A0 top_left_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_27_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_072_ chanx_right_in[14] VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
XFILLER_18_9 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l2_in_1_ mux_left_track_17.mux_l1_in_3_/X mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_055_ VGND VGND VPWR VPWR _055_/HI _055_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__084__A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_5__A1 right_bottom_grid_pin_15_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_107_ _107_/A VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
X_038_ VGND VGND VPWR VPWR _038_/HI _038_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_17.mux_l1_in_2_ left_bottom_grid_pin_3_ chanx_right_in[17] mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_18.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_27_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_9.mux_l2_in_1_ chanx_right_in[16] chanx_right_in[6] mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__D mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l2_in_1_ right_bottom_grid_pin_13_ right_bottom_grid_pin_9_
+ mux_right_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_20.mux_l1_in_1__A1 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__092__A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_12.mux_l1_in_0_ chanx_right_in[10] top_left_grid_pin_44_ mux_top_track_12.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A1 top_left_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_071_ chanx_right_in[13] VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
XANTENNA__087__A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_2.mux_l2_in_1__S mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_2.mux_l1_in_3_ _037_/HI chanx_left_in[4] mux_top_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_24.mux_l1_in_3_ _055_/HI chanx_left_in[18] mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_3__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclk_3_N_FTB01 clk_3_S_in VGND VGND VPWR VPWR clk_3_N_out sky130_fd_sc_hd__buf_4
Xmux_top_track_24.mux_l1_in_1_ _040_/HI chanx_left_in[18] mux_top_track_24.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_054_ VGND VGND VPWR VPWR _054_/HI _054_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_3.mux_l2_in_0__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_106_ _106_/A VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l1_in_1_ chanx_right_in[8] chany_top_in[17] mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_037_ VGND VGND VPWR VPWR _037_/HI _037_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.mux_l2_in_0_ chany_top_in[18] mux_left_track_9.mux_l1_in_0_/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l2_in_2__A0 left_bottom_grid_pin_13_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__095__A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_5_ right_bottom_grid_pin_1_
+ mux_right_track_0.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_1_ mux_right_track_24.mux_l1_in_3_/X mux_right_track_24.mux_l1_in_2_/X
+ mux_right_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_1_ mux_top_track_2.mux_l1_in_3_/X mux_top_track_2.mux_l1_in_2_/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_070_ chanx_right_in[12] VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_track_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _109_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l1_in_2_ chanx_left_in[9] right_bottom_grid_pin_13_ mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l1_in_2_ chanx_right_in[4] chanx_right_in[3] mux_top_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[18] top_left_grid_pin_42_ mux_top_track_24.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 top_left_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_053_ VGND VGND VPWR VPWR _053_/HI _053_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_18.sky130_fd_sc_hd__buf_4_0_ mux_top_track_18.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _106_/A sky130_fd_sc_hd__buf_4
XFILLER_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_105_ _105_/A VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l1_in_0_ chany_top_in[10] chany_top_in[3] mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_036_ VGND VGND VPWR VPWR _036_/HI _036_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_2__A1 left_bottom_grid_pin_9_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_2__A0 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__buf_4
Xmux_left_track_9.mux_l1_in_0_ chany_top_in[11] chany_top_in[4] mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_0_ chany_top_in[13] chany_top_in[6] mux_right_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _098_/A sky130_fd_sc_hd__buf_4
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_left_track_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 top_left_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_3__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_3__A1 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l1_in_1_ top_left_grid_pin_49_ top_left_grid_pin_47_ mux_top_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_24.mux_l1_in_1_ right_bottom_grid_pin_5_ chany_top_in[18] mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_83 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_052_ VGND VGND VPWR VPWR _052_/HI _052_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_5.mux_l1_in_0__S mux_left_track_5.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l1_in_2__S mux_top_track_4.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_104_ _104_/A VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
X_035_ VGND VGND VPWR VPWR _035_/HI _035_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_6_ left_bottom_grid_pin_17_ left_bottom_grid_pin_15_ mux_left_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_6.mux_l1_in_2__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_5.mux_l1_in_2__A0 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_track_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_5.mux_l1_in_3__S mux_left_track_5.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_9.mux_l2_in_1__S mux_left_track_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_45_ top_left_grid_pin_43_ mux_top_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l1_in_0_ chany_top_in[11] chany_top_in[4] mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l1_in_3__A1 chanx_left_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_051_ VGND VGND VPWR VPWR _051_/HI _051_/LO sky130_fd_sc_hd__conb_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_24.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_left_track_9.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_103_ _103_/A VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_6.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_6.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_034_ VGND VGND VPWR VPWR _034_/HI _034_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_5_ left_bottom_grid_pin_13_ left_bottom_grid_pin_11_ mux_left_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_52 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_6__S mux_left_track_5.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_18.mux_l1_in_1__A1 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_3__A1 chanx_left_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X ccff_head VGND VGND
+ VPWR VPWR mux_top_track_0.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_18_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l2_in_3__A1 left_bottom_grid_pin_15_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l2_in_3_ _050_/HI mux_left_track_5.mux_l1_in_6_/X mux_left_track_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_prog_clk_3_N_FTB01_A prog_clk_3_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_050_ VGND VGND VPWR VPWR _050_/HI _050_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_102_ _102_/A VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_17.mux_l1_in_1__S mux_left_track_17.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_6.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_033_ VGND VGND VPWR VPWR _033_/HI _033_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 right_bottom_grid_pin_13_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_4_ left_bottom_grid_pin_9_ left_bottom_grid_pin_7_ mux_left_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_22.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_22.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_4.mux_l2_in_0__S mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A1 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__112__A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_2_ mux_left_track_5.mux_l1_in_5_/X mux_left_track_5.mux_l1_in_4_/X
+ mux_left_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_4.mux_l1_in_3__S mux_right_track_4.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_101_ _101_/A VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_032_ VGND VGND VPWR VPWR _032_/HI _032_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_1__S mux_right_track_8.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 right_bottom_grid_pin_9_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_6.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l1_in_3_ left_bottom_grid_pin_5_ left_bottom_grid_pin_3_ mux_left_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_5.mux_l1_in_5__A0 left_bottom_grid_pin_13_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_20.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_22.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _065_/A sky130_fd_sc_hd__buf_4
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_38.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__115__A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_6__S mux_right_track_4.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l1_in_3__A1 left_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_100_ _100_/A VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_031_ VGND VGND VPWR VPWR _031_/HI _031_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_3_ _047_/HI left_bottom_grid_pin_13_ mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l1_in_2_ left_bottom_grid_pin_1_ chanx_right_in[14] mux_left_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_5__A1 left_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_18.mux_l2_in_0_ mux_top_track_18.mux_l1_in_1_/X mux_top_track_18.mux_l1_in_0_/X
+ mux_top_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_18.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_20.mux_l2_in_0_ mux_top_track_20.mux_l1_in_1_/X mux_top_track_20.mux_l1_in_0_/X
+ mux_top_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_20.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_25.mux_l1_in_3__A1 left_bottom_grid_pin_13_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_18.mux_l1_in_1_ _036_/HI chanx_left_in[14] mux_top_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_18.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_20.mux_l1_in_1_ _038_/HI chanx_left_in[16] mux_top_track_20.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_20.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_38.mux_l1_in_0__A0 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_2.mux_l2_in_2__A0 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_1__S mux_top_track_6.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l2_in_1_ mux_left_track_25.mux_l1_in_3_/X mux_left_track_25.mux_l1_in_2_/X
+ mux_left_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_030_ VGND VGND VPWR VPWR _030_/HI _030_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_1_ chanx_right_in[5] chany_top_in[19] mux_left_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_25.mux_l1_in_2_ left_bottom_grid_pin_5_ chanx_right_in[18] mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_20.sky130_fd_sc_hd__buf_4_0_ mux_top_track_20.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _107_/A sky130_fd_sc_hd__buf_4
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_3__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_0.mux_l2_in_0__A0 top_left_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_18.mux_l1_in_0_ chanx_right_in[14] top_left_grid_pin_47_ mux_top_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_18.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_14.sky130_fd_sc_hd__buf_4_0_ mux_top_track_14.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _104_/A sky130_fd_sc_hd__buf_4
XFILLER_29_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_20.mux_l1_in_0_ chanx_right_in[16] top_left_grid_pin_48_ mux_top_track_20.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_20.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_38.mux_l1_in_0__A1 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_2__A1 right_bottom_grid_pin_15_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_33.mux_l1_in_0__S mux_left_track_33.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_16.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_0_ chany_top_in[12] chany_top_in[5] mux_left_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l1_in_1_ chanx_right_in[9] chany_top_in[16] mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_089_ _089_/A VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__060__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_12.mux_l1_in_0__A0 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l2_in_1_ _044_/HI chanx_left_in[8] mux_top_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_32.mux_l2_in_1_ _028_/HI mux_right_track_32.mux_l1_in_2_/X mux_right_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__063__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l1_in_2_ chanx_left_in[10] right_bottom_grid_pin_15_ mux_right_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_2.mux_l1_in_1__S mux_top_track_2.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l2_in_3__A1 left_bottom_grid_pin_17_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_4__A0 right_bottom_grid_pin_13_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_25.mux_l1_in_0_ chany_top_in[9] chany_top_in[2] mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_088_ chanx_left_in[10] VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
XFILLER_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_14.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_14.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_20.mux_l1_in_0__A0 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__071__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_12.mux_l1_in_0__A1 top_left_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l2_in_0_ chanx_right_in[15] mux_top_track_8.mux_l1_in_0_/X mux_top_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__066__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 top_left_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _101_/A sky130_fd_sc_hd__buf_4
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_32.mux_l1_in_1_ right_bottom_grid_pin_7_ chany_top_in[19] mux_right_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_2.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_10.mux_l2_in_1__A1 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__074__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_4__A1 right_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_087_ chanx_left_in[9] VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
XFILLER_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_14.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_20.mux_l1_in_0__A1 top_left_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _089_/A sky130_fd_sc_hd__buf_4
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_3_ _045_/HI left_bottom_grid_pin_17_ mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA__082__A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[8] top_left_grid_pin_42_ mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_32.mux_l1_in_0_ chany_top_in[12] chany_top_in[5] mux_right_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l1_in_2__A0 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l1_in_2__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__090__A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_086_ chanx_left_in[8] VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_1.mux_l2_in_1__A0 left_bottom_grid_pin_5_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _058_/A sky130_fd_sc_hd__buf_4
XFILLER_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_069_ _069_/A VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XFILLER_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l2_in_3__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l2_in_2_ left_bottom_grid_pin_13_ left_bottom_grid_pin_9_ mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_8.mux_l2_in_2__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__088__A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l2_in_3_ _054_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_83 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_14.mux_l1_in_1__A1 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_085_ _085_/A VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_068_ chanx_right_in[10] VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
XFILLER_23_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_6.mux_l1_in_1__A0 top_left_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__096__A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ left_bottom_grid_pin_5_ mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_track_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_2__A1 right_bottom_grid_pin_17_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l1_in_2_ left_bottom_grid_pin_1_ chanx_right_in[12] mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_2.mux_l2_in_2_ chanx_left_in[4] right_bottom_grid_pin_15_ mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_14.mux_l2_in_0_ mux_top_track_14.mux_l1_in_1_/X mux_top_track_14.mux_l1_in_0_/X
+ mux_top_track_14.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_14.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_16.mux_l1_in_2__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_22.mux_l1_in_1__A1 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_17.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
X_084_ chanx_left_in[6] VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_14.mux_l1_in_1_ _034_/HI chanx_left_in[12] mux_top_track_14.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_14.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_38.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_38.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_1__A1 top_left_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_067_ chanx_right_in[9] VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_16.mux_l1_in_1__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l1_in_3__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_18.mux_l1_in_0__A0 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_24.mux_l1_in_2__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clk_3_N_FTB01_A clk_3_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l1_in_1_ chanx_right_in[2] chany_top_in[14] mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ right_bottom_grid_pin_11_ right_bottom_grid_pin_7_
+ mux_right_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l2_in_2__A0 left_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_2__A1 right_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_10.sky130_fd_sc_hd__buf_4_0_ mux_top_track_10.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _102_/A sky130_fd_sc_hd__buf_4
XFILLER_27_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_left_track_5.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_083_ chanx_left_in[5] VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
XFILLER_10_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_14.mux_l1_in_0_ chanx_right_in[12] top_left_grid_pin_45_ mux_top_track_14.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_1__S mux_left_track_5.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_38.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_4.mux_l1_in_3__S mux_top_track_4.mux_l1_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_066_ chanx_right_in[8] VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_32.mux_l1_in_2__A0 chanx_left_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_3_ _042_/HI chanx_left_in[5] mux_top_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
X_049_ VGND VGND VPWR VPWR _049_/HI _049_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_18.mux_l1_in_0__A1 top_left_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail VGND VGND VPWR VPWR mux_left_track_33.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_2__A1 right_bottom_grid_pin_13_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_0_ chany_top_in[7] chany_top_in[0] mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 right_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_4__S mux_left_track_5.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_2__A1 left_bottom_grid_pin_7_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l2_in_1_ _049_/HI mux_left_track_33.mux_l1_in_2_/X mux_left_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_track_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_9.mux_l2_in_2__S mux_left_track_9.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_082_ chanx_left_in[4] VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_2.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_18_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l1_in_3_/X mux_top_track_4.mux_l1_in_2_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_3_ chany_top_in[14] mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_2_ left_bottom_grid_pin_15_ left_bottom_grid_pin_7_ mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_065_ _065_/A VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l1_in_2_ chanx_right_in[7] chanx_right_in[5] mux_top_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_32.mux_l1_in_2__A1 right_bottom_grid_pin_15_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_048_ VGND VGND VPWR VPWR _048_/HI _048_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_38.mux_l2_in_0_ _041_/HI mux_top_track_38.mux_l1_in_0_/X mux_top_track_38.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_38.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_17.mux_l1_in_2__A0 left_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_194 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_17.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_081_ _081_/A VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__buf_4
XFILLER_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l1_in_0_ chany_top_in[7] chany_top_in[0] mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_1_ chanx_right_in[10] chany_top_in[15] mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XTest_en_N_FTB01 Test_en_S_in VGND VGND VPWR VPWR Test_en_N_out sky130_fd_sc_hd__buf_4
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l1_in_4__A0 left_bottom_grid_pin_9_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__110__A top_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _099_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_8.mux_l2_in_1__A1 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_064_ chanx_right_in[6] VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_17.mux_l1_in_2__S mux_left_track_17.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_track_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l1_in_1_ top_left_grid_pin_48_ top_left_grid_pin_46_ mux_top_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_116_ _116_/A VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_4.mux_l1_in_1__S mux_right_track_4.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_2__A0 left_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_047_ VGND VGND VPWR VPWR _047_/HI _047_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_4.mux_l2_in_1__S mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2__A1 chanx_right_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_24.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_38.mux_l1_in_0_ chanx_left_in[1] chanx_right_in[0] mux_top_track_38.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_38.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA__113__A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_6_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_080_ chanx_left_in[2] VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_33.mux_l1_in_0_ chany_top_in[8] chany_top_in[1] mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_4.mux_l1_in_4__S mux_right_track_4.mux_l1_in_6_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l1_in_4__A1 left_bottom_grid_pin_7_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_063_ chanx_right_in[5] VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_8.mux_l2_in_2__S mux_right_track_8.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l1_in_2__A0 left_bottom_grid_pin_15_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_44_ top_left_grid_pin_42_ mux_top_track_4.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_25.mux_l1_in_2__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_115_ chanx_left_in[3] VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
X_046_ VGND VGND VPWR VPWR _046_/HI _046_/LO sky130_fd_sc_hd__conb_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_6.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 right_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_029_ VGND VGND VPWR VPWR _029_/HI _029_/LO sky130_fd_sc_hd__conb_1
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_22.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_25_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

