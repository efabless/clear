magic
tech sky130A
magscale 1 2
timestamp 1656943158
<< viali >>
rect 4537 20553 4571 20587
rect 6377 20553 6411 20587
rect 8493 20553 8527 20587
rect 10333 20553 10367 20587
rect 5181 20485 5215 20519
rect 6745 20417 6779 20451
rect 7389 20417 7423 20451
rect 8309 20417 8343 20451
rect 9229 20417 9263 20451
rect 9505 20417 9539 20451
rect 10149 20417 10183 20451
rect 18889 20417 18923 20451
rect 20545 20417 20579 20451
rect 5917 20349 5951 20383
rect 6837 20349 6871 20383
rect 6929 20349 6963 20383
rect 21189 20349 21223 20383
rect 4905 20281 4939 20315
rect 7573 20281 7607 20315
rect 9689 20281 9723 20315
rect 5641 20213 5675 20247
rect 7941 20213 7975 20247
rect 9045 20213 9079 20247
rect 19257 20213 19291 20247
rect 19625 20213 19659 20247
rect 19993 20213 20027 20247
rect 1501 20009 1535 20043
rect 2053 20009 2087 20043
rect 2697 20009 2731 20043
rect 11437 20009 11471 20043
rect 4353 19941 4387 19975
rect 9413 19941 9447 19975
rect 10517 19941 10551 19975
rect 4813 19873 4847 19907
rect 5549 19873 5583 19907
rect 6469 19873 6503 19907
rect 8125 19873 8159 19907
rect 8953 19873 8987 19907
rect 1685 19805 1719 19839
rect 2237 19805 2271 19839
rect 2513 19805 2547 19839
rect 5089 19805 5123 19839
rect 6653 19805 6687 19839
rect 8033 19805 8067 19839
rect 9597 19805 9631 19839
rect 9873 19805 9907 19839
rect 10701 19805 10735 19839
rect 11253 19805 11287 19839
rect 18357 19805 18391 19839
rect 18613 19805 18647 19839
rect 19257 19805 19291 19839
rect 21373 19805 21407 19839
rect 3985 19737 4019 19771
rect 5641 19737 5675 19771
rect 7941 19737 7975 19771
rect 19717 19737 19751 19771
rect 21106 19737 21140 19771
rect 5733 19669 5767 19703
rect 6101 19669 6135 19703
rect 6745 19669 6779 19703
rect 7113 19669 7147 19703
rect 7573 19669 7607 19703
rect 10057 19669 10091 19703
rect 14197 19669 14231 19703
rect 14473 19669 14507 19703
rect 17233 19669 17267 19703
rect 19993 19669 20027 19703
rect 1961 19465 1995 19499
rect 5457 19465 5491 19499
rect 6009 19465 6043 19499
rect 6745 19465 6779 19499
rect 7481 19465 7515 19499
rect 9965 19465 9999 19499
rect 10609 19465 10643 19499
rect 14105 19465 14139 19499
rect 18061 19465 18095 19499
rect 3617 19397 3651 19431
rect 7389 19397 7423 19431
rect 8861 19397 8895 19431
rect 2145 19329 2179 19363
rect 3893 19329 3927 19363
rect 6561 19329 6595 19363
rect 8585 19329 8619 19363
rect 9597 19329 9631 19363
rect 10149 19329 10183 19363
rect 10425 19329 10459 19363
rect 13562 19329 13596 19363
rect 13829 19329 13863 19363
rect 15218 19329 15252 19363
rect 16937 19329 16971 19363
rect 20830 19329 20864 19363
rect 7297 19261 7331 19295
rect 15485 19261 15519 19295
rect 15761 19261 15795 19295
rect 16681 19261 16715 19295
rect 21097 19261 21131 19295
rect 9413 19193 9447 19227
rect 4537 19125 4571 19159
rect 4997 19125 5031 19159
rect 7849 19125 7883 19159
rect 8125 19125 8159 19159
rect 12449 19125 12483 19159
rect 18337 19125 18371 19159
rect 18981 19125 19015 19159
rect 19441 19125 19475 19159
rect 19717 19125 19751 19159
rect 5457 18921 5491 18955
rect 2329 18853 2363 18887
rect 16129 18853 16163 18887
rect 6285 18785 6319 18819
rect 6837 18785 6871 18819
rect 8493 18785 8527 18819
rect 2513 18717 2547 18751
rect 4721 18717 4755 18751
rect 9321 18717 9355 18751
rect 9781 18717 9815 18751
rect 10057 18717 10091 18751
rect 13737 18717 13771 18751
rect 15218 18717 15252 18751
rect 15485 18717 15519 18751
rect 15761 18717 15795 18751
rect 17509 18717 17543 18751
rect 17785 18717 17819 18751
rect 18797 18717 18831 18751
rect 19257 18717 19291 18751
rect 20913 18717 20947 18751
rect 21281 18717 21315 18751
rect 4445 18649 4479 18683
rect 6929 18649 6963 18683
rect 8309 18649 8343 18683
rect 13470 18649 13504 18683
rect 17242 18649 17276 18683
rect 19524 18649 19558 18683
rect 5089 18581 5123 18615
rect 5917 18581 5951 18615
rect 7021 18581 7055 18615
rect 7389 18581 7423 18615
rect 7849 18581 7883 18615
rect 8217 18581 8251 18615
rect 9137 18581 9171 18615
rect 12357 18581 12391 18615
rect 14105 18581 14139 18615
rect 18429 18581 18463 18615
rect 20637 18581 20671 18615
rect 5089 18377 5123 18411
rect 6377 18377 6411 18411
rect 7573 18377 7607 18411
rect 8309 18377 8343 18411
rect 10885 18377 10919 18411
rect 14105 18377 14139 18411
rect 21373 18377 21407 18411
rect 2513 18309 2547 18343
rect 4077 18309 4111 18343
rect 9689 18309 9723 18343
rect 12970 18309 13004 18343
rect 2789 18241 2823 18275
rect 4353 18241 4387 18275
rect 7665 18241 7699 18275
rect 9413 18241 9447 18275
rect 10793 18241 10827 18275
rect 15494 18241 15528 18275
rect 17794 18241 17828 18275
rect 19461 18241 19495 18275
rect 19717 18241 19751 18275
rect 19993 18241 20027 18275
rect 20260 18241 20294 18275
rect 4629 18173 4663 18207
rect 7481 18173 7515 18207
rect 10977 18173 11011 18207
rect 12725 18173 12759 18207
rect 15761 18173 15795 18207
rect 18061 18173 18095 18207
rect 3249 18105 3283 18139
rect 8033 18105 8067 18139
rect 14381 18105 14415 18139
rect 16681 18105 16715 18139
rect 3617 18037 3651 18071
rect 5641 18037 5675 18071
rect 6009 18037 6043 18071
rect 6929 18037 6963 18071
rect 8769 18037 8803 18071
rect 10425 18037 10459 18071
rect 12449 18037 12483 18071
rect 16037 18037 16071 18071
rect 18337 18037 18371 18071
rect 1961 17833 1995 17867
rect 2513 17833 2547 17867
rect 4077 17833 4111 17867
rect 5457 17833 5491 17867
rect 7113 17833 7147 17867
rect 4721 17697 4755 17731
rect 6101 17697 6135 17731
rect 8033 17697 8067 17731
rect 9597 17697 9631 17731
rect 10885 17697 10919 17731
rect 19625 17697 19659 17731
rect 2145 17629 2179 17663
rect 2697 17629 2731 17663
rect 4445 17629 4479 17663
rect 10609 17629 10643 17663
rect 11345 17629 11379 17663
rect 13737 17629 13771 17663
rect 15485 17629 15519 17663
rect 16129 17629 16163 17663
rect 21106 17629 21140 17663
rect 21373 17629 21407 17663
rect 5825 17561 5859 17595
rect 6469 17561 6503 17595
rect 8217 17561 8251 17595
rect 9413 17561 9447 17595
rect 13470 17561 13504 17595
rect 15218 17561 15252 17595
rect 16374 17561 16408 17595
rect 3433 17493 3467 17527
rect 4537 17493 4571 17527
rect 5181 17493 5215 17527
rect 5917 17493 5951 17527
rect 7573 17493 7607 17527
rect 8125 17493 8159 17527
rect 8585 17493 8619 17527
rect 8953 17493 8987 17527
rect 9321 17493 9355 17527
rect 10057 17493 10091 17527
rect 12357 17493 12391 17527
rect 14105 17493 14139 17527
rect 15761 17493 15795 17527
rect 17509 17493 17543 17527
rect 17877 17493 17911 17527
rect 18153 17493 18187 17527
rect 18889 17493 18923 17527
rect 19257 17493 19291 17527
rect 19993 17493 20027 17527
rect 1961 17289 1995 17323
rect 3249 17289 3283 17323
rect 3617 17289 3651 17323
rect 4537 17289 4571 17323
rect 4997 17289 5031 17323
rect 6377 17289 6411 17323
rect 6837 17289 6871 17323
rect 7573 17289 7607 17323
rect 7941 17289 7975 17323
rect 8033 17289 8067 17323
rect 2697 17221 2731 17255
rect 4905 17221 4939 17255
rect 5825 17221 5859 17255
rect 9229 17221 9263 17255
rect 9873 17221 9907 17255
rect 21106 17221 21140 17255
rect 2145 17153 2179 17187
rect 2973 17153 3007 17187
rect 5549 17153 5583 17187
rect 6745 17153 6779 17187
rect 8953 17153 8987 17187
rect 13378 17153 13412 17187
rect 17868 17153 17902 17187
rect 3709 17085 3743 17119
rect 3801 17085 3835 17119
rect 5181 17085 5215 17119
rect 6929 17085 6963 17119
rect 8125 17085 8159 17119
rect 10885 17085 10919 17119
rect 13645 17085 13679 17119
rect 17601 17085 17635 17119
rect 21373 17085 21407 17119
rect 10149 17017 10183 17051
rect 12265 17017 12299 17051
rect 17233 17017 17267 17051
rect 19993 17017 20027 17051
rect 8677 16949 8711 16983
rect 13921 16949 13955 16983
rect 14289 16949 14323 16983
rect 14657 16949 14691 16983
rect 15577 16949 15611 16983
rect 16957 16949 16991 16983
rect 18981 16949 19015 16983
rect 19257 16949 19291 16983
rect 19625 16949 19659 16983
rect 1961 16745 1995 16779
rect 3801 16745 3835 16779
rect 4169 16745 4203 16779
rect 8953 16745 8987 16779
rect 1593 16677 1627 16711
rect 15485 16677 15519 16711
rect 2697 16609 2731 16643
rect 4629 16609 4663 16643
rect 4813 16609 4847 16643
rect 7205 16609 7239 16643
rect 8033 16609 8067 16643
rect 10977 16609 11011 16643
rect 11161 16609 11195 16643
rect 12357 16609 12391 16643
rect 19441 16609 19475 16643
rect 2145 16541 2179 16575
rect 3157 16541 3191 16575
rect 3433 16541 3467 16575
rect 5825 16541 5859 16575
rect 6101 16541 6135 16575
rect 9781 16541 9815 16575
rect 10057 16541 10091 16575
rect 10885 16541 10919 16575
rect 14105 16541 14139 16575
rect 15761 16541 15795 16575
rect 18889 16541 18923 16575
rect 19697 16541 19731 16575
rect 21097 16541 21131 16575
rect 4537 16473 4571 16507
rect 5181 16473 5215 16507
rect 12624 16473 12658 16507
rect 14372 16473 14406 16507
rect 16028 16473 16062 16507
rect 18622 16473 18656 16507
rect 6561 16405 6595 16439
rect 6929 16405 6963 16439
rect 7021 16405 7055 16439
rect 8125 16405 8159 16439
rect 8217 16405 8251 16439
rect 8585 16405 8619 16439
rect 10517 16405 10551 16439
rect 11713 16405 11747 16439
rect 13737 16405 13771 16439
rect 17141 16405 17175 16439
rect 17509 16405 17543 16439
rect 20821 16405 20855 16439
rect 1961 16201 1995 16235
rect 3341 16201 3375 16235
rect 3801 16201 3835 16235
rect 5549 16201 5583 16235
rect 6377 16201 6411 16235
rect 7389 16201 7423 16235
rect 7941 16201 7975 16235
rect 8309 16201 8343 16235
rect 9045 16201 9079 16235
rect 11897 16201 11931 16235
rect 2789 16133 2823 16167
rect 3709 16133 3743 16167
rect 4537 16133 4571 16167
rect 6745 16133 6779 16167
rect 9965 16133 9999 16167
rect 10793 16133 10827 16167
rect 15209 16133 15243 16167
rect 17794 16133 17828 16167
rect 18705 16133 18739 16167
rect 19318 16133 19352 16167
rect 2145 16065 2179 16099
rect 3065 16065 3099 16099
rect 4813 16065 4847 16099
rect 5457 16065 5491 16099
rect 8401 16065 8435 16099
rect 9321 16065 9355 16099
rect 10241 16065 10275 16099
rect 10517 16065 10551 16099
rect 14309 16065 14343 16099
rect 14565 16065 14599 16099
rect 18061 16065 18095 16099
rect 19073 16065 19107 16099
rect 3893 15997 3927 16031
rect 5733 15997 5767 16031
rect 6837 15997 6871 16031
rect 7021 15997 7055 16031
rect 8493 15997 8527 16031
rect 11989 15997 12023 16031
rect 12173 15997 12207 16031
rect 21189 15929 21223 15963
rect 1593 15861 1627 15895
rect 5089 15861 5123 15895
rect 11529 15861 11563 15895
rect 13185 15861 13219 15895
rect 14933 15861 14967 15895
rect 15577 15861 15611 15895
rect 16681 15861 16715 15895
rect 18337 15861 18371 15895
rect 20453 15861 20487 15895
rect 20821 15861 20855 15895
rect 1961 15657 1995 15691
rect 2513 15657 2547 15691
rect 3341 15657 3375 15691
rect 4353 15657 4387 15691
rect 7389 15657 7423 15691
rect 8585 15657 8619 15691
rect 15485 15657 15519 15691
rect 1593 15589 1627 15623
rect 3985 15589 4019 15623
rect 5365 15589 5399 15623
rect 4813 15521 4847 15555
rect 6285 15521 6319 15555
rect 6837 15521 6871 15555
rect 8033 15521 8067 15555
rect 11437 15521 11471 15555
rect 2145 15453 2179 15487
rect 2697 15453 2731 15487
rect 4997 15453 5031 15487
rect 6009 15453 6043 15487
rect 6929 15453 6963 15487
rect 8953 15453 8987 15487
rect 10241 15453 10275 15487
rect 10517 15453 10551 15487
rect 14105 15453 14139 15487
rect 15761 15453 15795 15487
rect 16773 15453 16807 15487
rect 18429 15453 18463 15487
rect 18797 15453 18831 15487
rect 19625 15453 19659 15487
rect 21373 15453 21407 15487
rect 3065 15385 3099 15419
rect 4905 15385 4939 15419
rect 7021 15385 7055 15419
rect 11161 15385 11195 15419
rect 11805 15385 11839 15419
rect 14372 15385 14406 15419
rect 17040 15385 17074 15419
rect 21106 15385 21140 15419
rect 5641 15317 5675 15351
rect 6101 15317 6135 15351
rect 8125 15317 8159 15351
rect 8217 15317 8251 15351
rect 10793 15317 10827 15351
rect 11253 15317 11287 15351
rect 16405 15317 16439 15351
rect 18153 15317 18187 15351
rect 19349 15317 19383 15351
rect 19993 15317 20027 15351
rect 2789 15113 2823 15147
rect 3985 15113 4019 15147
rect 5549 15113 5583 15147
rect 6009 15113 6043 15147
rect 7573 15113 7607 15147
rect 7849 15113 7883 15147
rect 2053 15045 2087 15079
rect 4629 15045 4663 15079
rect 7113 15045 7147 15079
rect 8309 15045 8343 15079
rect 10517 15045 10551 15079
rect 11805 15045 11839 15079
rect 16068 15045 16102 15079
rect 2329 14977 2363 15011
rect 2605 14977 2639 15011
rect 3617 14977 3651 15011
rect 4537 14977 4571 15011
rect 5641 14977 5675 15011
rect 7205 14977 7239 15011
rect 8217 14977 8251 15011
rect 9229 14977 9263 15011
rect 9873 14977 9907 15011
rect 10793 14977 10827 15011
rect 11529 14977 11563 15011
rect 13185 14977 13219 15011
rect 13452 14977 13486 15011
rect 16313 14977 16347 15011
rect 17978 14977 18012 15011
rect 18245 14977 18279 15011
rect 18889 14977 18923 15011
rect 19625 14977 19659 15011
rect 21106 14977 21140 15011
rect 21373 14977 21407 15011
rect 1593 14909 1627 14943
rect 3341 14909 3375 14943
rect 3525 14909 3559 14943
rect 4445 14909 4479 14943
rect 5457 14909 5491 14943
rect 7021 14909 7055 14943
rect 8401 14909 8435 14943
rect 9321 14909 9355 14943
rect 9505 14909 9539 14943
rect 8861 14841 8895 14875
rect 4997 14773 5031 14807
rect 6469 14773 6503 14807
rect 14565 14773 14599 14807
rect 14933 14773 14967 14807
rect 16865 14773 16899 14807
rect 18521 14773 18555 14807
rect 19993 14773 20027 14807
rect 1961 14569 1995 14603
rect 2605 14569 2639 14603
rect 3985 14569 4019 14603
rect 5457 14569 5491 14603
rect 6285 14569 6319 14603
rect 7757 14569 7791 14603
rect 8953 14569 8987 14603
rect 11253 14569 11287 14603
rect 15853 14569 15887 14603
rect 3065 14501 3099 14535
rect 16589 14501 16623 14535
rect 19901 14501 19935 14535
rect 4537 14433 4571 14467
rect 7389 14433 7423 14467
rect 8309 14433 8343 14467
rect 9413 14433 9447 14467
rect 9597 14433 9631 14467
rect 10701 14433 10735 14467
rect 2145 14365 2179 14399
rect 2421 14365 2455 14399
rect 4445 14365 4479 14399
rect 5733 14365 5767 14399
rect 8125 14365 8159 14399
rect 9321 14365 9355 14399
rect 9965 14365 9999 14399
rect 14473 14365 14507 14399
rect 16129 14365 16163 14399
rect 17969 14365 18003 14399
rect 18245 14365 18279 14399
rect 19257 14365 19291 14399
rect 21281 14365 21315 14399
rect 5089 14297 5123 14331
rect 14718 14297 14752 14331
rect 17702 14297 17736 14331
rect 21014 14297 21048 14331
rect 3341 14229 3375 14263
rect 4353 14229 4387 14263
rect 6745 14229 6779 14263
rect 10793 14229 10827 14263
rect 10885 14229 10919 14263
rect 13737 14229 13771 14263
rect 14105 14229 14139 14263
rect 18797 14229 18831 14263
rect 1685 14025 1719 14059
rect 2421 14025 2455 14059
rect 3065 14025 3099 14059
rect 3433 14025 3467 14059
rect 4261 14025 4295 14059
rect 5641 14025 5675 14059
rect 7205 14025 7239 14059
rect 8033 14025 8067 14059
rect 8401 14025 8435 14059
rect 9045 14025 9079 14059
rect 9413 14025 9447 14059
rect 9873 14025 9907 14059
rect 10885 14025 10919 14059
rect 15209 14025 15243 14059
rect 17417 14025 17451 14059
rect 20729 14025 20763 14059
rect 5181 13957 5215 13991
rect 6009 13957 6043 13991
rect 15485 13957 15519 13991
rect 16681 13957 16715 13991
rect 18530 13957 18564 13991
rect 5273 13889 5307 13923
rect 6837 13889 6871 13923
rect 7481 13889 7515 13923
rect 8493 13889 8527 13923
rect 10241 13889 10275 13923
rect 13297 13889 13331 13923
rect 14096 13889 14130 13923
rect 20186 13889 20220 13923
rect 20453 13889 20487 13923
rect 21189 13889 21223 13923
rect 2145 13821 2179 13855
rect 2329 13821 2363 13855
rect 3525 13821 3559 13855
rect 3617 13821 3651 13855
rect 5089 13821 5123 13855
rect 6653 13821 6687 13855
rect 6745 13821 6779 13855
rect 8677 13821 8711 13855
rect 10333 13821 10367 13855
rect 10517 13821 10551 13855
rect 13553 13821 13587 13855
rect 13829 13821 13863 13855
rect 18797 13821 18831 13855
rect 2789 13753 2823 13787
rect 4629 13685 4663 13719
rect 12173 13685 12207 13719
rect 19073 13685 19107 13719
rect 2697 13481 2731 13515
rect 3985 13481 4019 13515
rect 6377 13481 6411 13515
rect 7849 13481 7883 13515
rect 8953 13481 8987 13515
rect 9321 13481 9355 13515
rect 10517 13481 10551 13515
rect 15485 13481 15519 13515
rect 19533 13481 19567 13515
rect 21189 13481 21223 13515
rect 2053 13413 2087 13447
rect 5825 13413 5859 13447
rect 18889 13413 18923 13447
rect 2329 13345 2363 13379
rect 3341 13345 3375 13379
rect 4537 13345 4571 13379
rect 5181 13345 5215 13379
rect 5365 13345 5399 13379
rect 7021 13345 7055 13379
rect 8309 13345 8343 13379
rect 8493 13345 8527 13379
rect 10241 13345 10275 13379
rect 11345 13345 11379 13379
rect 11529 13345 11563 13379
rect 3065 13277 3099 13311
rect 5457 13277 5491 13311
rect 12173 13277 12207 13311
rect 14105 13277 14139 13311
rect 15761 13277 15795 13311
rect 17509 13277 17543 13311
rect 20913 13277 20947 13311
rect 4445 13209 4479 13243
rect 6745 13209 6779 13243
rect 7389 13209 7423 13243
rect 11253 13209 11287 13243
rect 12418 13209 12452 13243
rect 14350 13209 14384 13243
rect 17754 13209 17788 13243
rect 20668 13209 20702 13243
rect 1685 13141 1719 13175
rect 3157 13141 3191 13175
rect 4353 13141 4387 13175
rect 6837 13141 6871 13175
rect 8217 13141 8251 13175
rect 10885 13141 10919 13175
rect 13553 13141 13587 13175
rect 1501 12937 1535 12971
rect 5273 12937 5307 12971
rect 7113 12937 7147 12971
rect 7665 12937 7699 12971
rect 8125 12937 8159 12971
rect 8677 12937 8711 12971
rect 9137 12937 9171 12971
rect 9689 12937 9723 12971
rect 10609 12937 10643 12971
rect 16681 12937 16715 12971
rect 19349 12937 19383 12971
rect 19809 12937 19843 12971
rect 1961 12869 1995 12903
rect 4169 12869 4203 12903
rect 17794 12869 17828 12903
rect 20922 12869 20956 12903
rect 2237 12801 2271 12835
rect 2881 12801 2915 12835
rect 3341 12801 3375 12835
rect 5365 12801 5399 12835
rect 6745 12801 6779 12835
rect 8033 12801 8067 12835
rect 9045 12801 9079 12835
rect 11161 12801 11195 12835
rect 11897 12801 11931 12835
rect 14217 12801 14251 12835
rect 18061 12801 18095 12835
rect 18337 12801 18371 12835
rect 18981 12801 19015 12835
rect 3617 12733 3651 12767
rect 4445 12733 4479 12767
rect 5181 12733 5215 12767
rect 6469 12733 6503 12767
rect 6653 12733 6687 12767
rect 8217 12733 8251 12767
rect 9321 12733 9355 12767
rect 11989 12733 12023 12767
rect 12173 12733 12207 12767
rect 14473 12733 14507 12767
rect 14749 12733 14783 12767
rect 21189 12733 21223 12767
rect 2605 12665 2639 12699
rect 5733 12665 5767 12699
rect 11529 12597 11563 12631
rect 12725 12597 12759 12631
rect 13093 12597 13127 12631
rect 1593 12393 1627 12427
rect 3433 12393 3467 12427
rect 4537 12393 4571 12427
rect 9689 12393 9723 12427
rect 11069 12393 11103 12427
rect 12081 12393 12115 12427
rect 5549 12325 5583 12359
rect 7297 12325 7331 12359
rect 2237 12257 2271 12291
rect 2881 12257 2915 12291
rect 3985 12257 4019 12291
rect 4997 12257 5031 12291
rect 6285 12257 6319 12291
rect 6745 12257 6779 12291
rect 8401 12257 8435 12291
rect 9137 12257 9171 12291
rect 11529 12257 11563 12291
rect 11621 12257 11655 12291
rect 2421 12189 2455 12223
rect 3065 12189 3099 12223
rect 4169 12189 4203 12223
rect 5181 12189 5215 12223
rect 13737 12189 13771 12223
rect 14197 12189 14231 12223
rect 15025 12189 15059 12223
rect 16681 12189 16715 12223
rect 17141 12189 17175 12223
rect 18797 12189 18831 12223
rect 19257 12189 19291 12223
rect 21373 12189 21407 12223
rect 2973 12121 3007 12155
rect 6837 12121 6871 12155
rect 13470 12121 13504 12155
rect 15292 12121 15326 12155
rect 17386 12121 17420 12155
rect 21106 12121 21140 12155
rect 4077 12053 4111 12087
rect 5089 12053 5123 12087
rect 6929 12053 6963 12087
rect 7665 12053 7699 12087
rect 8033 12053 8067 12087
rect 9229 12053 9263 12087
rect 9321 12053 9355 12087
rect 10609 12053 10643 12087
rect 11713 12053 11747 12087
rect 12357 12053 12391 12087
rect 14473 12053 14507 12087
rect 16405 12053 16439 12087
rect 18521 12053 18555 12087
rect 19625 12053 19659 12087
rect 19993 12053 20027 12087
rect 2053 11849 2087 11883
rect 3157 11849 3191 11883
rect 3617 11849 3651 11883
rect 6929 11849 6963 11883
rect 9229 11849 9263 11883
rect 10885 11849 10919 11883
rect 19625 11849 19659 11883
rect 21281 11849 21315 11883
rect 2605 11781 2639 11815
rect 13737 11781 13771 11815
rect 14105 11781 14139 11815
rect 14810 11781 14844 11815
rect 18806 11781 18840 11815
rect 2237 11713 2271 11747
rect 4445 11713 4479 11747
rect 4721 11713 4755 11747
rect 5365 11713 5399 11747
rect 6377 11713 6411 11747
rect 7665 11713 7699 11747
rect 10793 11713 10827 11747
rect 11529 11713 11563 11747
rect 13194 11713 13228 11747
rect 13461 11713 13495 11747
rect 14565 11713 14599 11747
rect 19073 11713 19107 11747
rect 20738 11713 20772 11747
rect 21005 11713 21039 11747
rect 5457 11645 5491 11679
rect 5641 11645 5675 11679
rect 10057 11645 10091 11679
rect 11069 11645 11103 11679
rect 16773 11645 16807 11679
rect 17233 11645 17267 11679
rect 10425 11577 10459 11611
rect 15945 11577 15979 11611
rect 3893 11509 3927 11543
rect 4997 11509 5031 11543
rect 7205 11509 7239 11543
rect 12081 11509 12115 11543
rect 16221 11509 16255 11543
rect 17693 11509 17727 11543
rect 2053 11305 2087 11339
rect 3065 11305 3099 11339
rect 5549 11305 5583 11339
rect 6745 11305 6779 11339
rect 8953 11305 8987 11339
rect 15485 11305 15519 11339
rect 17417 11305 17451 11339
rect 21005 11305 21039 11339
rect 21281 11305 21315 11339
rect 11253 11237 11287 11271
rect 12357 11237 12391 11271
rect 15761 11237 15795 11271
rect 3985 11169 4019 11203
rect 4997 11169 5031 11203
rect 6193 11169 6227 11203
rect 6285 11169 6319 11203
rect 7757 11169 7791 11203
rect 9505 11169 9539 11203
rect 10701 11169 10735 11203
rect 10885 11169 10919 11203
rect 13737 11169 13771 11203
rect 14105 11169 14139 11203
rect 19625 11169 19659 11203
rect 2237 11101 2271 11135
rect 4261 11101 4295 11135
rect 5089 11101 5123 11135
rect 5181 11101 5215 11135
rect 7481 11101 7515 11135
rect 10609 11101 10643 11135
rect 13470 11101 13504 11135
rect 14372 11101 14406 11135
rect 17141 11101 17175 11135
rect 18797 11101 18831 11135
rect 19881 11101 19915 11135
rect 3433 11033 3467 11067
rect 7205 11033 7239 11067
rect 8585 11033 8619 11067
rect 9321 11033 9355 11067
rect 16896 11033 16930 11067
rect 18552 11033 18586 11067
rect 19257 11033 19291 11067
rect 6377 10965 6411 10999
rect 9413 10965 9447 10999
rect 10241 10965 10275 10999
rect 2053 10761 2087 10795
rect 3985 10761 4019 10795
rect 4629 10761 4663 10795
rect 6745 10761 6779 10795
rect 7113 10761 7147 10795
rect 7757 10761 7791 10795
rect 7849 10761 7883 10795
rect 10333 10761 10367 10795
rect 13001 10761 13035 10795
rect 19717 10761 19751 10795
rect 19993 10761 20027 10795
rect 2605 10693 2639 10727
rect 5733 10693 5767 10727
rect 6653 10693 6687 10727
rect 8677 10693 8711 10727
rect 15770 10693 15804 10727
rect 18582 10693 18616 10727
rect 1869 10625 1903 10659
rect 2881 10625 2915 10659
rect 3617 10625 3651 10659
rect 4261 10625 4295 10659
rect 5273 10625 5307 10659
rect 6009 10625 6043 10659
rect 10241 10625 10275 10659
rect 10885 10625 10919 10659
rect 12633 10625 12667 10659
rect 14114 10625 14148 10659
rect 14381 10625 14415 10659
rect 16681 10625 16715 10659
rect 16948 10625 16982 10659
rect 18337 10625 18371 10659
rect 21106 10625 21140 10659
rect 21373 10625 21407 10659
rect 3341 10557 3375 10591
rect 6561 10557 6595 10591
rect 8033 10557 8067 10591
rect 9137 10557 9171 10591
rect 10517 10557 10551 10591
rect 16037 10557 16071 10591
rect 9873 10489 9907 10523
rect 14657 10489 14691 10523
rect 1501 10421 1535 10455
rect 7389 10421 7423 10455
rect 9413 10421 9447 10455
rect 18061 10421 18095 10455
rect 2053 10217 2087 10251
rect 4169 10217 4203 10251
rect 5549 10217 5583 10251
rect 6837 10217 6871 10251
rect 7849 10217 7883 10251
rect 9689 10217 9723 10251
rect 12357 10217 12391 10251
rect 15761 10217 15795 10251
rect 18797 10217 18831 10251
rect 19441 10217 19475 10251
rect 14105 10149 14139 10183
rect 3893 10081 3927 10115
rect 4813 10081 4847 10115
rect 7481 10081 7515 10115
rect 8493 10081 8527 10115
rect 9137 10081 9171 10115
rect 2237 10013 2271 10047
rect 9321 10013 9355 10047
rect 13470 10013 13504 10047
rect 13737 10013 13771 10047
rect 15485 10013 15519 10047
rect 17141 10013 17175 10047
rect 17417 10013 17451 10047
rect 19993 10013 20027 10047
rect 4537 9945 4571 9979
rect 6561 9945 6595 9979
rect 8217 9945 8251 9979
rect 9229 9945 9263 9979
rect 10701 9945 10735 9979
rect 15218 9945 15252 9979
rect 16874 9945 16908 9979
rect 17684 9945 17718 9979
rect 20238 9945 20272 9979
rect 4629 9877 4663 9911
rect 5825 9877 5859 9911
rect 7205 9877 7239 9911
rect 7297 9877 7331 9911
rect 8309 9877 8343 9911
rect 10241 9877 10275 9911
rect 21373 9877 21407 9911
rect 6745 9673 6779 9707
rect 7849 9673 7883 9707
rect 9413 9673 9447 9707
rect 9781 9673 9815 9707
rect 10425 9673 10459 9707
rect 10793 9673 10827 9707
rect 13921 9673 13955 9707
rect 16681 9673 16715 9707
rect 17141 9673 17175 9707
rect 17509 9673 17543 9707
rect 18245 9673 18279 9707
rect 18889 9673 18923 9707
rect 19809 9673 19843 9707
rect 20269 9673 20303 9707
rect 20913 9673 20947 9707
rect 21281 9673 21315 9707
rect 5733 9605 5767 9639
rect 7113 9605 7147 9639
rect 9873 9605 9907 9639
rect 13286 9605 13320 9639
rect 18521 9605 18555 9639
rect 19533 9605 19567 9639
rect 20545 9605 20579 9639
rect 2237 9537 2271 9571
rect 2513 9537 2547 9571
rect 3065 9537 3099 9571
rect 4537 9537 4571 9571
rect 6009 9537 6043 9571
rect 8769 9537 8803 9571
rect 11529 9537 11563 9571
rect 13553 9537 13587 9571
rect 14473 9537 14507 9571
rect 14729 9537 14763 9571
rect 4721 9469 4755 9503
rect 6377 9469 6411 9503
rect 7205 9469 7239 9503
rect 7297 9469 7331 9503
rect 8861 9469 8895 9503
rect 9045 9469 9079 9503
rect 10057 9469 10091 9503
rect 10885 9469 10919 9503
rect 10977 9469 11011 9503
rect 2053 9401 2087 9435
rect 8401 9401 8435 9435
rect 12173 9401 12207 9435
rect 15853 9401 15887 9435
rect 2697 9333 2731 9367
rect 16129 9333 16163 9367
rect 2145 9129 2179 9163
rect 4537 9129 4571 9163
rect 8033 9129 8067 9163
rect 9597 9129 9631 9163
rect 10609 9129 10643 9163
rect 19809 9129 19843 9163
rect 4261 8993 4295 9027
rect 5181 8993 5215 9027
rect 6193 8993 6227 9027
rect 10241 8993 10275 9027
rect 11253 8993 11287 9027
rect 12265 8993 12299 9027
rect 2329 8925 2363 8959
rect 4997 8925 5031 8959
rect 10057 8925 10091 8959
rect 11989 8925 12023 8959
rect 12633 8925 12667 8959
rect 4905 8857 4939 8891
rect 5917 8857 5951 8891
rect 6561 8857 6595 8891
rect 7665 8857 7699 8891
rect 9321 8857 9355 8891
rect 9965 8857 9999 8891
rect 10977 8857 11011 8891
rect 20361 8857 20395 8891
rect 20729 8857 20763 8891
rect 21097 8857 21131 8891
rect 5549 8789 5583 8823
rect 6009 8789 6043 8823
rect 7113 8789 7147 8823
rect 8585 8789 8619 8823
rect 11069 8789 11103 8823
rect 11621 8789 11655 8823
rect 12081 8789 12115 8823
rect 13737 8789 13771 8823
rect 16037 8789 16071 8823
rect 19257 8789 19291 8823
rect 5181 8585 5215 8619
rect 6837 8585 6871 8619
rect 7389 8585 7423 8619
rect 9045 8585 9079 8619
rect 9413 8585 9447 8619
rect 10425 8585 10459 8619
rect 10885 8585 10919 8619
rect 11713 8585 11747 8619
rect 12449 8585 12483 8619
rect 21005 8585 21039 8619
rect 21281 8585 21315 8619
rect 5641 8517 5675 8551
rect 7757 8517 7791 8551
rect 12173 8517 12207 8551
rect 12909 8517 12943 8551
rect 6745 8449 6779 8483
rect 7849 8449 7883 8483
rect 10793 8449 10827 8483
rect 12817 8449 12851 8483
rect 4905 8381 4939 8415
rect 7021 8381 7055 8415
rect 8033 8381 8067 8415
rect 9505 8381 9539 8415
rect 9689 8381 9723 8415
rect 10977 8381 11011 8415
rect 13093 8381 13127 8415
rect 6009 8313 6043 8347
rect 6377 8245 6411 8279
rect 8677 8245 8711 8279
rect 10057 8245 10091 8279
rect 6009 8041 6043 8075
rect 8953 8041 8987 8075
rect 10609 8041 10643 8075
rect 12265 8041 12299 8075
rect 13277 8041 13311 8075
rect 7297 7973 7331 8007
rect 11253 7973 11287 8007
rect 11897 7973 11931 8007
rect 6469 7905 6503 7939
rect 6653 7905 6687 7939
rect 7757 7905 7791 7939
rect 7941 7905 7975 7939
rect 9597 7905 9631 7939
rect 12725 7905 12759 7939
rect 12817 7905 12851 7939
rect 7665 7837 7699 7871
rect 10241 7837 10275 7871
rect 8585 7769 8619 7803
rect 9321 7769 9355 7803
rect 12633 7769 12667 7803
rect 5641 7701 5675 7735
rect 6377 7701 6411 7735
rect 9413 7701 9447 7735
rect 6009 7497 6043 7531
rect 7021 7497 7055 7531
rect 8125 7497 8159 7531
rect 8401 7497 8435 7531
rect 9505 7497 9539 7531
rect 9873 7497 9907 7531
rect 6745 7429 6779 7463
rect 8861 7429 8895 7463
rect 7389 7361 7423 7395
rect 8769 7361 8803 7395
rect 7481 7293 7515 7327
rect 7573 7293 7607 7327
rect 9045 7293 9079 7327
rect 5641 7157 5675 7191
rect 10241 7157 10275 7191
rect 4721 6953 4755 6987
rect 9045 6953 9079 6987
rect 10333 6953 10367 6987
rect 5273 6885 5307 6919
rect 7573 6817 7607 6851
rect 8309 6817 8343 6851
rect 9689 6817 9723 6851
rect 10977 6817 11011 6851
rect 11805 6817 11839 6851
rect 5089 6749 5123 6783
rect 5641 6749 5675 6783
rect 6193 6749 6227 6783
rect 5825 6613 5859 6647
rect 6377 6613 6411 6647
rect 7021 6613 7055 6647
rect 7389 6613 7423 6647
rect 7481 6613 7515 6647
rect 9413 6613 9447 6647
rect 9505 6613 9539 6647
rect 10701 6613 10735 6647
rect 10793 6613 10827 6647
rect 11437 6613 11471 6647
rect 5549 6409 5583 6443
rect 8125 6409 8159 6443
rect 9137 6409 9171 6443
rect 10149 6409 10183 6443
rect 10609 6409 10643 6443
rect 7757 6273 7791 6307
rect 9505 6273 9539 6307
rect 5917 6205 5951 6239
rect 6929 6205 6963 6239
rect 9597 6205 9631 6239
rect 9781 6205 9815 6239
rect 6469 6069 6503 6103
rect 7205 6069 7239 6103
rect 8769 6069 8803 6103
rect 8953 5865 8987 5899
rect 9321 5865 9355 5899
rect 8493 5797 8527 5831
rect 10885 5185 10919 5219
rect 11529 5185 11563 5219
rect 11069 5049 11103 5083
<< metal1 >>
rect 21174 20748 21180 20800
rect 21232 20788 21238 20800
rect 21818 20788 21824 20800
rect 21232 20760 21824 20788
rect 21232 20748 21238 20760
rect 21818 20748 21824 20760
rect 21876 20748 21882 20800
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 4525 20587 4583 20593
rect 4525 20553 4537 20587
rect 4571 20584 4583 20587
rect 5258 20584 5264 20596
rect 4571 20556 5264 20584
rect 4571 20553 4583 20556
rect 4525 20547 4583 20553
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 5350 20544 5356 20596
rect 5408 20584 5414 20596
rect 6365 20587 6423 20593
rect 6365 20584 6377 20587
rect 5408 20556 6377 20584
rect 5408 20544 5414 20556
rect 6365 20553 6377 20556
rect 6411 20553 6423 20587
rect 6365 20547 6423 20553
rect 8481 20587 8539 20593
rect 8481 20553 8493 20587
rect 8527 20553 8539 20587
rect 8481 20547 8539 20553
rect 10321 20587 10379 20593
rect 10321 20553 10333 20587
rect 10367 20584 10379 20587
rect 12526 20584 12532 20596
rect 10367 20556 12532 20584
rect 10367 20553 10379 20556
rect 10321 20547 10379 20553
rect 5169 20519 5227 20525
rect 5169 20485 5181 20519
rect 5215 20516 5227 20519
rect 8496 20516 8524 20547
rect 12526 20544 12532 20556
rect 12584 20544 12590 20596
rect 13078 20516 13084 20528
rect 5215 20488 6914 20516
rect 8496 20488 13084 20516
rect 5215 20485 5227 20488
rect 5169 20479 5227 20485
rect 5994 20408 6000 20460
rect 6052 20448 6058 20460
rect 6733 20451 6791 20457
rect 6733 20448 6745 20451
rect 6052 20420 6745 20448
rect 6052 20408 6058 20420
rect 6733 20417 6745 20420
rect 6779 20417 6791 20451
rect 6886 20448 6914 20488
rect 13078 20476 13084 20488
rect 13136 20476 13142 20528
rect 6886 20420 6960 20448
rect 6733 20411 6791 20417
rect 5534 20340 5540 20392
rect 5592 20380 5598 20392
rect 5905 20383 5963 20389
rect 5905 20380 5917 20383
rect 5592 20352 5917 20380
rect 5592 20340 5598 20352
rect 5905 20349 5917 20352
rect 5951 20349 5963 20383
rect 5905 20343 5963 20349
rect 4893 20315 4951 20321
rect 4893 20281 4905 20315
rect 4939 20312 4951 20315
rect 5810 20312 5816 20324
rect 4939 20284 5816 20312
rect 4939 20281 4951 20284
rect 4893 20275 4951 20281
rect 5810 20272 5816 20284
rect 5868 20272 5874 20324
rect 5920 20312 5948 20343
rect 6178 20340 6184 20392
rect 6236 20380 6242 20392
rect 6932 20389 6960 20420
rect 7006 20408 7012 20460
rect 7064 20448 7070 20460
rect 7377 20451 7435 20457
rect 7377 20448 7389 20451
rect 7064 20420 7389 20448
rect 7064 20408 7070 20420
rect 7377 20417 7389 20420
rect 7423 20417 7435 20451
rect 8294 20448 8300 20460
rect 8255 20420 8300 20448
rect 7377 20411 7435 20417
rect 8294 20408 8300 20420
rect 8352 20408 8358 20460
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20417 9275 20451
rect 9490 20448 9496 20460
rect 9451 20420 9496 20448
rect 9217 20411 9275 20417
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6236 20352 6837 20380
rect 6236 20340 6242 20352
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 6917 20383 6975 20389
rect 6917 20349 6929 20383
rect 6963 20349 6975 20383
rect 9232 20380 9260 20411
rect 9490 20408 9496 20420
rect 9548 20408 9554 20460
rect 10134 20448 10140 20460
rect 10095 20420 10140 20448
rect 10134 20408 10140 20420
rect 10192 20408 10198 20460
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20448 18935 20451
rect 20533 20451 20591 20457
rect 20533 20448 20545 20451
rect 18923 20420 20545 20448
rect 18923 20417 18935 20420
rect 18877 20411 18935 20417
rect 20533 20417 20545 20420
rect 20579 20448 20591 20451
rect 22278 20448 22284 20460
rect 20579 20420 22284 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 22278 20408 22284 20420
rect 22336 20408 22342 20460
rect 10042 20380 10048 20392
rect 9232 20352 10048 20380
rect 6917 20343 6975 20349
rect 6730 20312 6736 20324
rect 5920 20284 6736 20312
rect 6730 20272 6736 20284
rect 6788 20272 6794 20324
rect 6932 20312 6960 20343
rect 10042 20340 10048 20352
rect 10100 20340 10106 20392
rect 21177 20383 21235 20389
rect 21177 20349 21189 20383
rect 21223 20380 21235 20383
rect 21358 20380 21364 20392
rect 21223 20352 21364 20380
rect 21223 20349 21235 20352
rect 21177 20343 21235 20349
rect 21358 20340 21364 20352
rect 21416 20340 21422 20392
rect 6840 20284 6960 20312
rect 7561 20315 7619 20321
rect 6840 20256 6868 20284
rect 7561 20281 7573 20315
rect 7607 20312 7619 20315
rect 9677 20315 9735 20321
rect 7607 20284 9628 20312
rect 7607 20281 7619 20284
rect 7561 20275 7619 20281
rect 5626 20244 5632 20256
rect 5587 20216 5632 20244
rect 5626 20204 5632 20216
rect 5684 20204 5690 20256
rect 6822 20204 6828 20256
rect 6880 20204 6886 20256
rect 7926 20244 7932 20256
rect 7887 20216 7932 20244
rect 7926 20204 7932 20216
rect 7984 20204 7990 20256
rect 9033 20247 9091 20253
rect 9033 20213 9045 20247
rect 9079 20244 9091 20247
rect 9306 20244 9312 20256
rect 9079 20216 9312 20244
rect 9079 20213 9091 20216
rect 9033 20207 9091 20213
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 9600 20244 9628 20284
rect 9677 20281 9689 20315
rect 9723 20312 9735 20315
rect 14918 20312 14924 20324
rect 9723 20284 14924 20312
rect 9723 20281 9735 20284
rect 9677 20275 9735 20281
rect 14918 20272 14924 20284
rect 14976 20272 14982 20324
rect 13538 20244 13544 20256
rect 9600 20216 13544 20244
rect 13538 20204 13544 20216
rect 13596 20204 13602 20256
rect 19058 20204 19064 20256
rect 19116 20244 19122 20256
rect 19245 20247 19303 20253
rect 19245 20244 19257 20247
rect 19116 20216 19257 20244
rect 19116 20204 19122 20216
rect 19245 20213 19257 20216
rect 19291 20244 19303 20247
rect 19613 20247 19671 20253
rect 19613 20244 19625 20247
rect 19291 20216 19625 20244
rect 19291 20213 19303 20216
rect 19245 20207 19303 20213
rect 19613 20213 19625 20216
rect 19659 20244 19671 20247
rect 19981 20247 20039 20253
rect 19981 20244 19993 20247
rect 19659 20216 19993 20244
rect 19659 20213 19671 20216
rect 19613 20207 19671 20213
rect 19981 20213 19993 20216
rect 20027 20213 20039 20247
rect 19981 20207 20039 20213
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 1486 20040 1492 20052
rect 1447 20012 1492 20040
rect 1486 20000 1492 20012
rect 1544 20000 1550 20052
rect 2038 20040 2044 20052
rect 1999 20012 2044 20040
rect 2038 20000 2044 20012
rect 2096 20000 2102 20052
rect 2685 20043 2743 20049
rect 2685 20009 2697 20043
rect 2731 20040 2743 20043
rect 2774 20040 2780 20052
rect 2731 20012 2780 20040
rect 2731 20009 2743 20012
rect 2685 20003 2743 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 5166 20000 5172 20052
rect 5224 20040 5230 20052
rect 11425 20043 11483 20049
rect 5224 20012 6408 20040
rect 5224 20000 5230 20012
rect 1394 19932 1400 19984
rect 1452 19972 1458 19984
rect 2498 19972 2504 19984
rect 1452 19944 2504 19972
rect 1452 19932 1458 19944
rect 2498 19932 2504 19944
rect 2556 19932 2562 19984
rect 4154 19932 4160 19984
rect 4212 19972 4218 19984
rect 4341 19975 4399 19981
rect 4341 19972 4353 19975
rect 4212 19944 4353 19972
rect 4212 19932 4218 19944
rect 4341 19941 4353 19944
rect 4387 19972 4399 19975
rect 4387 19944 5948 19972
rect 4387 19941 4399 19944
rect 4341 19935 4399 19941
rect 4801 19907 4859 19913
rect 4801 19904 4813 19907
rect 2240 19876 4813 19904
rect 1670 19836 1676 19848
rect 1631 19808 1676 19836
rect 1670 19796 1676 19808
rect 1728 19796 1734 19848
rect 2240 19845 2268 19876
rect 4801 19873 4813 19876
rect 4847 19873 4859 19907
rect 4801 19867 4859 19873
rect 5537 19907 5595 19913
rect 5537 19873 5549 19907
rect 5583 19873 5595 19907
rect 5537 19867 5595 19873
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19805 2283 19839
rect 2498 19836 2504 19848
rect 2459 19808 2504 19836
rect 2225 19799 2283 19805
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 5077 19839 5135 19845
rect 5077 19805 5089 19839
rect 5123 19836 5135 19839
rect 5350 19836 5356 19848
rect 5123 19808 5356 19836
rect 5123 19805 5135 19808
rect 5077 19799 5135 19805
rect 5350 19796 5356 19808
rect 5408 19796 5414 19848
rect 5552 19836 5580 19867
rect 5810 19836 5816 19848
rect 5552 19808 5816 19836
rect 5810 19796 5816 19808
rect 5868 19796 5874 19848
rect 5920 19836 5948 19944
rect 6380 19904 6408 20012
rect 11425 20009 11437 20043
rect 11471 20040 11483 20043
rect 18966 20040 18972 20052
rect 11471 20012 18972 20040
rect 11471 20009 11483 20012
rect 11425 20003 11483 20009
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 9398 19972 9404 19984
rect 9359 19944 9404 19972
rect 9398 19932 9404 19944
rect 9456 19932 9462 19984
rect 9858 19932 9864 19984
rect 9916 19972 9922 19984
rect 10410 19972 10416 19984
rect 9916 19944 10416 19972
rect 9916 19932 9922 19944
rect 10410 19932 10416 19944
rect 10468 19932 10474 19984
rect 10505 19975 10563 19981
rect 10505 19941 10517 19975
rect 10551 19972 10563 19975
rect 15838 19972 15844 19984
rect 10551 19944 15844 19972
rect 10551 19941 10563 19944
rect 10505 19935 10563 19941
rect 15838 19932 15844 19944
rect 15896 19932 15902 19984
rect 6457 19907 6515 19913
rect 6457 19904 6469 19907
rect 6380 19876 6469 19904
rect 6457 19873 6469 19876
rect 6503 19904 6515 19907
rect 8113 19907 8171 19913
rect 8113 19904 8125 19907
rect 6503 19876 8125 19904
rect 6503 19873 6515 19876
rect 6457 19867 6515 19873
rect 8113 19873 8125 19876
rect 8159 19904 8171 19907
rect 8941 19907 8999 19913
rect 8941 19904 8953 19907
rect 8159 19876 8953 19904
rect 8159 19873 8171 19876
rect 8113 19867 8171 19873
rect 8941 19873 8953 19876
rect 8987 19904 8999 19907
rect 11974 19904 11980 19916
rect 8987 19876 9444 19904
rect 8987 19873 8999 19876
rect 8941 19867 8999 19873
rect 9416 19848 9444 19876
rect 9600 19876 11980 19904
rect 6641 19839 6699 19845
rect 6641 19836 6653 19839
rect 5920 19808 6653 19836
rect 6641 19805 6653 19808
rect 6687 19805 6699 19839
rect 6641 19799 6699 19805
rect 6730 19796 6736 19848
rect 6788 19836 6794 19848
rect 8021 19839 8079 19845
rect 8021 19836 8033 19839
rect 6788 19808 8033 19836
rect 6788 19796 6794 19808
rect 8021 19805 8033 19808
rect 8067 19805 8079 19839
rect 8021 19799 8079 19805
rect 9398 19796 9404 19848
rect 9456 19796 9462 19848
rect 9600 19845 9628 19876
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 12710 19864 12716 19916
rect 12768 19904 12774 19916
rect 16298 19904 16304 19916
rect 12768 19876 16304 19904
rect 12768 19864 12774 19876
rect 16298 19864 16304 19876
rect 16356 19864 16362 19916
rect 18524 19876 19748 19904
rect 18524 19848 18552 19876
rect 9585 19839 9643 19845
rect 9585 19805 9597 19839
rect 9631 19805 9643 19839
rect 9858 19836 9864 19848
rect 9819 19808 9864 19836
rect 9585 19799 9643 19805
rect 9858 19796 9864 19808
rect 9916 19796 9922 19848
rect 10686 19836 10692 19848
rect 10647 19808 10692 19836
rect 10686 19796 10692 19808
rect 10744 19796 10750 19848
rect 11238 19836 11244 19848
rect 11199 19808 11244 19836
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 12802 19796 12808 19848
rect 12860 19836 12866 19848
rect 15286 19836 15292 19848
rect 12860 19808 15292 19836
rect 12860 19796 12866 19808
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 18345 19839 18403 19845
rect 18345 19805 18357 19839
rect 18391 19836 18403 19839
rect 18506 19836 18512 19848
rect 18391 19808 18512 19836
rect 18391 19805 18403 19808
rect 18345 19799 18403 19805
rect 18506 19796 18512 19808
rect 18564 19796 18570 19848
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 19058 19836 19064 19848
rect 18647 19808 19064 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 3973 19771 4031 19777
rect 3973 19737 3985 19771
rect 4019 19768 4031 19771
rect 4019 19740 5212 19768
rect 4019 19737 4031 19740
rect 3973 19731 4031 19737
rect 5184 19700 5212 19740
rect 5258 19728 5264 19780
rect 5316 19768 5322 19780
rect 5629 19771 5687 19777
rect 5629 19768 5641 19771
rect 5316 19740 5641 19768
rect 5316 19728 5322 19740
rect 5629 19737 5641 19740
rect 5675 19737 5687 19771
rect 5629 19731 5687 19737
rect 6822 19728 6828 19780
rect 6880 19768 6886 19780
rect 7929 19771 7987 19777
rect 7929 19768 7941 19771
rect 6880 19740 7941 19768
rect 6880 19728 6886 19740
rect 7929 19737 7941 19740
rect 7975 19737 7987 19771
rect 15378 19768 15384 19780
rect 7929 19731 7987 19737
rect 10060 19740 15384 19768
rect 5442 19700 5448 19712
rect 5184 19672 5448 19700
rect 5442 19660 5448 19672
rect 5500 19700 5506 19712
rect 5721 19703 5779 19709
rect 5721 19700 5733 19703
rect 5500 19672 5733 19700
rect 5500 19660 5506 19672
rect 5721 19669 5733 19672
rect 5767 19669 5779 19703
rect 5721 19663 5779 19669
rect 6089 19703 6147 19709
rect 6089 19669 6101 19703
rect 6135 19700 6147 19703
rect 6178 19700 6184 19712
rect 6135 19672 6184 19700
rect 6135 19669 6147 19672
rect 6089 19663 6147 19669
rect 6178 19660 6184 19672
rect 6236 19660 6242 19712
rect 6546 19660 6552 19712
rect 6604 19700 6610 19712
rect 6733 19703 6791 19709
rect 6733 19700 6745 19703
rect 6604 19672 6745 19700
rect 6604 19660 6610 19672
rect 6733 19669 6745 19672
rect 6779 19669 6791 19703
rect 6733 19663 6791 19669
rect 7101 19703 7159 19709
rect 7101 19669 7113 19703
rect 7147 19700 7159 19703
rect 7466 19700 7472 19712
rect 7147 19672 7472 19700
rect 7147 19669 7159 19672
rect 7101 19663 7159 19669
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 7558 19660 7564 19712
rect 7616 19700 7622 19712
rect 10060 19709 10088 19740
rect 15378 19728 15384 19740
rect 15436 19728 15442 19780
rect 18616 19768 18644 19799
rect 19058 19796 19064 19808
rect 19116 19836 19122 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 19116 19808 19257 19836
rect 19116 19796 19122 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 19720 19777 19748 19876
rect 21358 19836 21364 19848
rect 21319 19808 21364 19836
rect 21358 19796 21364 19808
rect 21416 19796 21422 19848
rect 18340 19740 18644 19768
rect 19705 19771 19763 19777
rect 18340 19712 18368 19740
rect 19705 19737 19717 19771
rect 19751 19768 19763 19771
rect 20162 19768 20168 19780
rect 19751 19740 20168 19768
rect 19751 19737 19763 19740
rect 19705 19731 19763 19737
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 20990 19728 20996 19780
rect 21048 19768 21054 19780
rect 21094 19771 21152 19777
rect 21094 19768 21106 19771
rect 21048 19740 21106 19768
rect 21048 19728 21054 19740
rect 21094 19737 21106 19740
rect 21140 19737 21152 19771
rect 21094 19731 21152 19737
rect 10045 19703 10103 19709
rect 7616 19672 7661 19700
rect 7616 19660 7622 19672
rect 10045 19669 10057 19703
rect 10091 19669 10103 19703
rect 10045 19663 10103 19669
rect 13722 19660 13728 19712
rect 13780 19700 13786 19712
rect 14185 19703 14243 19709
rect 14185 19700 14197 19703
rect 13780 19672 14197 19700
rect 13780 19660 13786 19672
rect 14185 19669 14197 19672
rect 14231 19700 14243 19703
rect 14461 19703 14519 19709
rect 14461 19700 14473 19703
rect 14231 19672 14473 19700
rect 14231 19669 14243 19672
rect 14185 19663 14243 19669
rect 14461 19669 14473 19672
rect 14507 19669 14519 19703
rect 14461 19663 14519 19669
rect 14642 19660 14648 19712
rect 14700 19700 14706 19712
rect 17221 19703 17279 19709
rect 17221 19700 17233 19703
rect 14700 19672 17233 19700
rect 14700 19660 14706 19672
rect 17221 19669 17233 19672
rect 17267 19669 17279 19703
rect 17221 19663 17279 19669
rect 18322 19660 18328 19712
rect 18380 19660 18386 19712
rect 19426 19660 19432 19712
rect 19484 19700 19490 19712
rect 19981 19703 20039 19709
rect 19981 19700 19993 19703
rect 19484 19672 19993 19700
rect 19484 19660 19490 19672
rect 19981 19669 19993 19672
rect 20027 19700 20039 19703
rect 20714 19700 20720 19712
rect 20027 19672 20720 19700
rect 20027 19669 20039 19672
rect 19981 19663 20039 19669
rect 20714 19660 20720 19672
rect 20772 19660 20778 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 5445 19499 5503 19505
rect 5445 19496 5457 19499
rect 5224 19468 5457 19496
rect 5224 19456 5230 19468
rect 5445 19465 5457 19468
rect 5491 19465 5503 19499
rect 5994 19496 6000 19508
rect 5955 19468 6000 19496
rect 5445 19459 5503 19465
rect 5994 19456 6000 19468
rect 6052 19456 6058 19508
rect 6546 19456 6552 19508
rect 6604 19456 6610 19508
rect 6733 19499 6791 19505
rect 6733 19465 6745 19499
rect 6779 19465 6791 19499
rect 7466 19496 7472 19508
rect 7427 19468 7472 19496
rect 6733 19459 6791 19465
rect 1578 19388 1584 19440
rect 1636 19388 1642 19440
rect 1670 19388 1676 19440
rect 1728 19428 1734 19440
rect 3605 19431 3663 19437
rect 3605 19428 3617 19431
rect 1728 19400 3617 19428
rect 1728 19388 1734 19400
rect 3605 19397 3617 19400
rect 3651 19397 3663 19431
rect 3605 19391 3663 19397
rect 4522 19388 4528 19440
rect 4580 19428 4586 19440
rect 6564 19428 6592 19456
rect 4580 19400 6592 19428
rect 4580 19388 4586 19400
rect 1596 19292 1624 19388
rect 2133 19363 2191 19369
rect 2133 19329 2145 19363
rect 2179 19360 2191 19363
rect 3418 19360 3424 19372
rect 2179 19332 3424 19360
rect 2179 19329 2191 19332
rect 2133 19323 2191 19329
rect 3418 19320 3424 19332
rect 3476 19320 3482 19372
rect 3878 19360 3884 19372
rect 3839 19332 3884 19360
rect 3878 19320 3884 19332
rect 3936 19320 3942 19372
rect 6546 19360 6552 19372
rect 6507 19332 6552 19360
rect 6546 19320 6552 19332
rect 6604 19320 6610 19372
rect 6748 19360 6776 19459
rect 7466 19456 7472 19468
rect 7524 19456 7530 19508
rect 9953 19499 10011 19505
rect 9953 19465 9965 19499
rect 9999 19496 10011 19499
rect 10597 19499 10655 19505
rect 9999 19468 10548 19496
rect 9999 19465 10011 19468
rect 9953 19459 10011 19465
rect 7377 19431 7435 19437
rect 7377 19397 7389 19431
rect 7423 19428 7435 19431
rect 7558 19428 7564 19440
rect 7423 19400 7564 19428
rect 7423 19397 7435 19400
rect 7377 19391 7435 19397
rect 7558 19388 7564 19400
rect 7616 19388 7622 19440
rect 8849 19431 8907 19437
rect 8404 19400 8800 19428
rect 8404 19360 8432 19400
rect 8570 19360 8576 19372
rect 6748 19332 8432 19360
rect 8531 19332 8576 19360
rect 8570 19320 8576 19332
rect 8628 19320 8634 19372
rect 8772 19360 8800 19400
rect 8849 19397 8861 19431
rect 8895 19428 8907 19431
rect 8895 19400 10456 19428
rect 8895 19397 8907 19400
rect 8849 19391 8907 19397
rect 8772 19332 9536 19360
rect 3050 19292 3056 19304
rect 1596 19264 3056 19292
rect 3050 19252 3056 19264
rect 3108 19252 3114 19304
rect 7285 19295 7343 19301
rect 7285 19261 7297 19295
rect 7331 19292 7343 19295
rect 7558 19292 7564 19304
rect 7331 19264 7564 19292
rect 7331 19261 7343 19264
rect 7285 19255 7343 19261
rect 7558 19252 7564 19264
rect 7616 19292 7622 19304
rect 7926 19292 7932 19304
rect 7616 19264 7932 19292
rect 7616 19252 7622 19264
rect 7926 19252 7932 19264
rect 7984 19252 7990 19304
rect 9508 19292 9536 19332
rect 9582 19320 9588 19372
rect 9640 19360 9646 19372
rect 9640 19332 9685 19360
rect 9640 19320 9646 19332
rect 9950 19320 9956 19372
rect 10008 19360 10014 19372
rect 10428 19369 10456 19400
rect 10137 19363 10195 19369
rect 10137 19360 10149 19363
rect 10008 19332 10149 19360
rect 10008 19320 10014 19332
rect 10137 19329 10149 19332
rect 10183 19329 10195 19363
rect 10137 19323 10195 19329
rect 10413 19363 10471 19369
rect 10413 19329 10425 19363
rect 10459 19329 10471 19363
rect 10520 19360 10548 19468
rect 10597 19465 10609 19499
rect 10643 19496 10655 19499
rect 13630 19496 13636 19508
rect 10643 19468 13636 19496
rect 10643 19465 10655 19468
rect 10597 19459 10655 19465
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 13722 19456 13728 19508
rect 13780 19496 13786 19508
rect 14093 19499 14151 19505
rect 13780 19468 13871 19496
rect 13780 19456 13786 19468
rect 13565 19400 13768 19428
rect 12710 19360 12716 19372
rect 10520 19332 12716 19360
rect 10413 19323 10471 19329
rect 12710 19320 12716 19332
rect 12768 19320 12774 19372
rect 12986 19320 12992 19372
rect 13044 19360 13050 19372
rect 13565 19369 13593 19400
rect 13550 19363 13608 19369
rect 13550 19360 13562 19363
rect 13044 19332 13562 19360
rect 13044 19320 13050 19332
rect 13550 19329 13562 19332
rect 13596 19329 13608 19363
rect 13550 19323 13608 19329
rect 10226 19292 10232 19304
rect 9508 19264 10232 19292
rect 10226 19252 10232 19264
rect 10284 19252 10290 19304
rect 13740 19292 13768 19400
rect 13843 19369 13871 19468
rect 14093 19465 14105 19499
rect 14139 19496 14151 19499
rect 14274 19496 14280 19508
rect 14139 19468 14280 19496
rect 14139 19465 14151 19468
rect 14093 19459 14151 19465
rect 14274 19456 14280 19468
rect 14332 19456 14338 19508
rect 17494 19456 17500 19508
rect 17552 19496 17558 19508
rect 18049 19499 18107 19505
rect 18049 19496 18061 19499
rect 17552 19468 18061 19496
rect 17552 19456 17558 19468
rect 18049 19465 18061 19468
rect 18095 19465 18107 19499
rect 18049 19459 18107 19465
rect 16758 19428 16764 19440
rect 13924 19400 16764 19428
rect 13817 19363 13875 19369
rect 13817 19329 13829 19363
rect 13863 19329 13875 19363
rect 13817 19323 13875 19329
rect 13924 19292 13952 19400
rect 16758 19388 16764 19400
rect 16816 19388 16822 19440
rect 15194 19360 15200 19372
rect 15252 19369 15258 19372
rect 15164 19332 15200 19360
rect 15194 19320 15200 19332
rect 15252 19323 15264 19369
rect 15252 19320 15258 19323
rect 16574 19320 16580 19372
rect 16632 19360 16638 19372
rect 16925 19363 16983 19369
rect 16925 19360 16937 19363
rect 16632 19332 16937 19360
rect 16632 19320 16638 19332
rect 16925 19329 16937 19332
rect 16971 19329 16983 19363
rect 16925 19323 16983 19329
rect 20806 19320 20812 19372
rect 20864 19369 20870 19372
rect 20864 19360 20876 19369
rect 20864 19332 20909 19360
rect 20864 19323 20876 19332
rect 20864 19320 20870 19323
rect 13740 19264 13952 19292
rect 15473 19295 15531 19301
rect 15473 19261 15485 19295
rect 15519 19292 15531 19295
rect 15746 19292 15752 19304
rect 15519 19264 15752 19292
rect 15519 19261 15531 19264
rect 15473 19255 15531 19261
rect 15746 19252 15752 19264
rect 15804 19292 15810 19304
rect 16669 19295 16727 19301
rect 16669 19292 16681 19295
rect 15804 19264 16681 19292
rect 15804 19252 15810 19264
rect 16669 19261 16681 19264
rect 16715 19261 16727 19295
rect 16669 19255 16727 19261
rect 18230 19252 18236 19304
rect 18288 19292 18294 19304
rect 19886 19292 19892 19304
rect 18288 19264 19892 19292
rect 18288 19252 18294 19264
rect 19886 19252 19892 19264
rect 19944 19252 19950 19304
rect 21082 19292 21088 19304
rect 21043 19264 21088 19292
rect 21082 19252 21088 19264
rect 21140 19292 21146 19304
rect 21358 19292 21364 19304
rect 21140 19264 21364 19292
rect 21140 19252 21146 19264
rect 21358 19252 21364 19264
rect 21416 19252 21422 19304
rect 5626 19224 5632 19236
rect 2746 19196 5632 19224
rect 1118 19116 1124 19168
rect 1176 19156 1182 19168
rect 2746 19156 2774 19196
rect 5626 19184 5632 19196
rect 5684 19184 5690 19236
rect 9401 19227 9459 19233
rect 9401 19193 9413 19227
rect 9447 19224 9459 19227
rect 9447 19196 12940 19224
rect 9447 19193 9459 19196
rect 9401 19187 9459 19193
rect 1176 19128 2774 19156
rect 1176 19116 1182 19128
rect 3510 19116 3516 19168
rect 3568 19156 3574 19168
rect 4246 19156 4252 19168
rect 3568 19128 4252 19156
rect 3568 19116 3574 19128
rect 4246 19116 4252 19128
rect 4304 19116 4310 19168
rect 4522 19156 4528 19168
rect 4483 19128 4528 19156
rect 4522 19116 4528 19128
rect 4580 19116 4586 19168
rect 4985 19159 5043 19165
rect 4985 19125 4997 19159
rect 5031 19156 5043 19159
rect 5258 19156 5264 19168
rect 5031 19128 5264 19156
rect 5031 19125 5043 19128
rect 4985 19119 5043 19125
rect 5258 19116 5264 19128
rect 5316 19116 5322 19168
rect 7834 19156 7840 19168
rect 7795 19128 7840 19156
rect 7834 19116 7840 19128
rect 7892 19116 7898 19168
rect 7926 19116 7932 19168
rect 7984 19156 7990 19168
rect 8113 19159 8171 19165
rect 8113 19156 8125 19159
rect 7984 19128 8125 19156
rect 7984 19116 7990 19128
rect 8113 19125 8125 19128
rect 8159 19125 8171 19159
rect 8113 19119 8171 19125
rect 12437 19159 12495 19165
rect 12437 19125 12449 19159
rect 12483 19156 12495 19159
rect 12802 19156 12808 19168
rect 12483 19128 12808 19156
rect 12483 19125 12495 19128
rect 12437 19119 12495 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 12912 19156 12940 19196
rect 13832 19196 14596 19224
rect 13832 19156 13860 19196
rect 12912 19128 13860 19156
rect 14568 19156 14596 19196
rect 17954 19184 17960 19236
rect 18012 19224 18018 19236
rect 19334 19224 19340 19236
rect 18012 19196 19340 19224
rect 18012 19184 18018 19196
rect 19334 19184 19340 19196
rect 19392 19184 19398 19236
rect 16942 19156 16948 19168
rect 14568 19128 16948 19156
rect 16942 19116 16948 19128
rect 17000 19116 17006 19168
rect 18322 19156 18328 19168
rect 18283 19128 18328 19156
rect 18322 19116 18328 19128
rect 18380 19156 18386 19168
rect 18969 19159 19027 19165
rect 18969 19156 18981 19159
rect 18380 19128 18981 19156
rect 18380 19116 18386 19128
rect 18969 19125 18981 19128
rect 19015 19125 19027 19159
rect 18969 19119 19027 19125
rect 19429 19159 19487 19165
rect 19429 19125 19441 19159
rect 19475 19156 19487 19159
rect 19610 19156 19616 19168
rect 19475 19128 19616 19156
rect 19475 19125 19487 19128
rect 19429 19119 19487 19125
rect 19610 19116 19616 19128
rect 19668 19116 19674 19168
rect 19702 19116 19708 19168
rect 19760 19156 19766 19168
rect 19760 19128 19805 19156
rect 19760 19116 19766 19128
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 2130 18912 2136 18964
rect 2188 18952 2194 18964
rect 4154 18952 4160 18964
rect 2188 18924 4160 18952
rect 2188 18912 2194 18924
rect 4154 18912 4160 18924
rect 4212 18912 4218 18964
rect 4982 18912 4988 18964
rect 5040 18952 5046 18964
rect 5445 18955 5503 18961
rect 5445 18952 5457 18955
rect 5040 18924 5457 18952
rect 5040 18912 5046 18924
rect 5445 18921 5457 18924
rect 5491 18952 5503 18955
rect 5718 18952 5724 18964
rect 5491 18924 5724 18952
rect 5491 18921 5503 18924
rect 5445 18915 5503 18921
rect 5718 18912 5724 18924
rect 5776 18912 5782 18964
rect 12434 18952 12440 18964
rect 12406 18912 12440 18952
rect 12492 18912 12498 18964
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 18598 18952 18604 18964
rect 12584 18924 18604 18952
rect 12584 18912 12590 18924
rect 18598 18912 18604 18924
rect 18656 18912 18662 18964
rect 18690 18912 18696 18964
rect 18748 18952 18754 18964
rect 22738 18952 22744 18964
rect 18748 18924 22744 18952
rect 18748 18912 18754 18924
rect 22738 18912 22744 18924
rect 22796 18912 22802 18964
rect 2314 18884 2320 18896
rect 2275 18856 2320 18884
rect 2314 18844 2320 18856
rect 2372 18844 2378 18896
rect 2958 18844 2964 18896
rect 3016 18884 3022 18896
rect 4522 18884 4528 18896
rect 3016 18856 4528 18884
rect 3016 18844 3022 18856
rect 4522 18844 4528 18856
rect 4580 18844 4586 18896
rect 12406 18884 12434 18912
rect 8404 18856 12434 18884
rect 3142 18776 3148 18828
rect 3200 18816 3206 18828
rect 6270 18816 6276 18828
rect 3200 18788 6276 18816
rect 3200 18776 3206 18788
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 6825 18819 6883 18825
rect 6825 18785 6837 18819
rect 6871 18816 6883 18819
rect 8404 18816 8432 18856
rect 15562 18844 15568 18896
rect 15620 18884 15626 18896
rect 16117 18887 16175 18893
rect 16117 18884 16129 18887
rect 15620 18856 16129 18884
rect 15620 18844 15626 18856
rect 16117 18853 16129 18856
rect 16163 18884 16175 18887
rect 16482 18884 16488 18896
rect 16163 18856 16488 18884
rect 16163 18853 16175 18856
rect 16117 18847 16175 18853
rect 16482 18844 16488 18856
rect 16540 18844 16546 18896
rect 6871 18788 8432 18816
rect 8481 18819 8539 18825
rect 6871 18785 6883 18788
rect 6825 18779 6883 18785
rect 8481 18785 8493 18819
rect 8527 18816 8539 18819
rect 12526 18816 12532 18828
rect 8527 18788 12532 18816
rect 8527 18785 8539 18788
rect 8481 18779 8539 18785
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 2501 18751 2559 18757
rect 2501 18717 2513 18751
rect 2547 18717 2559 18751
rect 2501 18711 2559 18717
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 9309 18751 9367 18757
rect 4755 18720 7880 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 2516 18680 2544 18711
rect 4433 18683 4491 18689
rect 4433 18680 4445 18683
rect 2516 18652 4445 18680
rect 4433 18649 4445 18652
rect 4479 18649 4491 18683
rect 5534 18680 5540 18692
rect 4433 18643 4491 18649
rect 4540 18652 5540 18680
rect 198 18572 204 18624
rect 256 18612 262 18624
rect 4540 18612 4568 18652
rect 5534 18640 5540 18652
rect 5592 18640 5598 18692
rect 6822 18680 6828 18692
rect 5920 18652 6828 18680
rect 5074 18612 5080 18624
rect 256 18584 4568 18612
rect 5035 18584 5080 18612
rect 256 18572 262 18584
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 5718 18572 5724 18624
rect 5776 18612 5782 18624
rect 5920 18621 5948 18652
rect 6822 18640 6828 18652
rect 6880 18680 6886 18692
rect 6917 18683 6975 18689
rect 6917 18680 6929 18683
rect 6880 18652 6929 18680
rect 6880 18640 6886 18652
rect 6917 18649 6929 18652
rect 6963 18649 6975 18683
rect 6917 18643 6975 18649
rect 5905 18615 5963 18621
rect 5905 18612 5917 18615
rect 5776 18584 5917 18612
rect 5776 18572 5782 18584
rect 5905 18581 5917 18584
rect 5951 18581 5963 18615
rect 5905 18575 5963 18581
rect 6270 18572 6276 18624
rect 6328 18612 6334 18624
rect 7009 18615 7067 18621
rect 7009 18612 7021 18615
rect 6328 18584 7021 18612
rect 6328 18572 6334 18584
rect 7009 18581 7021 18584
rect 7055 18581 7067 18615
rect 7374 18612 7380 18624
rect 7335 18584 7380 18612
rect 7009 18575 7067 18581
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 7852 18621 7880 18720
rect 9309 18717 9321 18751
rect 9355 18717 9367 18751
rect 9766 18748 9772 18760
rect 9727 18720 9772 18748
rect 9309 18711 9367 18717
rect 8110 18640 8116 18692
rect 8168 18680 8174 18692
rect 8297 18683 8355 18689
rect 8297 18680 8309 18683
rect 8168 18652 8309 18680
rect 8168 18640 8174 18652
rect 8297 18649 8309 18652
rect 8343 18649 8355 18683
rect 9324 18680 9352 18711
rect 9766 18708 9772 18720
rect 9824 18708 9830 18760
rect 10042 18748 10048 18760
rect 10003 18720 10048 18748
rect 10042 18708 10048 18720
rect 10100 18708 10106 18760
rect 10226 18708 10232 18760
rect 10284 18748 10290 18760
rect 13722 18748 13728 18760
rect 10284 18720 13584 18748
rect 13683 18720 13728 18748
rect 10284 18708 10290 18720
rect 9674 18680 9680 18692
rect 9324 18652 9680 18680
rect 8297 18643 8355 18649
rect 9674 18640 9680 18652
rect 9732 18640 9738 18692
rect 12526 18640 12532 18692
rect 12584 18680 12590 18692
rect 13262 18680 13268 18692
rect 12584 18652 13268 18680
rect 12584 18640 12590 18652
rect 13262 18640 13268 18652
rect 13320 18640 13326 18692
rect 13446 18680 13452 18692
rect 13504 18689 13510 18692
rect 13416 18652 13452 18680
rect 13446 18640 13452 18652
rect 13504 18643 13516 18689
rect 13556 18680 13584 18720
rect 13722 18708 13728 18720
rect 13780 18708 13786 18760
rect 15206 18751 15264 18757
rect 15206 18717 15218 18751
rect 15252 18717 15264 18751
rect 15206 18711 15264 18717
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18748 15531 18751
rect 15746 18748 15752 18760
rect 15519 18720 15752 18748
rect 15519 18717 15531 18720
rect 15473 18711 15531 18717
rect 14458 18680 14464 18692
rect 13556 18652 14464 18680
rect 13504 18640 13510 18643
rect 14458 18640 14464 18652
rect 14516 18640 14522 18692
rect 15212 18680 15240 18711
rect 15746 18708 15752 18720
rect 15804 18748 15810 18760
rect 17497 18751 17555 18757
rect 17497 18748 17509 18751
rect 15804 18720 17509 18748
rect 15804 18708 15810 18720
rect 17497 18717 17509 18720
rect 17543 18748 17555 18751
rect 17773 18751 17831 18757
rect 17773 18748 17785 18751
rect 17543 18720 17785 18748
rect 17543 18717 17555 18720
rect 17497 18711 17555 18717
rect 17773 18717 17785 18720
rect 17819 18748 17831 18751
rect 18322 18748 18328 18760
rect 17819 18720 18328 18748
rect 17819 18717 17831 18720
rect 17773 18711 17831 18717
rect 18322 18708 18328 18720
rect 18380 18748 18386 18760
rect 18785 18751 18843 18757
rect 18785 18748 18797 18751
rect 18380 18720 18797 18748
rect 18380 18708 18386 18720
rect 18785 18717 18797 18720
rect 18831 18748 18843 18751
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 18831 18720 19257 18748
rect 18831 18717 18843 18720
rect 18785 18711 18843 18717
rect 19245 18717 19257 18720
rect 19291 18748 19303 18751
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 19291 18720 20913 18748
rect 19291 18717 19303 18720
rect 19245 18711 19303 18717
rect 20901 18717 20913 18720
rect 20947 18748 20959 18751
rect 21082 18748 21088 18760
rect 20947 18720 21088 18748
rect 20947 18717 20959 18720
rect 20901 18711 20959 18717
rect 21082 18708 21088 18720
rect 21140 18748 21146 18760
rect 21269 18751 21327 18757
rect 21269 18748 21281 18751
rect 21140 18720 21281 18748
rect 21140 18708 21146 18720
rect 21269 18717 21281 18720
rect 21315 18717 21327 18751
rect 21269 18711 21327 18717
rect 15286 18680 15292 18692
rect 15212 18652 15292 18680
rect 15286 18640 15292 18652
rect 15344 18640 15350 18692
rect 16114 18640 16120 18692
rect 16172 18680 16178 18692
rect 17230 18683 17288 18689
rect 17230 18680 17242 18683
rect 16172 18652 17242 18680
rect 16172 18640 16178 18652
rect 17230 18649 17242 18652
rect 17276 18649 17288 18683
rect 19334 18680 19340 18692
rect 17230 18643 17288 18649
rect 18340 18652 19340 18680
rect 7837 18615 7895 18621
rect 7837 18581 7849 18615
rect 7883 18581 7895 18615
rect 8202 18612 8208 18624
rect 8163 18584 8208 18612
rect 7837 18575 7895 18581
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 9125 18615 9183 18621
rect 9125 18581 9137 18615
rect 9171 18612 9183 18615
rect 11790 18612 11796 18624
rect 9171 18584 11796 18612
rect 9171 18581 9183 18584
rect 9125 18575 9183 18581
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 12066 18572 12072 18624
rect 12124 18612 12130 18624
rect 12345 18615 12403 18621
rect 12345 18612 12357 18615
rect 12124 18584 12357 18612
rect 12124 18572 12130 18584
rect 12345 18581 12357 18584
rect 12391 18581 12403 18615
rect 12345 18575 12403 18581
rect 12710 18572 12716 18624
rect 12768 18612 12774 18624
rect 14093 18615 14151 18621
rect 14093 18612 14105 18615
rect 12768 18584 14105 18612
rect 12768 18572 12774 18584
rect 14093 18581 14105 18584
rect 14139 18581 14151 18615
rect 14093 18575 14151 18581
rect 14182 18572 14188 18624
rect 14240 18612 14246 18624
rect 18340 18612 18368 18652
rect 19334 18640 19340 18652
rect 19392 18640 19398 18692
rect 19512 18683 19570 18689
rect 19512 18680 19524 18683
rect 19444 18652 19524 18680
rect 14240 18584 18368 18612
rect 14240 18572 14246 18584
rect 18414 18572 18420 18624
rect 18472 18612 18478 18624
rect 19444 18612 19472 18652
rect 19512 18649 19524 18652
rect 19558 18680 19570 18683
rect 19702 18680 19708 18692
rect 19558 18652 19708 18680
rect 19558 18649 19570 18652
rect 19512 18643 19570 18649
rect 19702 18640 19708 18652
rect 19760 18640 19766 18692
rect 18472 18584 19472 18612
rect 18472 18572 18478 18584
rect 20254 18572 20260 18624
rect 20312 18612 20318 18624
rect 20625 18615 20683 18621
rect 20625 18612 20637 18615
rect 20312 18584 20637 18612
rect 20312 18572 20318 18584
rect 20625 18581 20637 18584
rect 20671 18581 20683 18615
rect 20625 18575 20683 18581
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 5077 18411 5135 18417
rect 5077 18408 5089 18411
rect 4212 18380 5089 18408
rect 4212 18368 4218 18380
rect 5077 18377 5089 18380
rect 5123 18408 5135 18411
rect 5350 18408 5356 18420
rect 5123 18380 5356 18408
rect 5123 18377 5135 18380
rect 5077 18371 5135 18377
rect 5350 18368 5356 18380
rect 5408 18368 5414 18420
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 6365 18411 6423 18417
rect 6365 18408 6377 18411
rect 5960 18380 6377 18408
rect 5960 18368 5966 18380
rect 6365 18377 6377 18380
rect 6411 18408 6423 18411
rect 6822 18408 6828 18420
rect 6411 18380 6828 18408
rect 6411 18377 6423 18380
rect 6365 18371 6423 18377
rect 6822 18368 6828 18380
rect 6880 18368 6886 18420
rect 7561 18411 7619 18417
rect 7561 18377 7573 18411
rect 7607 18408 7619 18411
rect 7834 18408 7840 18420
rect 7607 18380 7840 18408
rect 7607 18377 7619 18380
rect 7561 18371 7619 18377
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 8202 18368 8208 18420
rect 8260 18408 8266 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 8260 18380 8309 18408
rect 8260 18368 8266 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 10873 18411 10931 18417
rect 10873 18408 10885 18411
rect 8297 18371 8355 18377
rect 9140 18380 10885 18408
rect 2498 18340 2504 18352
rect 2459 18312 2504 18340
rect 2498 18300 2504 18312
rect 2556 18300 2562 18352
rect 3418 18300 3424 18352
rect 3476 18340 3482 18352
rect 4065 18343 4123 18349
rect 4065 18340 4077 18343
rect 3476 18312 4077 18340
rect 3476 18300 3482 18312
rect 4065 18309 4077 18312
rect 4111 18309 4123 18343
rect 4065 18303 4123 18309
rect 7374 18300 7380 18352
rect 7432 18340 7438 18352
rect 9140 18340 9168 18380
rect 10873 18377 10885 18380
rect 10919 18377 10931 18411
rect 12434 18408 12440 18420
rect 10873 18371 10931 18377
rect 11716 18380 12440 18408
rect 7432 18312 9168 18340
rect 9677 18343 9735 18349
rect 7432 18300 7438 18312
rect 9677 18309 9689 18343
rect 9723 18340 9735 18343
rect 10134 18340 10140 18352
rect 9723 18312 10140 18340
rect 9723 18309 9735 18312
rect 9677 18303 9735 18309
rect 10134 18300 10140 18312
rect 10192 18300 10198 18352
rect 2774 18232 2780 18284
rect 2832 18272 2838 18284
rect 4341 18275 4399 18281
rect 2832 18244 2877 18272
rect 2832 18232 2838 18244
rect 4341 18241 4353 18275
rect 4387 18272 4399 18275
rect 5442 18272 5448 18284
rect 4387 18244 5448 18272
rect 4387 18241 4399 18244
rect 4341 18235 4399 18241
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 7650 18272 7656 18284
rect 7611 18244 7656 18272
rect 7650 18232 7656 18244
rect 7708 18232 7714 18284
rect 9398 18272 9404 18284
rect 9359 18244 9404 18272
rect 9398 18232 9404 18244
rect 9456 18232 9462 18284
rect 10778 18272 10784 18284
rect 10739 18244 10784 18272
rect 10778 18232 10784 18244
rect 10836 18232 10842 18284
rect 4430 18164 4436 18216
rect 4488 18204 4494 18216
rect 4617 18207 4675 18213
rect 4617 18204 4629 18207
rect 4488 18176 4629 18204
rect 4488 18164 4494 18176
rect 4617 18173 4629 18176
rect 4663 18173 4675 18207
rect 4617 18167 4675 18173
rect 4706 18164 4712 18216
rect 4764 18204 4770 18216
rect 7469 18207 7527 18213
rect 4764 18176 6960 18204
rect 4764 18164 4770 18176
rect 3234 18136 3240 18148
rect 3195 18108 3240 18136
rect 3234 18096 3240 18108
rect 3292 18096 3298 18148
rect 3418 18096 3424 18148
rect 3476 18136 3482 18148
rect 4798 18136 4804 18148
rect 3476 18108 4804 18136
rect 3476 18096 3482 18108
rect 4798 18096 4804 18108
rect 4856 18096 4862 18148
rect 6932 18136 6960 18176
rect 7469 18173 7481 18207
rect 7515 18204 7527 18207
rect 7834 18204 7840 18216
rect 7515 18176 7840 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 7834 18164 7840 18176
rect 7892 18164 7898 18216
rect 10965 18207 11023 18213
rect 10965 18173 10977 18207
rect 11011 18204 11023 18207
rect 11716 18204 11744 18380
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 12526 18368 12532 18420
rect 12584 18408 12590 18420
rect 14093 18411 14151 18417
rect 14093 18408 14105 18411
rect 12584 18380 14105 18408
rect 12584 18368 12590 18380
rect 14093 18377 14105 18380
rect 14139 18408 14151 18411
rect 15194 18408 15200 18420
rect 14139 18380 15200 18408
rect 14139 18377 14151 18380
rect 14093 18371 14151 18377
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 15378 18368 15384 18420
rect 15436 18408 15442 18420
rect 20990 18408 20996 18420
rect 15436 18380 20996 18408
rect 15436 18368 15442 18380
rect 20990 18368 20996 18380
rect 21048 18408 21054 18420
rect 21361 18411 21419 18417
rect 21361 18408 21373 18411
rect 21048 18380 21373 18408
rect 21048 18368 21054 18380
rect 21361 18377 21373 18380
rect 21407 18377 21419 18411
rect 21361 18371 21419 18377
rect 11790 18300 11796 18352
rect 11848 18340 11854 18352
rect 11848 18312 12664 18340
rect 11848 18300 11854 18312
rect 12636 18272 12664 18312
rect 12710 18300 12716 18352
rect 12768 18340 12774 18352
rect 12958 18343 13016 18349
rect 12958 18340 12970 18343
rect 12768 18312 12970 18340
rect 12768 18300 12774 18312
rect 12958 18309 12970 18312
rect 13004 18309 13016 18343
rect 17678 18340 17684 18352
rect 12958 18303 13016 18309
rect 13096 18312 17684 18340
rect 13096 18272 13124 18312
rect 17678 18300 17684 18312
rect 17736 18300 17742 18352
rect 18064 18312 19748 18340
rect 12636 18244 13124 18272
rect 13446 18232 13452 18284
rect 13504 18272 13510 18284
rect 13504 18244 14412 18272
rect 13504 18232 13510 18244
rect 11011 18176 11744 18204
rect 12713 18207 12771 18213
rect 11011 18173 11023 18176
rect 10965 18167 11023 18173
rect 12713 18173 12725 18207
rect 12759 18173 12771 18207
rect 12713 18167 12771 18173
rect 8021 18139 8079 18145
rect 6932 18108 7052 18136
rect 3605 18071 3663 18077
rect 3605 18037 3617 18071
rect 3651 18068 3663 18071
rect 4890 18068 4896 18080
rect 3651 18040 4896 18068
rect 3651 18037 3663 18040
rect 3605 18031 3663 18037
rect 4890 18028 4896 18040
rect 4948 18028 4954 18080
rect 5626 18068 5632 18080
rect 5587 18040 5632 18068
rect 5626 18028 5632 18040
rect 5684 18028 5690 18080
rect 5997 18071 6055 18077
rect 5997 18037 6009 18071
rect 6043 18068 6055 18071
rect 6086 18068 6092 18080
rect 6043 18040 6092 18068
rect 6043 18037 6055 18040
rect 5997 18031 6055 18037
rect 6086 18028 6092 18040
rect 6144 18028 6150 18080
rect 6914 18068 6920 18080
rect 6875 18040 6920 18068
rect 6914 18028 6920 18040
rect 6972 18028 6978 18080
rect 7024 18068 7052 18108
rect 8021 18105 8033 18139
rect 8067 18136 8079 18139
rect 8570 18136 8576 18148
rect 8067 18108 8576 18136
rect 8067 18105 8079 18108
rect 8021 18099 8079 18105
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 8662 18068 8668 18080
rect 7024 18040 8668 18068
rect 8662 18028 8668 18040
rect 8720 18068 8726 18080
rect 8757 18071 8815 18077
rect 8757 18068 8769 18071
rect 8720 18040 8769 18068
rect 8720 18028 8726 18040
rect 8757 18037 8769 18040
rect 8803 18037 8815 18071
rect 8757 18031 8815 18037
rect 10413 18071 10471 18077
rect 10413 18037 10425 18071
rect 10459 18068 10471 18071
rect 10502 18068 10508 18080
rect 10459 18040 10508 18068
rect 10459 18037 10471 18040
rect 10413 18031 10471 18037
rect 10502 18028 10508 18040
rect 10560 18028 10566 18080
rect 10870 18028 10876 18080
rect 10928 18068 10934 18080
rect 11790 18068 11796 18080
rect 10928 18040 11796 18068
rect 10928 18028 10934 18040
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 12437 18071 12495 18077
rect 12437 18037 12449 18071
rect 12483 18068 12495 18071
rect 12728 18068 12756 18167
rect 14384 18145 14412 18244
rect 15470 18232 15476 18284
rect 15528 18281 15534 18284
rect 15528 18272 15540 18281
rect 15528 18244 15573 18272
rect 15528 18235 15540 18244
rect 15528 18232 15534 18235
rect 17494 18232 17500 18284
rect 17552 18272 17558 18284
rect 17770 18272 17776 18284
rect 17828 18281 17834 18284
rect 17552 18244 17776 18272
rect 17552 18232 17558 18244
rect 17770 18232 17776 18244
rect 17828 18272 17840 18281
rect 17828 18244 17873 18272
rect 17828 18235 17840 18244
rect 17828 18232 17834 18235
rect 18064 18216 18092 18312
rect 19449 18275 19507 18281
rect 19449 18241 19461 18275
rect 19495 18272 19507 18275
rect 19610 18272 19616 18284
rect 19495 18244 19616 18272
rect 19495 18241 19507 18244
rect 19449 18235 19507 18241
rect 19610 18232 19616 18244
rect 19668 18232 19674 18284
rect 19720 18281 19748 18312
rect 20254 18281 20260 18284
rect 19705 18275 19763 18281
rect 19705 18241 19717 18275
rect 19751 18272 19763 18275
rect 19981 18275 20039 18281
rect 19981 18272 19993 18275
rect 19751 18244 19993 18272
rect 19751 18241 19763 18244
rect 19705 18235 19763 18241
rect 19981 18241 19993 18244
rect 20027 18241 20039 18275
rect 20248 18272 20260 18281
rect 20215 18244 20260 18272
rect 19981 18235 20039 18241
rect 20248 18235 20260 18244
rect 20254 18232 20260 18235
rect 20312 18232 20318 18284
rect 15749 18207 15807 18213
rect 15749 18173 15761 18207
rect 15795 18173 15807 18207
rect 18046 18204 18052 18216
rect 18007 18176 18052 18204
rect 15749 18167 15807 18173
rect 14369 18139 14427 18145
rect 14369 18105 14381 18139
rect 14415 18105 14427 18139
rect 14369 18099 14427 18105
rect 15764 18080 15792 18167
rect 18046 18164 18052 18176
rect 18104 18164 18110 18216
rect 16669 18139 16727 18145
rect 16669 18105 16681 18139
rect 16715 18136 16727 18139
rect 16942 18136 16948 18148
rect 16715 18108 16948 18136
rect 16715 18105 16727 18108
rect 16669 18099 16727 18105
rect 16942 18096 16948 18108
rect 17000 18096 17006 18148
rect 13722 18068 13728 18080
rect 12483 18040 13728 18068
rect 12483 18037 12495 18040
rect 12437 18031 12495 18037
rect 13722 18028 13728 18040
rect 13780 18028 13786 18080
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 15562 18068 15568 18080
rect 13872 18040 15568 18068
rect 13872 18028 13878 18040
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 15746 18028 15752 18080
rect 15804 18068 15810 18080
rect 16025 18071 16083 18077
rect 16025 18068 16037 18071
rect 15804 18040 16037 18068
rect 15804 18028 15810 18040
rect 16025 18037 16037 18040
rect 16071 18037 16083 18071
rect 16025 18031 16083 18037
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 18325 18071 18383 18077
rect 18325 18068 18337 18071
rect 16172 18040 18337 18068
rect 16172 18028 16178 18040
rect 18325 18037 18337 18040
rect 18371 18037 18383 18071
rect 18325 18031 18383 18037
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 2501 17867 2559 17873
rect 2501 17833 2513 17867
rect 2547 17864 2559 17867
rect 2866 17864 2872 17876
rect 2547 17836 2872 17864
rect 2547 17833 2559 17836
rect 2501 17827 2559 17833
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 3878 17824 3884 17876
rect 3936 17864 3942 17876
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3936 17836 4077 17864
rect 3936 17824 3942 17836
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 4522 17824 4528 17876
rect 4580 17864 4586 17876
rect 4706 17864 4712 17876
rect 4580 17836 4712 17864
rect 4580 17824 4586 17836
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 5442 17864 5448 17876
rect 5403 17836 5448 17864
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 7098 17864 7104 17876
rect 7059 17836 7104 17864
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 12250 17824 12256 17876
rect 12308 17864 12314 17876
rect 12526 17864 12532 17876
rect 12308 17836 12532 17864
rect 12308 17824 12314 17836
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 20254 17864 20260 17876
rect 12820 17836 20260 17864
rect 5074 17756 5080 17808
rect 5132 17796 5138 17808
rect 5132 17768 11376 17796
rect 5132 17756 5138 17768
rect 4709 17731 4767 17737
rect 4709 17697 4721 17731
rect 4755 17728 4767 17731
rect 5258 17728 5264 17740
rect 4755 17700 5264 17728
rect 4755 17697 4767 17700
rect 4709 17691 4767 17697
rect 5258 17688 5264 17700
rect 5316 17688 5322 17740
rect 6086 17728 6092 17740
rect 6047 17700 6092 17728
rect 6086 17688 6092 17700
rect 6144 17688 6150 17740
rect 8021 17731 8079 17737
rect 8021 17697 8033 17731
rect 8067 17728 8079 17731
rect 9030 17728 9036 17740
rect 8067 17700 9036 17728
rect 8067 17697 8079 17700
rect 8021 17691 8079 17697
rect 9030 17688 9036 17700
rect 9088 17688 9094 17740
rect 9306 17688 9312 17740
rect 9364 17728 9370 17740
rect 9585 17731 9643 17737
rect 9585 17728 9597 17731
rect 9364 17700 9597 17728
rect 9364 17688 9370 17700
rect 9585 17697 9597 17700
rect 9631 17728 9643 17731
rect 10873 17731 10931 17737
rect 9631 17700 10088 17728
rect 9631 17697 9643 17700
rect 9585 17691 9643 17697
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17629 2191 17663
rect 2682 17660 2688 17672
rect 2643 17632 2688 17660
rect 2133 17623 2191 17629
rect 2148 17592 2176 17623
rect 2682 17620 2688 17632
rect 2740 17620 2746 17672
rect 4430 17660 4436 17672
rect 4391 17632 4436 17660
rect 4430 17620 4436 17632
rect 4488 17620 4494 17672
rect 4890 17620 4896 17672
rect 4948 17660 4954 17672
rect 8662 17660 8668 17672
rect 4948 17632 8668 17660
rect 4948 17620 4954 17632
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 8754 17620 8760 17672
rect 8812 17660 8818 17672
rect 8812 17632 9536 17660
rect 8812 17620 8818 17632
rect 4062 17592 4068 17604
rect 2148 17564 4068 17592
rect 4062 17552 4068 17564
rect 4120 17552 4126 17604
rect 5813 17595 5871 17601
rect 5813 17561 5825 17595
rect 5859 17592 5871 17595
rect 6457 17595 6515 17601
rect 6457 17592 6469 17595
rect 5859 17564 6469 17592
rect 5859 17561 5871 17564
rect 5813 17555 5871 17561
rect 6457 17561 6469 17564
rect 6503 17561 6515 17595
rect 6457 17555 6515 17561
rect 7282 17552 7288 17604
rect 7340 17592 7346 17604
rect 8205 17595 8263 17601
rect 8205 17592 8217 17595
rect 7340 17564 8217 17592
rect 7340 17552 7346 17564
rect 8205 17561 8217 17564
rect 8251 17561 8263 17595
rect 8205 17555 8263 17561
rect 8846 17552 8852 17604
rect 8904 17592 8910 17604
rect 9401 17595 9459 17601
rect 9401 17592 9413 17595
rect 8904 17564 9413 17592
rect 8904 17552 8910 17564
rect 9401 17561 9413 17564
rect 9447 17561 9459 17595
rect 9401 17555 9459 17561
rect 3421 17527 3479 17533
rect 3421 17493 3433 17527
rect 3467 17524 3479 17527
rect 3602 17524 3608 17536
rect 3467 17496 3608 17524
rect 3467 17493 3479 17496
rect 3421 17487 3479 17493
rect 3602 17484 3608 17496
rect 3660 17484 3666 17536
rect 4522 17484 4528 17536
rect 4580 17524 4586 17536
rect 5166 17524 5172 17536
rect 4580 17496 4625 17524
rect 5127 17496 5172 17524
rect 4580 17484 4586 17496
rect 5166 17484 5172 17496
rect 5224 17484 5230 17536
rect 5902 17484 5908 17536
rect 5960 17524 5966 17536
rect 7561 17527 7619 17533
rect 5960 17496 6005 17524
rect 5960 17484 5966 17496
rect 7561 17493 7573 17527
rect 7607 17524 7619 17527
rect 7926 17524 7932 17536
rect 7607 17496 7932 17524
rect 7607 17493 7619 17496
rect 7561 17487 7619 17493
rect 7926 17484 7932 17496
rect 7984 17484 7990 17536
rect 8018 17484 8024 17536
rect 8076 17524 8082 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 8076 17496 8125 17524
rect 8076 17484 8082 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 8570 17524 8576 17536
rect 8531 17496 8576 17524
rect 8113 17487 8171 17493
rect 8570 17484 8576 17496
rect 8628 17484 8634 17536
rect 8938 17524 8944 17536
rect 8899 17496 8944 17524
rect 8938 17484 8944 17496
rect 8996 17484 9002 17536
rect 9309 17527 9367 17533
rect 9309 17493 9321 17527
rect 9355 17524 9367 17527
rect 9508 17524 9536 17632
rect 10060 17533 10088 17700
rect 10873 17697 10885 17731
rect 10919 17728 10931 17731
rect 11238 17728 11244 17740
rect 10919 17700 11244 17728
rect 10919 17697 10931 17700
rect 10873 17691 10931 17697
rect 11238 17688 11244 17700
rect 11296 17688 11302 17740
rect 11348 17728 11376 17768
rect 12434 17756 12440 17808
rect 12492 17796 12498 17808
rect 12820 17796 12848 17836
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 12492 17768 12848 17796
rect 12492 17756 12498 17768
rect 14458 17728 14464 17740
rect 11348 17700 12434 17728
rect 10597 17663 10655 17669
rect 10597 17629 10609 17663
rect 10643 17629 10655 17663
rect 10597 17623 10655 17629
rect 10612 17592 10640 17623
rect 10778 17620 10784 17672
rect 10836 17660 10842 17672
rect 11333 17663 11391 17669
rect 11333 17660 11345 17663
rect 10836 17632 11345 17660
rect 10836 17620 10842 17632
rect 11333 17629 11345 17632
rect 11379 17629 11391 17663
rect 12406 17660 12434 17700
rect 13924 17700 14464 17728
rect 13722 17660 13728 17672
rect 12406 17632 13584 17660
rect 13683 17632 13728 17660
rect 11333 17623 11391 17629
rect 11146 17592 11152 17604
rect 10612 17564 11152 17592
rect 11146 17552 11152 17564
rect 11204 17552 11210 17604
rect 11238 17552 11244 17604
rect 11296 17592 11302 17604
rect 12066 17592 12072 17604
rect 11296 17564 12072 17592
rect 11296 17552 11302 17564
rect 12066 17552 12072 17564
rect 12124 17592 12130 17604
rect 13458 17595 13516 17601
rect 13458 17592 13470 17595
rect 12124 17564 13470 17592
rect 12124 17552 12130 17564
rect 13458 17561 13470 17564
rect 13504 17561 13516 17595
rect 13556 17592 13584 17632
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 13924 17592 13952 17700
rect 14458 17688 14464 17700
rect 14516 17688 14522 17740
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 19610 17728 19616 17740
rect 17184 17700 19616 17728
rect 17184 17688 17190 17700
rect 19610 17688 19616 17700
rect 19668 17688 19674 17740
rect 15473 17663 15531 17669
rect 13556 17564 13952 17592
rect 14016 17632 15332 17660
rect 13458 17555 13516 17561
rect 9355 17496 9536 17524
rect 10045 17527 10103 17533
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 10045 17493 10057 17527
rect 10091 17524 10103 17527
rect 11882 17524 11888 17536
rect 10091 17496 11888 17524
rect 10091 17493 10103 17496
rect 10045 17487 10103 17493
rect 11882 17484 11888 17496
rect 11940 17484 11946 17536
rect 12345 17527 12403 17533
rect 12345 17493 12357 17527
rect 12391 17524 12403 17527
rect 12618 17524 12624 17536
rect 12391 17496 12624 17524
rect 12391 17493 12403 17496
rect 12345 17487 12403 17493
rect 12618 17484 12624 17496
rect 12676 17484 12682 17536
rect 13262 17484 13268 17536
rect 13320 17524 13326 17536
rect 14016 17524 14044 17632
rect 14734 17552 14740 17604
rect 14792 17592 14798 17604
rect 15206 17595 15264 17601
rect 15206 17592 15218 17595
rect 14792 17564 15218 17592
rect 14792 17552 14798 17564
rect 15206 17561 15218 17564
rect 15252 17561 15264 17595
rect 15206 17555 15264 17561
rect 15304 17536 15332 17632
rect 15473 17629 15485 17663
rect 15519 17660 15531 17663
rect 16117 17663 16175 17669
rect 16117 17660 16129 17663
rect 15519 17632 16129 17660
rect 15519 17629 15531 17632
rect 15473 17623 15531 17629
rect 15764 17536 15792 17632
rect 16117 17629 16129 17632
rect 16163 17629 16175 17663
rect 16117 17623 16175 17629
rect 20714 17620 20720 17672
rect 20772 17660 20778 17672
rect 21094 17663 21152 17669
rect 21094 17660 21106 17663
rect 20772 17632 21106 17660
rect 20772 17620 20778 17632
rect 21094 17629 21106 17632
rect 21140 17629 21152 17663
rect 21358 17660 21364 17672
rect 21319 17632 21364 17660
rect 21094 17623 21152 17629
rect 21358 17620 21364 17632
rect 21416 17620 21422 17672
rect 15838 17552 15844 17604
rect 15896 17592 15902 17604
rect 16362 17595 16420 17601
rect 16362 17592 16374 17595
rect 15896 17564 16374 17592
rect 15896 17552 15902 17564
rect 16362 17561 16374 17564
rect 16408 17561 16420 17595
rect 20806 17592 20812 17604
rect 16362 17555 16420 17561
rect 17512 17564 20812 17592
rect 13320 17496 14044 17524
rect 14093 17527 14151 17533
rect 13320 17484 13326 17496
rect 14093 17493 14105 17527
rect 14139 17524 14151 17527
rect 14550 17524 14556 17536
rect 14139 17496 14556 17524
rect 14139 17493 14151 17496
rect 14093 17487 14151 17493
rect 14550 17484 14556 17496
rect 14608 17484 14614 17536
rect 15286 17484 15292 17536
rect 15344 17484 15350 17536
rect 15746 17524 15752 17536
rect 15707 17496 15752 17524
rect 15746 17484 15752 17496
rect 15804 17484 15810 17536
rect 17402 17484 17408 17536
rect 17460 17524 17466 17536
rect 17512 17533 17540 17564
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 17497 17527 17555 17533
rect 17497 17524 17509 17527
rect 17460 17496 17509 17524
rect 17460 17484 17466 17496
rect 17497 17493 17509 17496
rect 17543 17493 17555 17527
rect 17497 17487 17555 17493
rect 17865 17527 17923 17533
rect 17865 17493 17877 17527
rect 17911 17524 17923 17527
rect 18046 17524 18052 17536
rect 17911 17496 18052 17524
rect 17911 17493 17923 17496
rect 17865 17487 17923 17493
rect 18046 17484 18052 17496
rect 18104 17524 18110 17536
rect 18141 17527 18199 17533
rect 18141 17524 18153 17527
rect 18104 17496 18153 17524
rect 18104 17484 18110 17496
rect 18141 17493 18153 17496
rect 18187 17524 18199 17527
rect 18877 17527 18935 17533
rect 18877 17524 18889 17527
rect 18187 17496 18889 17524
rect 18187 17493 18199 17496
rect 18141 17487 18199 17493
rect 18877 17493 18889 17496
rect 18923 17524 18935 17527
rect 19058 17524 19064 17536
rect 18923 17496 19064 17524
rect 18923 17493 18935 17496
rect 18877 17487 18935 17493
rect 19058 17484 19064 17496
rect 19116 17524 19122 17536
rect 19245 17527 19303 17533
rect 19245 17524 19257 17527
rect 19116 17496 19257 17524
rect 19116 17484 19122 17496
rect 19245 17493 19257 17496
rect 19291 17493 19303 17527
rect 19245 17487 19303 17493
rect 19702 17484 19708 17536
rect 19760 17524 19766 17536
rect 19981 17527 20039 17533
rect 19981 17524 19993 17527
rect 19760 17496 19993 17524
rect 19760 17484 19766 17496
rect 19981 17493 19993 17496
rect 20027 17493 20039 17527
rect 19981 17487 20039 17493
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 2774 17280 2780 17332
rect 2832 17320 2838 17332
rect 3237 17323 3295 17329
rect 3237 17320 3249 17323
rect 2832 17292 3249 17320
rect 2832 17280 2838 17292
rect 3237 17289 3249 17292
rect 3283 17289 3295 17323
rect 3602 17320 3608 17332
rect 3563 17292 3608 17320
rect 3237 17283 3295 17289
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 4522 17320 4528 17332
rect 4483 17292 4528 17320
rect 4522 17280 4528 17292
rect 4580 17280 4586 17332
rect 4982 17320 4988 17332
rect 4943 17292 4988 17320
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 6365 17323 6423 17329
rect 6365 17320 6377 17323
rect 5960 17292 6377 17320
rect 5960 17280 5966 17292
rect 6365 17289 6377 17292
rect 6411 17289 6423 17323
rect 6822 17320 6828 17332
rect 6783 17292 6828 17320
rect 6365 17283 6423 17289
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 7561 17323 7619 17329
rect 7561 17289 7573 17323
rect 7607 17320 7619 17323
rect 7650 17320 7656 17332
rect 7607 17292 7656 17320
rect 7607 17289 7619 17292
rect 7561 17283 7619 17289
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 7926 17320 7932 17332
rect 7887 17292 7932 17320
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 8021 17323 8079 17329
rect 8021 17289 8033 17323
rect 8067 17320 8079 17323
rect 8938 17320 8944 17332
rect 8067 17292 8944 17320
rect 8067 17289 8079 17292
rect 8021 17283 8079 17289
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 9030 17280 9036 17332
rect 9088 17320 9094 17332
rect 17402 17320 17408 17332
rect 9088 17292 17408 17320
rect 9088 17280 9094 17292
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 20898 17280 20904 17332
rect 20956 17320 20962 17332
rect 21542 17320 21548 17332
rect 20956 17292 21548 17320
rect 20956 17280 20962 17292
rect 21542 17280 21548 17292
rect 21600 17280 21606 17332
rect 2682 17252 2688 17264
rect 2643 17224 2688 17252
rect 2682 17212 2688 17224
rect 2740 17212 2746 17264
rect 4890 17252 4896 17264
rect 4851 17224 4896 17252
rect 4890 17212 4896 17224
rect 4948 17212 4954 17264
rect 5166 17212 5172 17264
rect 5224 17252 5230 17264
rect 5813 17255 5871 17261
rect 5224 17224 5764 17252
rect 5224 17212 5230 17224
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17184 2191 17187
rect 2866 17184 2872 17196
rect 2179 17156 2872 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 2961 17187 3019 17193
rect 2961 17153 2973 17187
rect 3007 17184 3019 17187
rect 4154 17184 4160 17196
rect 3007 17156 4160 17184
rect 3007 17153 3019 17156
rect 2961 17147 3019 17153
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 5534 17184 5540 17196
rect 5495 17156 5540 17184
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 5736 17184 5764 17224
rect 5813 17221 5825 17255
rect 5859 17252 5871 17255
rect 7006 17252 7012 17264
rect 5859 17224 7012 17252
rect 5859 17221 5871 17224
rect 5813 17215 5871 17221
rect 7006 17212 7012 17224
rect 7064 17212 7070 17264
rect 8846 17212 8852 17264
rect 8904 17252 8910 17264
rect 9217 17255 9275 17261
rect 8904 17224 9076 17252
rect 8904 17212 8910 17224
rect 6733 17187 6791 17193
rect 6733 17184 6745 17187
rect 5736 17156 6745 17184
rect 6733 17153 6745 17156
rect 6779 17184 6791 17187
rect 6779 17156 8524 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 3326 17076 3332 17128
rect 3384 17116 3390 17128
rect 3697 17119 3755 17125
rect 3697 17116 3709 17119
rect 3384 17088 3709 17116
rect 3384 17076 3390 17088
rect 3697 17085 3709 17088
rect 3743 17085 3755 17119
rect 3697 17079 3755 17085
rect 3789 17119 3847 17125
rect 3789 17085 3801 17119
rect 3835 17085 3847 17119
rect 5166 17116 5172 17128
rect 5127 17088 5172 17116
rect 3789 17079 3847 17085
rect 3234 17008 3240 17060
rect 3292 17048 3298 17060
rect 3804 17048 3832 17079
rect 5166 17076 5172 17088
rect 5224 17116 5230 17128
rect 5626 17116 5632 17128
rect 5224 17088 5632 17116
rect 5224 17076 5230 17088
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 5902 17076 5908 17128
rect 5960 17116 5966 17128
rect 6914 17116 6920 17128
rect 5960 17088 6920 17116
rect 5960 17076 5966 17088
rect 6914 17076 6920 17088
rect 6972 17076 6978 17128
rect 7558 17076 7564 17128
rect 7616 17116 7622 17128
rect 8113 17119 8171 17125
rect 8113 17116 8125 17119
rect 7616 17088 8125 17116
rect 7616 17076 7622 17088
rect 8113 17085 8125 17088
rect 8159 17085 8171 17119
rect 8496 17116 8524 17156
rect 8570 17144 8576 17196
rect 8628 17184 8634 17196
rect 8941 17187 8999 17193
rect 8941 17184 8953 17187
rect 8628 17156 8953 17184
rect 8628 17144 8634 17156
rect 8941 17153 8953 17156
rect 8987 17153 8999 17187
rect 9048 17184 9076 17224
rect 9217 17221 9229 17255
rect 9263 17252 9275 17255
rect 9490 17252 9496 17264
rect 9263 17224 9496 17252
rect 9263 17221 9275 17224
rect 9217 17215 9275 17221
rect 9490 17212 9496 17224
rect 9548 17212 9554 17264
rect 9861 17255 9919 17261
rect 9861 17252 9873 17255
rect 9646 17224 9873 17252
rect 9306 17184 9312 17196
rect 9048 17156 9312 17184
rect 8941 17147 8999 17153
rect 9306 17144 9312 17156
rect 9364 17184 9370 17196
rect 9646 17184 9674 17224
rect 9861 17221 9873 17224
rect 9907 17252 9919 17255
rect 10594 17252 10600 17264
rect 9907 17224 10600 17252
rect 9907 17221 9919 17224
rect 9861 17215 9919 17221
rect 10594 17212 10600 17224
rect 10652 17212 10658 17264
rect 11698 17212 11704 17264
rect 11756 17252 11762 17264
rect 12342 17252 12348 17264
rect 11756 17224 12348 17252
rect 11756 17212 11762 17224
rect 12342 17212 12348 17224
rect 12400 17212 12406 17264
rect 14458 17212 14464 17264
rect 14516 17252 14522 17264
rect 17218 17252 17224 17264
rect 14516 17224 17224 17252
rect 14516 17212 14522 17224
rect 17218 17212 17224 17224
rect 17276 17212 17282 17264
rect 19610 17212 19616 17264
rect 19668 17252 19674 17264
rect 21094 17255 21152 17261
rect 21094 17252 21106 17255
rect 19668 17224 21106 17252
rect 19668 17212 19674 17224
rect 21094 17221 21106 17224
rect 21140 17221 21152 17255
rect 21094 17215 21152 17221
rect 9364 17156 9674 17184
rect 9364 17144 9370 17156
rect 13354 17144 13360 17196
rect 13412 17193 13418 17196
rect 13412 17184 13424 17193
rect 14274 17184 14280 17196
rect 13412 17156 14280 17184
rect 13412 17147 13424 17156
rect 13412 17144 13418 17147
rect 14274 17144 14280 17156
rect 14332 17144 14338 17196
rect 17856 17187 17914 17193
rect 17856 17153 17868 17187
rect 17902 17184 17914 17187
rect 18138 17184 18144 17196
rect 17902 17156 18144 17184
rect 17902 17153 17914 17156
rect 17856 17147 17914 17153
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 10594 17116 10600 17128
rect 8496 17088 10600 17116
rect 8113 17079 8171 17085
rect 3292 17020 3832 17048
rect 3292 17008 3298 17020
rect 8128 16980 8156 17079
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 10870 17116 10876 17128
rect 10831 17088 10876 17116
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 13633 17119 13691 17125
rect 13633 17085 13645 17119
rect 13679 17116 13691 17119
rect 13722 17116 13728 17128
rect 13679 17088 13728 17116
rect 13679 17085 13691 17088
rect 13633 17079 13691 17085
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 17589 17119 17647 17125
rect 17589 17116 17601 17119
rect 17236 17088 17601 17116
rect 8202 17008 8208 17060
rect 8260 17048 8266 17060
rect 10137 17051 10195 17057
rect 10137 17048 10149 17051
rect 8260 17020 10149 17048
rect 8260 17008 8266 17020
rect 10137 17017 10149 17020
rect 10183 17017 10195 17051
rect 10137 17011 10195 17017
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 12253 17051 12311 17057
rect 12253 17048 12265 17051
rect 10836 17020 12265 17048
rect 10836 17008 10842 17020
rect 12253 17017 12265 17020
rect 12299 17017 12311 17051
rect 14366 17048 14372 17060
rect 12253 17011 12311 17017
rect 13648 17020 14372 17048
rect 8665 16983 8723 16989
rect 8665 16980 8677 16983
rect 8128 16952 8677 16980
rect 8665 16949 8677 16952
rect 8711 16980 8723 16983
rect 11698 16980 11704 16992
rect 8711 16952 11704 16980
rect 8711 16949 8723 16952
rect 8665 16943 8723 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 12268 16980 12296 17011
rect 13648 16980 13676 17020
rect 14366 17008 14372 17020
rect 14424 17008 14430 17060
rect 15746 17048 15752 17060
rect 15580 17020 15752 17048
rect 12268 16952 13676 16980
rect 13722 16940 13728 16992
rect 13780 16980 13786 16992
rect 15580 16989 15608 17020
rect 15746 17008 15752 17020
rect 15804 17048 15810 17060
rect 17236 17057 17264 17088
rect 17589 17085 17601 17088
rect 17635 17085 17647 17119
rect 21358 17116 21364 17128
rect 21319 17088 21364 17116
rect 17589 17079 17647 17085
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 17221 17051 17279 17057
rect 17221 17048 17233 17051
rect 15804 17020 17233 17048
rect 15804 17008 15810 17020
rect 17221 17017 17233 17020
rect 17267 17017 17279 17051
rect 17221 17011 17279 17017
rect 18690 17008 18696 17060
rect 18748 17048 18754 17060
rect 19981 17051 20039 17057
rect 19981 17048 19993 17051
rect 18748 17020 19993 17048
rect 18748 17008 18754 17020
rect 19981 17017 19993 17020
rect 20027 17017 20039 17051
rect 19981 17011 20039 17017
rect 13909 16983 13967 16989
rect 13909 16980 13921 16983
rect 13780 16952 13921 16980
rect 13780 16940 13786 16952
rect 13909 16949 13921 16952
rect 13955 16980 13967 16983
rect 14277 16983 14335 16989
rect 14277 16980 14289 16983
rect 13955 16952 14289 16980
rect 13955 16949 13967 16952
rect 13909 16943 13967 16949
rect 14277 16949 14289 16952
rect 14323 16980 14335 16983
rect 14645 16983 14703 16989
rect 14645 16980 14657 16983
rect 14323 16952 14657 16980
rect 14323 16949 14335 16952
rect 14277 16943 14335 16949
rect 14645 16949 14657 16952
rect 14691 16980 14703 16983
rect 15565 16983 15623 16989
rect 15565 16980 15577 16983
rect 14691 16952 15577 16980
rect 14691 16949 14703 16952
rect 14645 16943 14703 16949
rect 15565 16949 15577 16952
rect 15611 16949 15623 16983
rect 15565 16943 15623 16949
rect 16945 16983 17003 16989
rect 16945 16949 16957 16983
rect 16991 16980 17003 16983
rect 18230 16980 18236 16992
rect 16991 16952 18236 16980
rect 16991 16949 17003 16952
rect 16945 16943 17003 16949
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 18966 16980 18972 16992
rect 18927 16952 18972 16980
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 19058 16940 19064 16992
rect 19116 16980 19122 16992
rect 19245 16983 19303 16989
rect 19245 16980 19257 16983
rect 19116 16952 19257 16980
rect 19116 16940 19122 16952
rect 19245 16949 19257 16952
rect 19291 16949 19303 16983
rect 19245 16943 19303 16949
rect 19518 16940 19524 16992
rect 19576 16980 19582 16992
rect 19613 16983 19671 16989
rect 19613 16980 19625 16983
rect 19576 16952 19625 16980
rect 19576 16940 19582 16952
rect 19613 16949 19625 16952
rect 19659 16949 19671 16983
rect 19613 16943 19671 16949
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 1946 16776 1952 16788
rect 1907 16748 1952 16776
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 3050 16736 3056 16788
rect 3108 16776 3114 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 3108 16748 3801 16776
rect 3108 16736 3114 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 4154 16776 4160 16788
rect 4115 16748 4160 16776
rect 3789 16739 3847 16745
rect 4154 16736 4160 16748
rect 4212 16736 4218 16788
rect 4706 16776 4712 16788
rect 4540 16748 4712 16776
rect 1581 16711 1639 16717
rect 1581 16677 1593 16711
rect 1627 16708 1639 16711
rect 3694 16708 3700 16720
rect 1627 16680 3700 16708
rect 1627 16677 1639 16680
rect 1581 16671 1639 16677
rect 3694 16668 3700 16680
rect 3752 16668 3758 16720
rect 2685 16643 2743 16649
rect 2685 16609 2697 16643
rect 2731 16640 2743 16643
rect 4540 16640 4568 16748
rect 4706 16736 4712 16748
rect 4764 16776 4770 16788
rect 5166 16776 5172 16788
rect 4764 16748 5172 16776
rect 4764 16736 4770 16748
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 6638 16736 6644 16788
rect 6696 16776 6702 16788
rect 8941 16779 8999 16785
rect 8941 16776 8953 16779
rect 6696 16748 8953 16776
rect 6696 16736 6702 16748
rect 8941 16745 8953 16748
rect 8987 16745 8999 16779
rect 13722 16776 13728 16788
rect 8941 16739 8999 16745
rect 12360 16748 13728 16776
rect 5994 16708 6000 16720
rect 4632 16680 6000 16708
rect 4632 16649 4660 16680
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 7098 16668 7104 16720
rect 7156 16708 7162 16720
rect 7156 16680 7880 16708
rect 7156 16668 7162 16680
rect 2731 16612 4568 16640
rect 4617 16643 4675 16649
rect 2731 16609 2743 16612
rect 2685 16603 2743 16609
rect 4617 16609 4629 16643
rect 4663 16609 4675 16643
rect 4617 16603 4675 16609
rect 4801 16643 4859 16649
rect 4801 16609 4813 16643
rect 4847 16640 4859 16643
rect 5074 16640 5080 16652
rect 4847 16612 5080 16640
rect 4847 16609 4859 16612
rect 4801 16603 4859 16609
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 7190 16640 7196 16652
rect 7151 16612 7196 16640
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16572 2191 16575
rect 2774 16572 2780 16584
rect 2179 16544 2780 16572
rect 2179 16541 2191 16544
rect 2133 16535 2191 16541
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 2866 16532 2872 16584
rect 2924 16572 2930 16584
rect 3145 16575 3203 16581
rect 3145 16572 3157 16575
rect 2924 16544 3157 16572
rect 2924 16532 2930 16544
rect 3145 16541 3157 16544
rect 3191 16541 3203 16575
rect 3145 16535 3203 16541
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16572 3479 16575
rect 5810 16572 5816 16584
rect 3467 16544 5304 16572
rect 5771 16544 5816 16572
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 4525 16507 4583 16513
rect 4525 16473 4537 16507
rect 4571 16504 4583 16507
rect 5169 16507 5227 16513
rect 5169 16504 5181 16507
rect 4571 16476 5181 16504
rect 4571 16473 4583 16476
rect 4525 16467 4583 16473
rect 5169 16473 5181 16476
rect 5215 16473 5227 16507
rect 5169 16467 5227 16473
rect 5276 16436 5304 16544
rect 5810 16532 5816 16544
rect 5868 16532 5874 16584
rect 6089 16575 6147 16581
rect 6089 16541 6101 16575
rect 6135 16572 6147 16575
rect 6546 16572 6552 16584
rect 6135 16544 6552 16572
rect 6135 16541 6147 16544
rect 6089 16535 6147 16541
rect 6546 16532 6552 16544
rect 6604 16532 6610 16584
rect 6549 16439 6607 16445
rect 6549 16436 6561 16439
rect 5276 16408 6561 16436
rect 6549 16405 6561 16408
rect 6595 16405 6607 16439
rect 6914 16436 6920 16448
rect 6875 16408 6920 16436
rect 6549 16399 6607 16405
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 7009 16439 7067 16445
rect 7009 16405 7021 16439
rect 7055 16436 7067 16439
rect 7558 16436 7564 16448
rect 7055 16408 7564 16436
rect 7055 16405 7067 16408
rect 7009 16399 7067 16405
rect 7558 16396 7564 16408
rect 7616 16396 7622 16448
rect 7852 16436 7880 16680
rect 8018 16640 8024 16652
rect 7979 16612 8024 16640
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 8386 16600 8392 16652
rect 8444 16640 8450 16652
rect 12360 16649 12388 16748
rect 13722 16736 13728 16748
rect 13780 16776 13786 16788
rect 13780 16748 13860 16776
rect 13780 16736 13786 16748
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 8444 16612 10977 16640
rect 8444 16600 8450 16612
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11149 16643 11207 16649
rect 11149 16609 11161 16643
rect 11195 16640 11207 16643
rect 12345 16643 12403 16649
rect 11195 16612 12296 16640
rect 11195 16609 11207 16612
rect 11149 16603 11207 16609
rect 8110 16532 8116 16584
rect 8168 16532 8174 16584
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 9769 16575 9827 16581
rect 9769 16572 9781 16575
rect 9732 16544 9781 16572
rect 9732 16532 9738 16544
rect 9769 16541 9781 16544
rect 9815 16541 9827 16575
rect 10042 16572 10048 16584
rect 10003 16544 10048 16572
rect 9769 16535 9827 16541
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 10870 16572 10876 16584
rect 10831 16544 10876 16572
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 12268 16572 12296 16612
rect 12345 16609 12357 16643
rect 12391 16609 12403 16643
rect 12345 16603 12403 16609
rect 13832 16584 13860 16748
rect 13998 16736 14004 16788
rect 14056 16776 14062 16788
rect 17770 16776 17776 16788
rect 14056 16748 17776 16776
rect 14056 16736 14062 16748
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 15470 16708 15476 16720
rect 15431 16680 15476 16708
rect 15470 16668 15476 16680
rect 15528 16668 15534 16720
rect 19058 16640 19064 16652
rect 18892 16612 19064 16640
rect 18892 16584 18920 16612
rect 19058 16600 19064 16612
rect 19116 16640 19122 16652
rect 19429 16643 19487 16649
rect 19429 16640 19441 16643
rect 19116 16612 19441 16640
rect 19116 16600 19122 16612
rect 19429 16609 19441 16612
rect 19475 16609 19487 16643
rect 19429 16603 19487 16609
rect 12268 16544 12434 16572
rect 8128 16504 8156 16532
rect 8128 16476 8616 16504
rect 8113 16439 8171 16445
rect 8113 16436 8125 16439
rect 7852 16408 8125 16436
rect 8113 16405 8125 16408
rect 8159 16405 8171 16439
rect 8113 16399 8171 16405
rect 8202 16396 8208 16448
rect 8260 16436 8266 16448
rect 8588 16445 8616 16476
rect 12406 16448 12434 16544
rect 13814 16532 13820 16584
rect 13872 16572 13878 16584
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 13872 16544 14105 16572
rect 13872 16532 13878 16544
rect 14093 16541 14105 16544
rect 14139 16572 14151 16575
rect 15749 16575 15807 16581
rect 15749 16572 15761 16575
rect 14139 16544 15761 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 15749 16541 15761 16544
rect 15795 16541 15807 16575
rect 18874 16572 18880 16584
rect 15749 16535 15807 16541
rect 15856 16544 17540 16572
rect 18835 16544 18880 16572
rect 12618 16513 12624 16516
rect 12612 16504 12624 16513
rect 12579 16476 12624 16504
rect 12612 16467 12624 16476
rect 12618 16464 12624 16467
rect 12676 16464 12682 16516
rect 13262 16464 13268 16516
rect 13320 16504 13326 16516
rect 14366 16513 14372 16516
rect 14360 16504 14372 16513
rect 13320 16476 14228 16504
rect 14327 16476 14372 16504
rect 13320 16464 13326 16476
rect 8573 16439 8631 16445
rect 8260 16408 8305 16436
rect 8260 16396 8266 16408
rect 8573 16405 8585 16439
rect 8619 16405 8631 16439
rect 8573 16399 8631 16405
rect 10226 16396 10232 16448
rect 10284 16436 10290 16448
rect 10505 16439 10563 16445
rect 10505 16436 10517 16439
rect 10284 16408 10517 16436
rect 10284 16396 10290 16408
rect 10505 16405 10517 16408
rect 10551 16405 10563 16439
rect 10505 16399 10563 16405
rect 11701 16439 11759 16445
rect 11701 16405 11713 16439
rect 11747 16436 11759 16439
rect 11882 16436 11888 16448
rect 11747 16408 11888 16436
rect 11747 16405 11759 16408
rect 11701 16399 11759 16405
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 12406 16408 12440 16448
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 13722 16436 13728 16448
rect 13683 16408 13728 16436
rect 13722 16396 13728 16408
rect 13780 16396 13786 16448
rect 14200 16436 14228 16476
rect 14360 16467 14372 16476
rect 14366 16464 14372 16467
rect 14424 16464 14430 16516
rect 14458 16464 14464 16516
rect 14516 16504 14522 16516
rect 15856 16504 15884 16544
rect 16016 16507 16074 16513
rect 16016 16504 16028 16507
rect 14516 16476 15884 16504
rect 15948 16476 16028 16504
rect 14516 16464 14522 16476
rect 15948 16436 15976 16476
rect 16016 16473 16028 16476
rect 16062 16473 16074 16507
rect 16016 16467 16074 16473
rect 17126 16436 17132 16448
rect 14200 16408 15976 16436
rect 17087 16408 17132 16436
rect 17126 16396 17132 16408
rect 17184 16396 17190 16448
rect 17512 16445 17540 16544
rect 18874 16532 18880 16544
rect 18932 16532 18938 16584
rect 19518 16532 19524 16584
rect 19576 16572 19582 16584
rect 19685 16575 19743 16581
rect 19685 16572 19697 16575
rect 19576 16544 19697 16572
rect 19576 16532 19582 16544
rect 19685 16541 19697 16544
rect 19731 16541 19743 16575
rect 19685 16535 19743 16541
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 20864 16544 21097 16572
rect 20864 16532 20870 16544
rect 21085 16541 21097 16544
rect 21131 16572 21143 16575
rect 21358 16572 21364 16584
rect 21131 16544 21364 16572
rect 21131 16541 21143 16544
rect 21085 16535 21143 16541
rect 21358 16532 21364 16544
rect 21416 16532 21422 16584
rect 18230 16464 18236 16516
rect 18288 16504 18294 16516
rect 18610 16507 18668 16513
rect 18610 16504 18622 16507
rect 18288 16476 18622 16504
rect 18288 16464 18294 16476
rect 18610 16473 18622 16476
rect 18656 16473 18668 16507
rect 18610 16467 18668 16473
rect 17497 16439 17555 16445
rect 17497 16405 17509 16439
rect 17543 16405 17555 16439
rect 17497 16399 17555 16405
rect 20622 16396 20628 16448
rect 20680 16436 20686 16448
rect 20809 16439 20867 16445
rect 20809 16436 20821 16439
rect 20680 16408 20821 16436
rect 20680 16396 20686 16408
rect 20809 16405 20821 16408
rect 20855 16405 20867 16439
rect 20809 16399 20867 16405
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 1949 16235 2007 16241
rect 1949 16201 1961 16235
rect 1995 16232 2007 16235
rect 2038 16232 2044 16244
rect 1995 16204 2044 16232
rect 1995 16201 2007 16204
rect 1949 16195 2007 16201
rect 2038 16192 2044 16204
rect 2096 16192 2102 16244
rect 3326 16232 3332 16244
rect 3287 16204 3332 16232
rect 3326 16192 3332 16204
rect 3384 16192 3390 16244
rect 3418 16192 3424 16244
rect 3476 16232 3482 16244
rect 3789 16235 3847 16241
rect 3789 16232 3801 16235
rect 3476 16204 3801 16232
rect 3476 16192 3482 16204
rect 3789 16201 3801 16204
rect 3835 16201 3847 16235
rect 3789 16195 3847 16201
rect 5350 16192 5356 16244
rect 5408 16232 5414 16244
rect 5537 16235 5595 16241
rect 5537 16232 5549 16235
rect 5408 16204 5549 16232
rect 5408 16192 5414 16204
rect 5537 16201 5549 16204
rect 5583 16201 5595 16235
rect 5537 16195 5595 16201
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6365 16235 6423 16241
rect 6365 16232 6377 16235
rect 6052 16204 6377 16232
rect 6052 16192 6058 16204
rect 6365 16201 6377 16204
rect 6411 16201 6423 16235
rect 6365 16195 6423 16201
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 7377 16235 7435 16241
rect 7377 16232 7389 16235
rect 6972 16204 7389 16232
rect 6972 16192 6978 16204
rect 7377 16201 7389 16204
rect 7423 16201 7435 16235
rect 7926 16232 7932 16244
rect 7887 16204 7932 16232
rect 7377 16195 7435 16201
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 8297 16235 8355 16241
rect 8297 16201 8309 16235
rect 8343 16232 8355 16235
rect 8570 16232 8576 16244
rect 8343 16204 8576 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 8570 16192 8576 16204
rect 8628 16232 8634 16244
rect 9033 16235 9091 16241
rect 9033 16232 9045 16235
rect 8628 16204 9045 16232
rect 8628 16192 8634 16204
rect 9033 16201 9045 16204
rect 9079 16232 9091 16235
rect 9306 16232 9312 16244
rect 9079 16204 9312 16232
rect 9079 16201 9091 16204
rect 9033 16195 9091 16201
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 11882 16232 11888 16244
rect 11843 16204 11888 16232
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 19518 16232 19524 16244
rect 13780 16204 19524 16232
rect 13780 16192 13786 16204
rect 19518 16192 19524 16204
rect 19576 16192 19582 16244
rect 2774 16124 2780 16176
rect 2832 16164 2838 16176
rect 3694 16164 3700 16176
rect 2832 16136 2877 16164
rect 3655 16136 3700 16164
rect 2832 16124 2838 16136
rect 3694 16124 3700 16136
rect 3752 16124 3758 16176
rect 4062 16124 4068 16176
rect 4120 16164 4126 16176
rect 4525 16167 4583 16173
rect 4525 16164 4537 16167
rect 4120 16136 4537 16164
rect 4120 16124 4126 16136
rect 4525 16133 4537 16136
rect 4571 16133 4583 16167
rect 4525 16127 4583 16133
rect 6733 16167 6791 16173
rect 6733 16133 6745 16167
rect 6779 16164 6791 16167
rect 6822 16164 6828 16176
rect 6779 16136 6828 16164
rect 6779 16133 6791 16136
rect 6733 16127 6791 16133
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 9674 16164 9680 16176
rect 7024 16136 9680 16164
rect 1486 16056 1492 16108
rect 1544 16096 1550 16108
rect 2133 16099 2191 16105
rect 2133 16096 2145 16099
rect 1544 16068 2145 16096
rect 1544 16056 1550 16068
rect 2133 16065 2145 16068
rect 2179 16065 2191 16099
rect 2133 16059 2191 16065
rect 3053 16099 3111 16105
rect 3053 16065 3065 16099
rect 3099 16096 3111 16099
rect 3326 16096 3332 16108
rect 3099 16068 3332 16096
rect 3099 16065 3111 16068
rect 3053 16059 3111 16065
rect 3326 16056 3332 16068
rect 3384 16056 3390 16108
rect 3712 16096 3740 16124
rect 4801 16099 4859 16105
rect 3712 16068 4108 16096
rect 4080 16040 4108 16068
rect 4801 16065 4813 16099
rect 4847 16065 4859 16099
rect 4801 16059 4859 16065
rect 3142 15988 3148 16040
rect 3200 16028 3206 16040
rect 3881 16031 3939 16037
rect 3881 16028 3893 16031
rect 3200 16000 3893 16028
rect 3200 15988 3206 16000
rect 3881 15997 3893 16000
rect 3927 15997 3939 16031
rect 3881 15991 3939 15997
rect 4062 15988 4068 16040
rect 4120 15988 4126 16040
rect 4816 15960 4844 16059
rect 5166 16056 5172 16108
rect 5224 16096 5230 16108
rect 5445 16099 5503 16105
rect 5445 16096 5457 16099
rect 5224 16068 5457 16096
rect 5224 16056 5230 16068
rect 5445 16065 5457 16068
rect 5491 16065 5503 16099
rect 5445 16059 5503 16065
rect 5721 16031 5779 16037
rect 5721 15997 5733 16031
rect 5767 16028 5779 16031
rect 6270 16028 6276 16040
rect 5767 16000 6276 16028
rect 5767 15997 5779 16000
rect 5721 15991 5779 15997
rect 6270 15988 6276 16000
rect 6328 15988 6334 16040
rect 6638 15988 6644 16040
rect 6696 16028 6702 16040
rect 7024 16037 7052 16136
rect 9674 16124 9680 16136
rect 9732 16124 9738 16176
rect 9858 16124 9864 16176
rect 9916 16164 9922 16176
rect 9953 16167 10011 16173
rect 9953 16164 9965 16167
rect 9916 16136 9965 16164
rect 9916 16124 9922 16136
rect 9953 16133 9965 16136
rect 9999 16133 10011 16167
rect 9953 16127 10011 16133
rect 10686 16124 10692 16176
rect 10744 16164 10750 16176
rect 10781 16167 10839 16173
rect 10781 16164 10793 16167
rect 10744 16136 10793 16164
rect 10744 16124 10750 16136
rect 10781 16133 10793 16136
rect 10827 16133 10839 16167
rect 10781 16127 10839 16133
rect 13814 16124 13820 16176
rect 13872 16164 13878 16176
rect 15197 16167 15255 16173
rect 15197 16164 15209 16167
rect 13872 16136 15209 16164
rect 13872 16124 13878 16136
rect 8389 16099 8447 16105
rect 8389 16065 8401 16099
rect 8435 16096 8447 16099
rect 9030 16096 9036 16108
rect 8435 16068 9036 16096
rect 8435 16065 8447 16068
rect 8389 16059 8447 16065
rect 9030 16056 9036 16068
rect 9088 16096 9094 16108
rect 9309 16099 9367 16105
rect 9309 16096 9321 16099
rect 9088 16068 9321 16096
rect 9088 16056 9094 16068
rect 9309 16065 9321 16068
rect 9355 16065 9367 16099
rect 10226 16096 10232 16108
rect 10187 16068 10232 16096
rect 9309 16059 9367 16065
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 10502 16096 10508 16108
rect 10463 16068 10508 16096
rect 10502 16056 10508 16068
rect 10560 16056 10566 16108
rect 13998 16096 14004 16108
rect 12176 16068 14004 16096
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6696 16000 6837 16028
rect 6696 15988 6702 16000
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 7009 16031 7067 16037
rect 7009 15997 7021 16031
rect 7055 15997 7067 16031
rect 7009 15991 7067 15997
rect 8481 16031 8539 16037
rect 8481 15997 8493 16031
rect 8527 15997 8539 16031
rect 11330 16028 11336 16040
rect 8481 15991 8539 15997
rect 8772 16000 11336 16028
rect 5994 15960 6000 15972
rect 4816 15932 6000 15960
rect 5994 15920 6000 15932
rect 6052 15920 6058 15972
rect 7190 15920 7196 15972
rect 7248 15960 7254 15972
rect 8496 15960 8524 15991
rect 8772 15960 8800 16000
rect 11330 15988 11336 16000
rect 11388 15988 11394 16040
rect 12176 16037 12204 16068
rect 13998 16056 14004 16068
rect 14056 16056 14062 16108
rect 14568 16105 14596 16136
rect 15197 16133 15209 16136
rect 15243 16133 15255 16167
rect 15197 16127 15255 16133
rect 16482 16124 16488 16176
rect 16540 16164 16546 16176
rect 17782 16167 17840 16173
rect 17782 16164 17794 16167
rect 16540 16136 17794 16164
rect 16540 16124 16546 16136
rect 17782 16133 17794 16136
rect 17828 16164 17840 16167
rect 18690 16164 18696 16176
rect 17828 16136 18696 16164
rect 17828 16133 17840 16136
rect 17782 16127 17840 16133
rect 18690 16124 18696 16136
rect 18748 16124 18754 16176
rect 18966 16124 18972 16176
rect 19024 16164 19030 16176
rect 19306 16167 19364 16173
rect 19306 16164 19318 16167
rect 19024 16136 19318 16164
rect 19024 16124 19030 16136
rect 19306 16133 19318 16136
rect 19352 16133 19364 16167
rect 19306 16127 19364 16133
rect 14297 16099 14355 16105
rect 14297 16065 14309 16099
rect 14343 16096 14355 16099
rect 14553 16099 14611 16105
rect 14343 16068 14504 16096
rect 14343 16065 14355 16068
rect 14297 16059 14355 16065
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 12161 16031 12219 16037
rect 12161 15997 12173 16031
rect 12207 15997 12219 16031
rect 14476 16028 14504 16068
rect 14553 16065 14565 16099
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18322 16096 18328 16108
rect 18095 16068 18328 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 18322 16056 18328 16068
rect 18380 16096 18386 16108
rect 18874 16096 18880 16108
rect 18380 16068 18880 16096
rect 18380 16056 18386 16068
rect 18874 16056 18880 16068
rect 18932 16096 18938 16108
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 18932 16068 19073 16096
rect 18932 16056 18938 16068
rect 19061 16065 19073 16068
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 14476 16000 14596 16028
rect 12161 15991 12219 15997
rect 11992 15960 12020 15991
rect 7248 15932 8800 15960
rect 9646 15932 12020 15960
rect 14568 15960 14596 16000
rect 14568 15932 15148 15960
rect 7248 15920 7254 15932
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 3050 15892 3056 15904
rect 1627 15864 3056 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5077 15895 5135 15901
rect 5077 15892 5089 15895
rect 5040 15864 5089 15892
rect 5040 15852 5046 15864
rect 5077 15861 5089 15864
rect 5123 15861 5135 15895
rect 5077 15855 5135 15861
rect 7374 15852 7380 15904
rect 7432 15892 7438 15904
rect 9646 15892 9674 15932
rect 15120 15904 15148 15932
rect 15378 15920 15384 15972
rect 15436 15960 15442 15972
rect 16482 15960 16488 15972
rect 15436 15932 16488 15960
rect 15436 15920 15442 15932
rect 16482 15920 16488 15932
rect 16540 15920 16546 15972
rect 21082 15920 21088 15972
rect 21140 15960 21146 15972
rect 21177 15963 21235 15969
rect 21177 15960 21189 15963
rect 21140 15932 21189 15960
rect 21140 15920 21146 15932
rect 21177 15929 21189 15932
rect 21223 15929 21235 15963
rect 21177 15923 21235 15929
rect 7432 15864 9674 15892
rect 7432 15852 7438 15864
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 10560 15864 11529 15892
rect 10560 15852 10566 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11517 15855 11575 15861
rect 13173 15895 13231 15901
rect 13173 15861 13185 15895
rect 13219 15892 13231 15895
rect 13262 15892 13268 15904
rect 13219 15864 13268 15892
rect 13219 15861 13231 15864
rect 13173 15855 13231 15861
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 14918 15852 14924 15904
rect 14976 15892 14982 15904
rect 14976 15864 15021 15892
rect 14976 15852 14982 15864
rect 15102 15852 15108 15904
rect 15160 15892 15166 15904
rect 15565 15895 15623 15901
rect 15565 15892 15577 15895
rect 15160 15864 15577 15892
rect 15160 15852 15166 15864
rect 15565 15861 15577 15864
rect 15611 15861 15623 15895
rect 15565 15855 15623 15861
rect 16669 15895 16727 15901
rect 16669 15861 16681 15895
rect 16715 15892 16727 15895
rect 16942 15892 16948 15904
rect 16715 15864 16948 15892
rect 16715 15861 16727 15864
rect 16669 15855 16727 15861
rect 16942 15852 16948 15864
rect 17000 15852 17006 15904
rect 18322 15892 18328 15904
rect 18283 15864 18328 15892
rect 18322 15852 18328 15864
rect 18380 15852 18386 15904
rect 20438 15892 20444 15904
rect 20399 15864 20444 15892
rect 20438 15852 20444 15864
rect 20496 15852 20502 15904
rect 20806 15892 20812 15904
rect 20767 15864 20812 15892
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 1949 15691 2007 15697
rect 1949 15688 1961 15691
rect 1912 15660 1961 15688
rect 1912 15648 1918 15660
rect 1949 15657 1961 15660
rect 1995 15657 2007 15691
rect 1949 15651 2007 15657
rect 2406 15648 2412 15700
rect 2464 15688 2470 15700
rect 2501 15691 2559 15697
rect 2501 15688 2513 15691
rect 2464 15660 2513 15688
rect 2464 15648 2470 15660
rect 2501 15657 2513 15660
rect 2547 15657 2559 15691
rect 2501 15651 2559 15657
rect 2958 15648 2964 15700
rect 3016 15688 3022 15700
rect 3142 15688 3148 15700
rect 3016 15660 3148 15688
rect 3016 15648 3022 15660
rect 3142 15648 3148 15660
rect 3200 15688 3206 15700
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 3200 15660 3341 15688
rect 3200 15648 3206 15660
rect 3329 15657 3341 15660
rect 3375 15657 3387 15691
rect 3329 15651 3387 15657
rect 4341 15691 4399 15697
rect 4341 15657 4353 15691
rect 4387 15688 4399 15691
rect 6730 15688 6736 15700
rect 4387 15660 6736 15688
rect 4387 15657 4399 15660
rect 4341 15651 4399 15657
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 7374 15688 7380 15700
rect 7335 15660 7380 15688
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 8573 15691 8631 15697
rect 8573 15657 8585 15691
rect 8619 15688 8631 15691
rect 9398 15688 9404 15700
rect 8619 15660 9404 15688
rect 8619 15657 8631 15660
rect 8573 15651 8631 15657
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 13722 15688 13728 15700
rect 9548 15660 13728 15688
rect 9548 15648 9554 15660
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 14090 15648 14096 15700
rect 14148 15688 14154 15700
rect 15473 15691 15531 15697
rect 15473 15688 15485 15691
rect 14148 15660 15485 15688
rect 14148 15648 14154 15660
rect 15473 15657 15485 15660
rect 15519 15688 15531 15691
rect 15838 15688 15844 15700
rect 15519 15660 15844 15688
rect 15519 15657 15531 15660
rect 15473 15651 15531 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 1581 15623 1639 15629
rect 1581 15589 1593 15623
rect 1627 15620 1639 15623
rect 3418 15620 3424 15632
rect 1627 15592 3424 15620
rect 1627 15589 1639 15592
rect 1581 15583 1639 15589
rect 3418 15580 3424 15592
rect 3476 15580 3482 15632
rect 3973 15623 4031 15629
rect 3973 15589 3985 15623
rect 4019 15620 4031 15623
rect 5353 15623 5411 15629
rect 4019 15592 5304 15620
rect 4019 15589 4031 15592
rect 3973 15583 4031 15589
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 5074 15552 5080 15564
rect 4847 15524 5080 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 2130 15484 2136 15496
rect 2091 15456 2136 15484
rect 2130 15444 2136 15456
rect 2188 15444 2194 15496
rect 2682 15484 2688 15496
rect 2643 15456 2688 15484
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 4982 15484 4988 15496
rect 4943 15456 4988 15484
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 5276 15484 5304 15592
rect 5353 15589 5365 15623
rect 5399 15620 5411 15623
rect 7098 15620 7104 15632
rect 5399 15592 7104 15620
rect 5399 15589 5411 15592
rect 5353 15583 5411 15589
rect 7098 15580 7104 15592
rect 7156 15580 7162 15632
rect 7944 15592 8248 15620
rect 6270 15552 6276 15564
rect 6231 15524 6276 15552
rect 6270 15512 6276 15524
rect 6328 15512 6334 15564
rect 6825 15555 6883 15561
rect 6825 15521 6837 15555
rect 6871 15552 6883 15555
rect 7944 15552 7972 15592
rect 6871 15524 7972 15552
rect 6871 15521 6883 15524
rect 6825 15515 6883 15521
rect 8018 15512 8024 15564
rect 8076 15552 8082 15564
rect 8220 15552 8248 15592
rect 8662 15580 8668 15632
rect 8720 15620 8726 15632
rect 13446 15620 13452 15632
rect 8720 15592 13452 15620
rect 8720 15580 8726 15592
rect 13446 15580 13452 15592
rect 13504 15580 13510 15632
rect 11425 15555 11483 15561
rect 8076 15524 8121 15552
rect 8220 15524 8340 15552
rect 8076 15512 8082 15524
rect 5718 15484 5724 15496
rect 5276 15456 5724 15484
rect 5718 15444 5724 15456
rect 5776 15484 5782 15496
rect 5997 15487 6055 15493
rect 5997 15484 6009 15487
rect 5776 15456 6009 15484
rect 5776 15444 5782 15456
rect 5997 15453 6009 15456
rect 6043 15453 6055 15487
rect 6917 15487 6975 15493
rect 6917 15484 6929 15487
rect 5997 15447 6055 15453
rect 6104 15456 6929 15484
rect 3053 15419 3111 15425
rect 3053 15385 3065 15419
rect 3099 15416 3111 15419
rect 3418 15416 3424 15428
rect 3099 15388 3424 15416
rect 3099 15385 3111 15388
rect 3053 15379 3111 15385
rect 3418 15376 3424 15388
rect 3476 15376 3482 15428
rect 4893 15419 4951 15425
rect 4893 15385 4905 15419
rect 4939 15385 4951 15419
rect 4893 15379 4951 15385
rect 4908 15348 4936 15379
rect 5350 15376 5356 15428
rect 5408 15416 5414 15428
rect 6104 15416 6132 15456
rect 6917 15453 6929 15456
rect 6963 15453 6975 15487
rect 6917 15447 6975 15453
rect 8202 15444 8208 15496
rect 8260 15444 8266 15496
rect 6638 15416 6644 15428
rect 5408 15388 6132 15416
rect 6196 15388 6644 15416
rect 5408 15376 5414 15388
rect 5736 15360 5764 15388
rect 5629 15351 5687 15357
rect 5629 15348 5641 15351
rect 4908 15320 5641 15348
rect 5629 15317 5641 15320
rect 5675 15317 5687 15351
rect 5629 15311 5687 15317
rect 5718 15308 5724 15360
rect 5776 15308 5782 15360
rect 6089 15351 6147 15357
rect 6089 15317 6101 15351
rect 6135 15348 6147 15351
rect 6196 15348 6224 15388
rect 6638 15376 6644 15388
rect 6696 15376 6702 15428
rect 6730 15376 6736 15428
rect 6788 15416 6794 15428
rect 7009 15419 7067 15425
rect 7009 15416 7021 15419
rect 6788 15388 7021 15416
rect 6788 15376 6794 15388
rect 7009 15385 7021 15388
rect 7055 15385 7067 15419
rect 7009 15379 7067 15385
rect 7374 15376 7380 15428
rect 7432 15416 7438 15428
rect 8220 15416 8248 15444
rect 7432 15388 8248 15416
rect 8312 15416 8340 15524
rect 9048 15524 10640 15552
rect 8478 15444 8484 15496
rect 8536 15484 8542 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8536 15456 8953 15484
rect 8536 15444 8542 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9048 15416 9076 15524
rect 9582 15444 9588 15496
rect 9640 15484 9646 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 9640 15456 10241 15484
rect 9640 15444 9646 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 10502 15484 10508 15496
rect 10463 15456 10508 15484
rect 10229 15447 10287 15453
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 10612 15484 10640 15524
rect 11425 15521 11437 15555
rect 11471 15552 11483 15555
rect 11471 15524 13676 15552
rect 11471 15521 11483 15524
rect 11425 15515 11483 15521
rect 13538 15484 13544 15496
rect 10612 15456 13544 15484
rect 13538 15444 13544 15456
rect 13596 15444 13602 15496
rect 8312 15388 9076 15416
rect 11149 15419 11207 15425
rect 7432 15376 7438 15388
rect 11149 15385 11161 15419
rect 11195 15416 11207 15419
rect 11793 15419 11851 15425
rect 11793 15416 11805 15419
rect 11195 15388 11805 15416
rect 11195 15385 11207 15388
rect 11149 15379 11207 15385
rect 11793 15385 11805 15388
rect 11839 15385 11851 15419
rect 13648 15416 13676 15524
rect 13814 15444 13820 15496
rect 13872 15484 13878 15496
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13872 15456 14105 15484
rect 13872 15444 13878 15456
rect 14093 15453 14105 15456
rect 14139 15484 14151 15487
rect 15749 15487 15807 15493
rect 15749 15484 15761 15487
rect 14139 15456 15761 15484
rect 14139 15453 14151 15456
rect 14093 15447 14151 15453
rect 15749 15453 15761 15456
rect 15795 15484 15807 15487
rect 16761 15487 16819 15493
rect 16761 15484 16773 15487
rect 15795 15456 16773 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 16761 15453 16773 15456
rect 16807 15484 16819 15487
rect 18322 15484 18328 15496
rect 16807 15456 18328 15484
rect 16807 15453 16819 15456
rect 16761 15447 16819 15453
rect 18322 15444 18328 15456
rect 18380 15484 18386 15496
rect 18417 15487 18475 15493
rect 18417 15484 18429 15487
rect 18380 15456 18429 15484
rect 18380 15444 18386 15456
rect 18417 15453 18429 15456
rect 18463 15484 18475 15487
rect 18785 15487 18843 15493
rect 18785 15484 18797 15487
rect 18463 15456 18797 15484
rect 18463 15453 18475 15456
rect 18417 15447 18475 15453
rect 18785 15453 18797 15456
rect 18831 15453 18843 15487
rect 19610 15484 19616 15496
rect 19571 15456 19616 15484
rect 18785 15447 18843 15453
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 20806 15444 20812 15496
rect 20864 15484 20870 15496
rect 21361 15487 21419 15493
rect 21361 15484 21373 15487
rect 20864 15456 21373 15484
rect 20864 15444 20870 15456
rect 21361 15453 21373 15456
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 14360 15419 14418 15425
rect 13648 15388 14320 15416
rect 11793 15379 11851 15385
rect 6135 15320 6224 15348
rect 6135 15317 6147 15320
rect 6089 15311 6147 15317
rect 6270 15308 6276 15360
rect 6328 15348 6334 15360
rect 6914 15348 6920 15360
rect 6328 15320 6920 15348
rect 6328 15308 6334 15320
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 7558 15308 7564 15360
rect 7616 15348 7622 15360
rect 7926 15348 7932 15360
rect 7616 15320 7932 15348
rect 7616 15308 7622 15320
rect 7926 15308 7932 15320
rect 7984 15308 7990 15360
rect 8110 15348 8116 15360
rect 8071 15320 8116 15348
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 8205 15351 8263 15357
rect 8205 15317 8217 15351
rect 8251 15348 8263 15351
rect 8662 15348 8668 15360
rect 8251 15320 8668 15348
rect 8251 15317 8263 15320
rect 8205 15311 8263 15317
rect 8662 15308 8668 15320
rect 8720 15308 8726 15360
rect 10778 15348 10784 15360
rect 10739 15320 10784 15348
rect 10778 15308 10784 15320
rect 10836 15308 10842 15360
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 11241 15351 11299 15357
rect 11241 15348 11253 15351
rect 10928 15320 11253 15348
rect 10928 15308 10934 15320
rect 11241 15317 11253 15320
rect 11287 15317 11299 15351
rect 11241 15311 11299 15317
rect 11330 15308 11336 15360
rect 11388 15348 11394 15360
rect 14090 15348 14096 15360
rect 11388 15320 14096 15348
rect 11388 15308 11394 15320
rect 14090 15308 14096 15320
rect 14148 15308 14154 15360
rect 14292 15348 14320 15388
rect 14360 15385 14372 15419
rect 14406 15416 14418 15419
rect 14458 15416 14464 15428
rect 14406 15388 14464 15416
rect 14406 15385 14418 15388
rect 14360 15379 14418 15385
rect 14458 15376 14464 15388
rect 14516 15376 14522 15428
rect 17034 15425 17040 15428
rect 17028 15379 17040 15425
rect 17092 15416 17098 15428
rect 19628 15416 19656 15444
rect 20622 15416 20628 15428
rect 17092 15388 17128 15416
rect 19628 15388 20628 15416
rect 17034 15376 17040 15379
rect 17092 15376 17098 15388
rect 20622 15376 20628 15388
rect 20680 15416 20686 15428
rect 21094 15419 21152 15425
rect 21094 15416 21106 15419
rect 20680 15388 21106 15416
rect 20680 15376 20686 15388
rect 21094 15385 21106 15388
rect 21140 15385 21152 15419
rect 21094 15379 21152 15385
rect 16114 15348 16120 15360
rect 14292 15320 16120 15348
rect 16114 15308 16120 15320
rect 16172 15308 16178 15360
rect 16390 15348 16396 15360
rect 16351 15320 16396 15348
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 18138 15348 18144 15360
rect 18099 15320 18144 15348
rect 18138 15308 18144 15320
rect 18196 15308 18202 15360
rect 18966 15308 18972 15360
rect 19024 15348 19030 15360
rect 19337 15351 19395 15357
rect 19337 15348 19349 15351
rect 19024 15320 19349 15348
rect 19024 15308 19030 15320
rect 19337 15317 19349 15320
rect 19383 15317 19395 15351
rect 19337 15311 19395 15317
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 19981 15351 20039 15357
rect 19981 15348 19993 15351
rect 19852 15320 19993 15348
rect 19852 15308 19858 15320
rect 19981 15317 19993 15320
rect 20027 15317 20039 15351
rect 19981 15311 20039 15317
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 2777 15147 2835 15153
rect 2777 15113 2789 15147
rect 2823 15144 2835 15147
rect 2866 15144 2872 15156
rect 2823 15116 2872 15144
rect 2823 15113 2835 15116
rect 2777 15107 2835 15113
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 3973 15147 4031 15153
rect 3973 15113 3985 15147
rect 4019 15144 4031 15147
rect 5537 15147 5595 15153
rect 5537 15144 5549 15147
rect 4019 15116 5549 15144
rect 4019 15113 4031 15116
rect 3973 15107 4031 15113
rect 5537 15113 5549 15116
rect 5583 15113 5595 15147
rect 5537 15107 5595 15113
rect 5810 15104 5816 15156
rect 5868 15144 5874 15156
rect 5997 15147 6055 15153
rect 5997 15144 6009 15147
rect 5868 15116 6009 15144
rect 5868 15104 5874 15116
rect 5997 15113 6009 15116
rect 6043 15113 6055 15147
rect 5997 15107 6055 15113
rect 7561 15147 7619 15153
rect 7561 15113 7573 15147
rect 7607 15113 7619 15147
rect 7561 15107 7619 15113
rect 7837 15147 7895 15153
rect 7837 15113 7849 15147
rect 7883 15144 7895 15147
rect 8018 15144 8024 15156
rect 7883 15116 8024 15144
rect 7883 15113 7895 15116
rect 7837 15107 7895 15113
rect 2041 15079 2099 15085
rect 2041 15045 2053 15079
rect 2087 15076 2099 15079
rect 2130 15076 2136 15088
rect 2087 15048 2136 15076
rect 2087 15045 2099 15048
rect 2041 15039 2099 15045
rect 2130 15036 2136 15048
rect 2188 15036 2194 15088
rect 3418 15036 3424 15088
rect 3476 15076 3482 15088
rect 4617 15079 4675 15085
rect 4617 15076 4629 15079
rect 3476 15048 4629 15076
rect 3476 15036 3482 15048
rect 4617 15045 4629 15048
rect 4663 15045 4675 15079
rect 7098 15076 7104 15088
rect 7059 15048 7104 15076
rect 4617 15039 4675 15045
rect 7098 15036 7104 15048
rect 7156 15036 7162 15088
rect 7208 15048 7512 15076
rect 2314 15008 2320 15020
rect 2275 14980 2320 15008
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 2590 15008 2596 15020
rect 2551 14980 2596 15008
rect 2590 14968 2596 14980
rect 2648 14968 2654 15020
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 15008 3663 15011
rect 3878 15008 3884 15020
rect 3651 14980 3884 15008
rect 3651 14977 3663 14980
rect 3605 14971 3663 14977
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 5626 15008 5632 15020
rect 4571 14980 4660 15008
rect 5587 14980 5632 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14940 1639 14943
rect 3326 14940 3332 14952
rect 1627 14912 3332 14940
rect 1627 14909 1639 14912
rect 1581 14903 1639 14909
rect 3326 14900 3332 14912
rect 3384 14900 3390 14952
rect 3513 14943 3571 14949
rect 3513 14909 3525 14943
rect 3559 14940 3571 14943
rect 3970 14940 3976 14952
rect 3559 14912 3976 14940
rect 3559 14909 3571 14912
rect 3513 14903 3571 14909
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 4430 14940 4436 14952
rect 4391 14912 4436 14940
rect 4430 14900 4436 14912
rect 4488 14900 4494 14952
rect 4632 14884 4660 14980
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 7208 15017 7236 15048
rect 7193 15011 7251 15017
rect 7193 14977 7205 15011
rect 7239 14977 7251 15011
rect 7193 14971 7251 14977
rect 5445 14943 5503 14949
rect 5445 14909 5457 14943
rect 5491 14940 5503 14943
rect 6086 14940 6092 14952
rect 5491 14912 6092 14940
rect 5491 14909 5503 14912
rect 5445 14903 5503 14909
rect 6086 14900 6092 14912
rect 6144 14900 6150 14952
rect 7006 14940 7012 14952
rect 6967 14912 7012 14940
rect 7006 14900 7012 14912
rect 7064 14900 7070 14952
rect 4614 14832 4620 14884
rect 4672 14832 4678 14884
rect 6638 14872 6644 14884
rect 4816 14844 6644 14872
rect 2314 14764 2320 14816
rect 2372 14804 2378 14816
rect 4816 14804 4844 14844
rect 6638 14832 6644 14844
rect 6696 14832 6702 14884
rect 4982 14804 4988 14816
rect 2372 14776 4844 14804
rect 4943 14776 4988 14804
rect 2372 14764 2378 14776
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 5718 14764 5724 14816
rect 5776 14804 5782 14816
rect 6457 14807 6515 14813
rect 6457 14804 6469 14807
rect 5776 14776 6469 14804
rect 5776 14764 5782 14776
rect 6457 14773 6469 14776
rect 6503 14804 6515 14807
rect 6730 14804 6736 14816
rect 6503 14776 6736 14804
rect 6503 14773 6515 14776
rect 6457 14767 6515 14773
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 7484 14804 7512 15048
rect 7576 15020 7604 15107
rect 8018 15104 8024 15116
rect 8076 15104 8082 15156
rect 8386 15104 8392 15156
rect 8444 15144 8450 15156
rect 14458 15144 14464 15156
rect 8444 15116 14464 15144
rect 8444 15104 8450 15116
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 8297 15079 8355 15085
rect 8297 15045 8309 15079
rect 8343 15076 8355 15079
rect 8478 15076 8484 15088
rect 8343 15048 8484 15076
rect 8343 15045 8355 15048
rect 8297 15039 8355 15045
rect 8478 15036 8484 15048
rect 8536 15036 8542 15088
rect 9950 15036 9956 15088
rect 10008 15076 10014 15088
rect 10505 15079 10563 15085
rect 10505 15076 10517 15079
rect 10008 15048 10517 15076
rect 10008 15036 10014 15048
rect 10505 15045 10517 15048
rect 10551 15045 10563 15079
rect 10505 15039 10563 15045
rect 11793 15079 11851 15085
rect 11793 15045 11805 15079
rect 11839 15076 11851 15079
rect 11974 15076 11980 15088
rect 11839 15048 11980 15076
rect 11839 15045 11851 15048
rect 11793 15039 11851 15045
rect 11974 15036 11980 15048
rect 12032 15036 12038 15088
rect 13722 15076 13728 15088
rect 13188 15048 13728 15076
rect 7558 14968 7564 15020
rect 7616 14968 7622 15020
rect 8018 14968 8024 15020
rect 8076 15008 8082 15020
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 8076 14980 8217 15008
rect 8076 14968 8082 14980
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 8205 14971 8263 14977
rect 9217 15011 9275 15017
rect 9217 14977 9229 15011
rect 9263 15008 9275 15011
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 9263 14980 9873 15008
rect 9263 14977 9275 14980
rect 9217 14971 9275 14977
rect 9861 14977 9873 14980
rect 9907 14977 9919 15011
rect 10778 15008 10784 15020
rect 10739 14980 10784 15008
rect 9861 14971 9919 14977
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 11514 15008 11520 15020
rect 11475 14980 11520 15008
rect 11514 14968 11520 14980
rect 11572 14968 11578 15020
rect 11698 14968 11704 15020
rect 11756 15008 11762 15020
rect 13188 15017 13216 15048
rect 13722 15036 13728 15048
rect 13780 15036 13786 15088
rect 14274 15036 14280 15088
rect 14332 15076 14338 15088
rect 16056 15079 16114 15085
rect 14332 15048 15976 15076
rect 14332 15036 14338 15048
rect 13173 15011 13231 15017
rect 11756 14980 13124 15008
rect 11756 14968 11762 14980
rect 8389 14943 8447 14949
rect 8389 14909 8401 14943
rect 8435 14909 8447 14943
rect 9306 14940 9312 14952
rect 9267 14912 9312 14940
rect 8389 14903 8447 14909
rect 8202 14832 8208 14884
rect 8260 14872 8266 14884
rect 8404 14872 8432 14903
rect 9306 14900 9312 14912
rect 9364 14900 9370 14952
rect 9493 14943 9551 14949
rect 9493 14909 9505 14943
rect 9539 14909 9551 14943
rect 12986 14940 12992 14952
rect 9493 14903 9551 14909
rect 12406 14912 12992 14940
rect 8846 14872 8852 14884
rect 8260 14844 8432 14872
rect 8807 14844 8852 14872
rect 8260 14832 8266 14844
rect 8846 14832 8852 14844
rect 8904 14832 8910 14884
rect 9508 14872 9536 14903
rect 12406 14872 12434 14912
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 13096 14940 13124 14980
rect 13173 14977 13185 15011
rect 13219 14977 13231 15011
rect 13440 15011 13498 15017
rect 13440 15008 13452 15011
rect 13173 14971 13231 14977
rect 13280 14980 13452 15008
rect 13280 14940 13308 14980
rect 13440 14977 13452 14980
rect 13486 15008 13498 15011
rect 14918 15008 14924 15020
rect 13486 14980 14924 15008
rect 13486 14977 13498 14980
rect 13440 14971 13498 14977
rect 14918 14968 14924 14980
rect 14976 14968 14982 15020
rect 15948 15008 15976 15048
rect 16056 15045 16068 15079
rect 16102 15076 16114 15079
rect 16390 15076 16396 15088
rect 16102 15048 16396 15076
rect 16102 15045 16114 15048
rect 16056 15039 16114 15045
rect 16390 15036 16396 15048
rect 16448 15036 16454 15088
rect 17144 15048 18276 15076
rect 16301 15011 16359 15017
rect 15948 14980 16252 15008
rect 13096 14912 13308 14940
rect 16224 14940 16252 14980
rect 16301 14977 16313 15011
rect 16347 15008 16359 15011
rect 17144 15008 17172 15048
rect 17954 15008 17960 15020
rect 18012 15017 18018 15020
rect 18248 15017 18276 15048
rect 20806 15036 20812 15088
rect 20864 15076 20870 15088
rect 20864 15048 21404 15076
rect 20864 15036 20870 15048
rect 16347 14980 17172 15008
rect 17924 14980 17960 15008
rect 16347 14977 16359 14980
rect 16301 14971 16359 14977
rect 17954 14968 17960 14980
rect 18012 14971 18024 15017
rect 18233 15011 18291 15017
rect 18233 14977 18245 15011
rect 18279 15008 18291 15011
rect 18322 15008 18328 15020
rect 18279 14980 18328 15008
rect 18279 14977 18291 14980
rect 18233 14971 18291 14977
rect 18012 14968 18018 14971
rect 18322 14968 18328 14980
rect 18380 15008 18386 15020
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 18380 14980 18889 15008
rect 18380 14968 18386 14980
rect 18877 14977 18889 14980
rect 18923 15008 18935 15011
rect 19613 15011 19671 15017
rect 19613 15008 19625 15011
rect 18923 14980 19625 15008
rect 18923 14977 18935 14980
rect 18877 14971 18935 14977
rect 19613 14977 19625 14980
rect 19659 14977 19671 15011
rect 19613 14971 19671 14977
rect 19702 14968 19708 15020
rect 19760 15008 19766 15020
rect 21376 15017 21404 15048
rect 21094 15011 21152 15017
rect 21094 15008 21106 15011
rect 19760 14980 21106 15008
rect 19760 14968 19766 14980
rect 21094 14977 21106 14980
rect 21140 14977 21152 15011
rect 21094 14971 21152 14977
rect 21361 15011 21419 15017
rect 21361 14977 21373 15011
rect 21407 14977 21419 15011
rect 21361 14971 21419 14977
rect 16574 14940 16580 14952
rect 16224 14912 16580 14940
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 9508 14844 12434 14872
rect 14458 14832 14464 14884
rect 14516 14872 14522 14884
rect 14516 14844 15056 14872
rect 14516 14832 14522 14844
rect 7156 14776 7512 14804
rect 7156 14764 7162 14776
rect 10686 14764 10692 14816
rect 10744 14804 10750 14816
rect 12802 14804 12808 14816
rect 10744 14776 12808 14804
rect 10744 14764 10750 14776
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 14274 14764 14280 14816
rect 14332 14804 14338 14816
rect 14553 14807 14611 14813
rect 14553 14804 14565 14807
rect 14332 14776 14565 14804
rect 14332 14764 14338 14776
rect 14553 14773 14565 14776
rect 14599 14773 14611 14807
rect 14553 14767 14611 14773
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 14921 14807 14979 14813
rect 14921 14804 14933 14807
rect 14792 14776 14933 14804
rect 14792 14764 14798 14776
rect 14921 14773 14933 14776
rect 14967 14773 14979 14807
rect 15028 14804 15056 14844
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 15028 14776 16865 14804
rect 14921 14767 14979 14773
rect 16853 14773 16865 14776
rect 16899 14773 16911 14807
rect 16853 14767 16911 14773
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18322 14804 18328 14816
rect 18012 14776 18328 14804
rect 18012 14764 18018 14776
rect 18322 14764 18328 14776
rect 18380 14804 18386 14816
rect 18509 14807 18567 14813
rect 18509 14804 18521 14807
rect 18380 14776 18521 14804
rect 18380 14764 18386 14776
rect 18509 14773 18521 14776
rect 18555 14804 18567 14807
rect 19794 14804 19800 14816
rect 18555 14776 19800 14804
rect 18555 14773 18567 14776
rect 18509 14767 18567 14773
rect 19794 14764 19800 14776
rect 19852 14764 19858 14816
rect 19978 14804 19984 14816
rect 19939 14776 19984 14804
rect 19978 14764 19984 14776
rect 20036 14764 20042 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2498 14560 2504 14612
rect 2556 14600 2562 14612
rect 2593 14603 2651 14609
rect 2593 14600 2605 14603
rect 2556 14572 2605 14600
rect 2556 14560 2562 14572
rect 2593 14569 2605 14572
rect 2639 14569 2651 14603
rect 3970 14600 3976 14612
rect 3931 14572 3976 14600
rect 2593 14563 2651 14569
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 5442 14600 5448 14612
rect 4212 14572 4936 14600
rect 5403 14572 5448 14600
rect 4212 14560 4218 14572
rect 3053 14535 3111 14541
rect 3053 14501 3065 14535
rect 3099 14532 3111 14535
rect 3510 14532 3516 14544
rect 3099 14504 3516 14532
rect 3099 14501 3111 14504
rect 3053 14495 3111 14501
rect 3510 14492 3516 14504
rect 3568 14532 3574 14544
rect 4246 14532 4252 14544
rect 3568 14504 4252 14532
rect 3568 14492 3574 14504
rect 4246 14492 4252 14504
rect 4304 14532 4310 14544
rect 4430 14532 4436 14544
rect 4304 14504 4436 14532
rect 4304 14492 4310 14504
rect 4430 14492 4436 14504
rect 4488 14492 4494 14544
rect 4525 14467 4583 14473
rect 4525 14464 4537 14467
rect 4356 14436 4537 14464
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14365 2191 14399
rect 2133 14359 2191 14365
rect 2148 14328 2176 14359
rect 2222 14356 2228 14408
rect 2280 14396 2286 14408
rect 2409 14399 2467 14405
rect 2409 14396 2421 14399
rect 2280 14368 2421 14396
rect 2280 14356 2286 14368
rect 2409 14365 2421 14368
rect 2455 14365 2467 14399
rect 2409 14359 2467 14365
rect 3326 14356 3332 14408
rect 3384 14396 3390 14408
rect 3694 14396 3700 14408
rect 3384 14368 3700 14396
rect 3384 14356 3390 14368
rect 3694 14356 3700 14368
rect 3752 14356 3758 14408
rect 2498 14328 2504 14340
rect 2148 14300 2504 14328
rect 2498 14288 2504 14300
rect 2556 14288 2562 14340
rect 3142 14288 3148 14340
rect 3200 14328 3206 14340
rect 3200 14300 4200 14328
rect 3200 14288 3206 14300
rect 3326 14260 3332 14272
rect 3287 14232 3332 14260
rect 3326 14220 3332 14232
rect 3384 14220 3390 14272
rect 4172 14260 4200 14300
rect 4246 14288 4252 14340
rect 4304 14328 4310 14340
rect 4356 14328 4384 14436
rect 4525 14433 4537 14436
rect 4571 14433 4583 14467
rect 4908 14464 4936 14572
rect 5442 14560 5448 14572
rect 5500 14560 5506 14612
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 6273 14603 6331 14609
rect 6273 14600 6285 14603
rect 5868 14572 6285 14600
rect 5868 14560 5874 14572
rect 6273 14569 6285 14572
rect 6319 14569 6331 14603
rect 6273 14563 6331 14569
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 7745 14603 7803 14609
rect 7745 14600 7757 14603
rect 7708 14572 7757 14600
rect 7708 14560 7714 14572
rect 7745 14569 7757 14572
rect 7791 14600 7803 14603
rect 8386 14600 8392 14612
rect 7791 14572 8392 14600
rect 7791 14569 7803 14572
rect 7745 14563 7803 14569
rect 8386 14560 8392 14572
rect 8444 14560 8450 14612
rect 8941 14603 8999 14609
rect 8941 14569 8953 14603
rect 8987 14600 8999 14603
rect 9306 14600 9312 14612
rect 8987 14572 9312 14600
rect 8987 14569 8999 14572
rect 8941 14563 8999 14569
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 10870 14600 10876 14612
rect 9416 14572 10876 14600
rect 4982 14492 4988 14544
rect 5040 14532 5046 14544
rect 9416 14532 9444 14572
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 11241 14603 11299 14609
rect 11241 14569 11253 14603
rect 11287 14600 11299 14603
rect 11514 14600 11520 14612
rect 11287 14572 11520 14600
rect 11287 14569 11299 14572
rect 11241 14563 11299 14569
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 15838 14600 15844 14612
rect 15751 14572 15844 14600
rect 15838 14560 15844 14572
rect 15896 14600 15902 14612
rect 19702 14600 19708 14612
rect 15896 14572 19708 14600
rect 15896 14560 15902 14572
rect 19702 14560 19708 14572
rect 19760 14560 19766 14612
rect 13814 14532 13820 14544
rect 5040 14504 9444 14532
rect 9600 14504 13820 14532
rect 5040 14492 5046 14504
rect 7377 14467 7435 14473
rect 7377 14464 7389 14467
rect 4908 14436 7389 14464
rect 4525 14427 4583 14433
rect 7377 14433 7389 14436
rect 7423 14464 7435 14467
rect 7650 14464 7656 14476
rect 7423 14436 7656 14464
rect 7423 14433 7435 14436
rect 7377 14427 7435 14433
rect 7650 14424 7656 14436
rect 7708 14464 7714 14476
rect 8018 14464 8024 14476
rect 7708 14436 8024 14464
rect 7708 14424 7714 14436
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 8294 14464 8300 14476
rect 8255 14436 8300 14464
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 9122 14424 9128 14476
rect 9180 14464 9186 14476
rect 9600 14473 9628 14504
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 16574 14532 16580 14544
rect 16535 14504 16580 14532
rect 16574 14492 16580 14504
rect 16632 14492 16638 14544
rect 17954 14492 17960 14544
rect 18012 14532 18018 14544
rect 19889 14535 19947 14541
rect 19889 14532 19901 14535
rect 18012 14504 19901 14532
rect 18012 14492 18018 14504
rect 19889 14501 19901 14504
rect 19935 14501 19947 14535
rect 19889 14495 19947 14501
rect 9401 14467 9459 14473
rect 9401 14464 9413 14467
rect 9180 14436 9413 14464
rect 9180 14424 9186 14436
rect 9401 14433 9413 14436
rect 9447 14433 9459 14467
rect 9401 14427 9459 14433
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14433 9643 14467
rect 10686 14464 10692 14476
rect 10647 14436 10692 14464
rect 9585 14427 9643 14433
rect 4433 14399 4491 14405
rect 4433 14365 4445 14399
rect 4479 14396 4491 14399
rect 5350 14396 5356 14408
rect 4479 14368 5356 14396
rect 4479 14365 4491 14368
rect 4433 14359 4491 14365
rect 5350 14356 5356 14368
rect 5408 14396 5414 14408
rect 5721 14399 5779 14405
rect 5721 14396 5733 14399
rect 5408 14368 5733 14396
rect 5408 14356 5414 14368
rect 5721 14365 5733 14368
rect 5767 14365 5779 14399
rect 5721 14359 5779 14365
rect 7558 14356 7564 14408
rect 7616 14396 7622 14408
rect 8113 14399 8171 14405
rect 8113 14396 8125 14399
rect 7616 14368 8125 14396
rect 7616 14356 7622 14368
rect 8113 14365 8125 14368
rect 8159 14365 8171 14399
rect 8113 14359 8171 14365
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 9306 14396 9312 14408
rect 8536 14368 9312 14396
rect 8536 14356 8542 14368
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9416 14396 9444 14427
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 19702 14424 19708 14476
rect 19760 14464 19766 14476
rect 20162 14464 20168 14476
rect 19760 14436 20168 14464
rect 19760 14424 19766 14436
rect 20162 14424 20168 14436
rect 20220 14424 20226 14476
rect 9953 14399 10011 14405
rect 9953 14396 9965 14399
rect 9416 14368 9965 14396
rect 9953 14365 9965 14368
rect 9999 14365 10011 14399
rect 13538 14396 13544 14408
rect 9953 14359 10011 14365
rect 10060 14368 13544 14396
rect 5077 14331 5135 14337
rect 5077 14328 5089 14331
rect 4304 14300 5089 14328
rect 4304 14288 4310 14300
rect 5077 14297 5089 14300
rect 5123 14328 5135 14331
rect 10060 14328 10088 14368
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 13722 14356 13728 14408
rect 13780 14396 13786 14408
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 13780 14368 14473 14396
rect 13780 14356 13786 14368
rect 14461 14365 14473 14368
rect 14507 14396 14519 14399
rect 15010 14396 15016 14408
rect 14507 14368 15016 14396
rect 14507 14365 14519 14368
rect 14461 14359 14519 14365
rect 15010 14356 15016 14368
rect 15068 14396 15074 14408
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 15068 14368 16129 14396
rect 15068 14356 15074 14368
rect 16117 14365 16129 14368
rect 16163 14396 16175 14399
rect 17957 14399 18015 14405
rect 17957 14396 17969 14399
rect 16163 14368 17969 14396
rect 16163 14365 16175 14368
rect 16117 14359 16175 14365
rect 17957 14365 17969 14368
rect 18003 14396 18015 14399
rect 18233 14399 18291 14405
rect 18233 14396 18245 14399
rect 18003 14368 18245 14396
rect 18003 14365 18015 14368
rect 17957 14359 18015 14365
rect 18233 14365 18245 14368
rect 18279 14396 18291 14399
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 18279 14368 19257 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 19245 14365 19257 14368
rect 19291 14396 19303 14399
rect 21269 14399 21327 14405
rect 21269 14396 21281 14399
rect 19291 14368 21281 14396
rect 19291 14365 19303 14368
rect 19245 14359 19303 14365
rect 20824 14340 20852 14368
rect 21269 14365 21281 14368
rect 21315 14365 21327 14399
rect 21269 14359 21327 14365
rect 5123 14300 10088 14328
rect 10152 14300 14504 14328
rect 5123 14297 5135 14300
rect 5077 14291 5135 14297
rect 4341 14263 4399 14269
rect 4341 14260 4353 14263
rect 4172 14232 4353 14260
rect 4341 14229 4353 14232
rect 4387 14260 4399 14263
rect 4614 14260 4620 14272
rect 4387 14232 4620 14260
rect 4387 14229 4399 14232
rect 4341 14223 4399 14229
rect 4614 14220 4620 14232
rect 4672 14220 4678 14272
rect 6733 14263 6791 14269
rect 6733 14229 6745 14263
rect 6779 14260 6791 14263
rect 6822 14260 6828 14272
rect 6779 14232 6828 14260
rect 6779 14229 6791 14232
rect 6733 14223 6791 14229
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 7006 14220 7012 14272
rect 7064 14260 7070 14272
rect 10152 14260 10180 14300
rect 10778 14260 10784 14272
rect 7064 14232 10180 14260
rect 10739 14232 10784 14260
rect 7064 14220 7070 14232
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 10870 14220 10876 14272
rect 10928 14260 10934 14272
rect 13722 14260 13728 14272
rect 10928 14232 10973 14260
rect 13683 14232 13728 14260
rect 10928 14220 10934 14232
rect 13722 14220 13728 14232
rect 13780 14260 13786 14272
rect 14093 14263 14151 14269
rect 14093 14260 14105 14263
rect 13780 14232 14105 14260
rect 13780 14220 13786 14232
rect 14093 14229 14105 14232
rect 14139 14229 14151 14263
rect 14476 14260 14504 14300
rect 14550 14288 14556 14340
rect 14608 14328 14614 14340
rect 14706 14331 14764 14337
rect 14706 14328 14718 14331
rect 14608 14300 14718 14328
rect 14608 14288 14614 14300
rect 14706 14297 14718 14300
rect 14752 14297 14764 14331
rect 17402 14328 17408 14340
rect 14706 14291 14764 14297
rect 16500 14300 17408 14328
rect 16500 14260 16528 14300
rect 17402 14288 17408 14300
rect 17460 14288 17466 14340
rect 17678 14288 17684 14340
rect 17736 14337 17742 14340
rect 17736 14328 17748 14337
rect 20438 14328 20444 14340
rect 17736 14300 17781 14328
rect 18800 14300 20444 14328
rect 17736 14291 17748 14300
rect 17736 14288 17742 14291
rect 14476 14232 16528 14260
rect 14093 14223 14151 14229
rect 16574 14220 16580 14272
rect 16632 14260 16638 14272
rect 17310 14260 17316 14272
rect 16632 14232 17316 14260
rect 16632 14220 16638 14232
rect 17310 14220 17316 14232
rect 17368 14220 17374 14272
rect 17420 14260 17448 14288
rect 18230 14260 18236 14272
rect 17420 14232 18236 14260
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 18690 14220 18696 14272
rect 18748 14260 18754 14272
rect 18800 14269 18828 14300
rect 20438 14288 20444 14300
rect 20496 14328 20502 14340
rect 20496 14300 20760 14328
rect 20496 14288 20502 14300
rect 18785 14263 18843 14269
rect 18785 14260 18797 14263
rect 18748 14232 18797 14260
rect 18748 14220 18754 14232
rect 18785 14229 18797 14232
rect 18831 14229 18843 14263
rect 20732 14260 20760 14300
rect 20806 14288 20812 14340
rect 20864 14288 20870 14340
rect 21002 14331 21060 14337
rect 21002 14328 21014 14331
rect 20916 14300 21014 14328
rect 20916 14260 20944 14300
rect 21002 14297 21014 14300
rect 21048 14297 21060 14331
rect 21002 14291 21060 14297
rect 20732 14232 20944 14260
rect 18785 14223 18843 14229
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 1673 14059 1731 14065
rect 1673 14056 1685 14059
rect 1452 14028 1685 14056
rect 1452 14016 1458 14028
rect 1673 14025 1685 14028
rect 1719 14025 1731 14059
rect 1673 14019 1731 14025
rect 2409 14059 2467 14065
rect 2409 14025 2421 14059
rect 2455 14056 2467 14059
rect 3053 14059 3111 14065
rect 3053 14056 3065 14059
rect 2455 14028 3065 14056
rect 2455 14025 2467 14028
rect 2409 14019 2467 14025
rect 3053 14025 3065 14028
rect 3099 14025 3111 14059
rect 3053 14019 3111 14025
rect 3421 14059 3479 14065
rect 3421 14025 3433 14059
rect 3467 14056 3479 14059
rect 3510 14056 3516 14068
rect 3467 14028 3516 14056
rect 3467 14025 3479 14028
rect 3421 14019 3479 14025
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 4246 14056 4252 14068
rect 4207 14028 4252 14056
rect 4246 14016 4252 14028
rect 4304 14016 4310 14068
rect 4798 14016 4804 14068
rect 4856 14056 4862 14068
rect 4856 14028 5304 14056
rect 4856 14016 4862 14028
rect 5169 13991 5227 13997
rect 5169 13988 5181 13991
rect 3712 13960 5181 13988
rect 3712 13920 3740 13960
rect 5169 13957 5181 13960
rect 5215 13957 5227 13991
rect 5276 13988 5304 14028
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 5592 14028 5641 14056
rect 5592 14016 5598 14028
rect 5629 14025 5641 14028
rect 5675 14025 5687 14059
rect 7006 14056 7012 14068
rect 5629 14019 5687 14025
rect 5736 14028 7012 14056
rect 5736 13988 5764 14028
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7098 14016 7104 14068
rect 7156 14056 7162 14068
rect 7193 14059 7251 14065
rect 7193 14056 7205 14059
rect 7156 14028 7205 14056
rect 7156 14016 7162 14028
rect 7193 14025 7205 14028
rect 7239 14025 7251 14059
rect 7193 14019 7251 14025
rect 8021 14059 8079 14065
rect 8021 14025 8033 14059
rect 8067 14056 8079 14059
rect 8110 14056 8116 14068
rect 8067 14028 8116 14056
rect 8067 14025 8079 14028
rect 8021 14019 8079 14025
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 8389 14059 8447 14065
rect 8389 14025 8401 14059
rect 8435 14056 8447 14059
rect 8570 14056 8576 14068
rect 8435 14028 8576 14056
rect 8435 14025 8447 14028
rect 8389 14019 8447 14025
rect 8570 14016 8576 14028
rect 8628 14056 8634 14068
rect 9033 14059 9091 14065
rect 9033 14056 9045 14059
rect 8628 14028 9045 14056
rect 8628 14016 8634 14028
rect 9033 14025 9045 14028
rect 9079 14025 9091 14059
rect 9033 14019 9091 14025
rect 9122 14016 9128 14068
rect 9180 14056 9186 14068
rect 9306 14056 9312 14068
rect 9180 14028 9312 14056
rect 9180 14016 9186 14028
rect 9306 14016 9312 14028
rect 9364 14056 9370 14068
rect 9401 14059 9459 14065
rect 9401 14056 9413 14059
rect 9364 14028 9413 14056
rect 9364 14016 9370 14028
rect 9401 14025 9413 14028
rect 9447 14025 9459 14059
rect 9401 14019 9459 14025
rect 9861 14059 9919 14065
rect 9861 14025 9873 14059
rect 9907 14056 9919 14059
rect 10042 14056 10048 14068
rect 9907 14028 10048 14056
rect 9907 14025 9919 14028
rect 9861 14019 9919 14025
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 10870 14056 10876 14068
rect 10831 14028 10876 14056
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 13538 14016 13544 14068
rect 13596 14056 13602 14068
rect 13596 14028 14872 14056
rect 13596 14016 13602 14028
rect 5276 13960 5764 13988
rect 5997 13991 6055 13997
rect 5169 13951 5227 13957
rect 5997 13957 6009 13991
rect 6043 13988 6055 13991
rect 10962 13988 10968 14000
rect 6043 13960 10968 13988
rect 6043 13957 6055 13960
rect 5997 13951 6055 13957
rect 2884 13892 3740 13920
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13821 2191 13855
rect 2314 13852 2320 13864
rect 2275 13824 2320 13852
rect 2133 13815 2191 13821
rect 1854 13744 1860 13796
rect 1912 13784 1918 13796
rect 2148 13784 2176 13815
rect 2314 13812 2320 13824
rect 2372 13812 2378 13864
rect 1912 13756 2176 13784
rect 2777 13787 2835 13793
rect 1912 13744 1918 13756
rect 2777 13753 2789 13787
rect 2823 13784 2835 13787
rect 2884 13784 2912 13892
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 4212 13892 5273 13920
rect 4212 13880 4218 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 3513 13855 3571 13861
rect 3513 13852 3525 13855
rect 2823 13756 2912 13784
rect 3160 13824 3525 13852
rect 2823 13753 2835 13756
rect 2777 13747 2835 13753
rect 2406 13676 2412 13728
rect 2464 13716 2470 13728
rect 3160 13716 3188 13824
rect 3513 13821 3525 13824
rect 3559 13821 3571 13855
rect 3513 13815 3571 13821
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13821 3663 13855
rect 3605 13815 3663 13821
rect 3326 13744 3332 13796
rect 3384 13784 3390 13796
rect 3620 13784 3648 13815
rect 3694 13812 3700 13864
rect 3752 13852 3758 13864
rect 4798 13852 4804 13864
rect 3752 13824 4804 13852
rect 3752 13812 3758 13824
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13821 5135 13855
rect 5077 13815 5135 13821
rect 3384 13756 3648 13784
rect 3384 13744 3390 13756
rect 4062 13744 4068 13796
rect 4120 13784 4126 13796
rect 4706 13784 4712 13796
rect 4120 13756 4712 13784
rect 4120 13744 4126 13756
rect 4706 13744 4712 13756
rect 4764 13744 4770 13796
rect 5092 13784 5120 13815
rect 5166 13812 5172 13864
rect 5224 13852 5230 13864
rect 6012 13852 6040 13951
rect 10962 13948 10968 13960
rect 11020 13948 11026 14000
rect 12526 13948 12532 14000
rect 12584 13988 12590 14000
rect 12584 13960 13584 13988
rect 12584 13948 12590 13960
rect 6825 13923 6883 13929
rect 6825 13889 6837 13923
rect 6871 13920 6883 13923
rect 7469 13923 7527 13929
rect 7469 13920 7481 13923
rect 6871 13892 7481 13920
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 7469 13889 7481 13892
rect 7515 13889 7527 13923
rect 7469 13883 7527 13889
rect 8386 13880 8392 13932
rect 8444 13920 8450 13932
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 8444 13892 8493 13920
rect 8444 13880 8450 13892
rect 8481 13889 8493 13892
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 10042 13920 10048 13932
rect 9732 13892 10048 13920
rect 9732 13880 9738 13892
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10226 13920 10232 13932
rect 10187 13892 10232 13920
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 13285 13923 13343 13929
rect 13285 13889 13297 13923
rect 13331 13920 13343 13923
rect 13446 13920 13452 13932
rect 13331 13892 13452 13920
rect 13331 13889 13343 13892
rect 13285 13883 13343 13889
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 13556 13920 13584 13960
rect 14084 13923 14142 13929
rect 14084 13920 14096 13923
rect 13556 13892 14096 13920
rect 14084 13889 14096 13892
rect 14130 13920 14142 13923
rect 14458 13920 14464 13932
rect 14130 13892 14464 13920
rect 14130 13889 14142 13892
rect 14084 13883 14142 13889
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 14844 13920 14872 14028
rect 14918 14016 14924 14068
rect 14976 14056 14982 14068
rect 15197 14059 15255 14065
rect 15197 14056 15209 14059
rect 14976 14028 15209 14056
rect 14976 14016 14982 14028
rect 15197 14025 15209 14028
rect 15243 14056 15255 14059
rect 17034 14056 17040 14068
rect 15243 14028 17040 14056
rect 15243 14025 15255 14028
rect 15197 14019 15255 14025
rect 17034 14016 17040 14028
rect 17092 14016 17098 14068
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 17678 14016 17684 14068
rect 17736 14056 17742 14068
rect 19794 14056 19800 14068
rect 17736 14028 19800 14056
rect 17736 14016 17742 14028
rect 19794 14016 19800 14028
rect 19852 14016 19858 14068
rect 20714 14056 20720 14068
rect 20088 14028 20720 14056
rect 15010 13948 15016 14000
rect 15068 13988 15074 14000
rect 15473 13991 15531 13997
rect 15473 13988 15485 13991
rect 15068 13960 15485 13988
rect 15068 13948 15074 13960
rect 15473 13957 15485 13960
rect 15519 13988 15531 13991
rect 16669 13991 16727 13997
rect 16669 13988 16681 13991
rect 15519 13960 16681 13988
rect 15519 13957 15531 13960
rect 15473 13951 15531 13957
rect 16669 13957 16681 13960
rect 16715 13957 16727 13991
rect 18518 13991 18576 13997
rect 18518 13988 18530 13991
rect 16669 13951 16727 13957
rect 16776 13960 18530 13988
rect 16776 13920 16804 13960
rect 18518 13957 18530 13960
rect 18564 13988 18576 13991
rect 18564 13960 19334 13988
rect 18564 13957 18576 13960
rect 18518 13951 18576 13957
rect 14844 13892 16804 13920
rect 19306 13920 19334 13960
rect 20088 13920 20116 14028
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 19306 13892 20116 13920
rect 20162 13880 20168 13932
rect 20220 13929 20226 13932
rect 20220 13920 20232 13929
rect 20441 13923 20499 13929
rect 20220 13892 20265 13920
rect 20220 13883 20232 13892
rect 20441 13889 20453 13923
rect 20487 13920 20499 13923
rect 20806 13920 20812 13932
rect 20487 13892 20812 13920
rect 20487 13889 20499 13892
rect 20441 13883 20499 13889
rect 20220 13880 20226 13883
rect 20806 13880 20812 13892
rect 20864 13920 20870 13932
rect 21177 13923 21235 13929
rect 21177 13920 21189 13923
rect 20864 13892 21189 13920
rect 20864 13880 20870 13892
rect 21177 13889 21189 13892
rect 21223 13889 21235 13923
rect 21177 13883 21235 13889
rect 5224 13824 6040 13852
rect 6641 13855 6699 13861
rect 5224 13812 5230 13824
rect 6641 13821 6653 13855
rect 6687 13821 6699 13855
rect 6641 13815 6699 13821
rect 6733 13855 6791 13861
rect 6733 13821 6745 13855
rect 6779 13852 6791 13855
rect 7834 13852 7840 13864
rect 6779 13824 7840 13852
rect 6779 13821 6791 13824
rect 6733 13815 6791 13821
rect 5442 13784 5448 13796
rect 5092 13756 5448 13784
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 6656 13784 6684 13815
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13821 8723 13855
rect 10318 13852 10324 13864
rect 10279 13824 10324 13852
rect 8665 13815 8723 13821
rect 7098 13784 7104 13796
rect 6656 13756 7104 13784
rect 4614 13716 4620 13728
rect 2464 13688 3188 13716
rect 4575 13688 4620 13716
rect 2464 13676 2470 13688
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 5074 13676 5080 13728
rect 5132 13716 5138 13728
rect 6656 13716 6684 13756
rect 7098 13744 7104 13756
rect 7156 13744 7162 13796
rect 8680 13784 8708 13815
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13852 10563 13855
rect 12250 13852 12256 13864
rect 10551 13824 12256 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 13541 13855 13599 13861
rect 13541 13821 13553 13855
rect 13587 13852 13599 13855
rect 13722 13852 13728 13864
rect 13587 13824 13728 13852
rect 13587 13821 13599 13824
rect 13541 13815 13599 13821
rect 13722 13812 13728 13824
rect 13780 13852 13786 13864
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 13780 13824 13829 13852
rect 13780 13812 13786 13824
rect 13817 13821 13829 13824
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 18785 13855 18843 13861
rect 18785 13821 18797 13855
rect 18831 13821 18843 13855
rect 18785 13815 18843 13821
rect 9490 13784 9496 13796
rect 8680 13756 9496 13784
rect 9490 13744 9496 13756
rect 9548 13784 9554 13796
rect 9548 13756 12434 13784
rect 9548 13744 9554 13756
rect 5132 13688 6684 13716
rect 5132 13676 5138 13688
rect 6914 13676 6920 13728
rect 6972 13716 6978 13728
rect 8386 13716 8392 13728
rect 6972 13688 8392 13716
rect 6972 13676 6978 13688
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 12161 13719 12219 13725
rect 12161 13685 12173 13719
rect 12207 13716 12219 13719
rect 12250 13716 12256 13728
rect 12207 13688 12256 13716
rect 12207 13685 12219 13688
rect 12161 13679 12219 13685
rect 12250 13676 12256 13688
rect 12308 13676 12314 13728
rect 12406 13716 12434 13756
rect 15470 13716 15476 13728
rect 12406 13688 15476 13716
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 18046 13676 18052 13728
rect 18104 13716 18110 13728
rect 18800 13716 18828 13815
rect 19058 13716 19064 13728
rect 18104 13688 18828 13716
rect 19019 13688 19064 13716
rect 18104 13676 18110 13688
rect 19058 13676 19064 13688
rect 19116 13676 19122 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 2685 13515 2743 13521
rect 2685 13512 2697 13515
rect 2372 13484 2697 13512
rect 2372 13472 2378 13484
rect 2685 13481 2697 13484
rect 2731 13481 2743 13515
rect 2685 13475 2743 13481
rect 3878 13472 3884 13524
rect 3936 13512 3942 13524
rect 3973 13515 4031 13521
rect 3973 13512 3985 13515
rect 3936 13484 3985 13512
rect 3936 13472 3942 13484
rect 3973 13481 3985 13484
rect 4019 13481 4031 13515
rect 3973 13475 4031 13481
rect 4062 13472 4068 13524
rect 4120 13512 4126 13524
rect 4522 13512 4528 13524
rect 4120 13484 4528 13512
rect 4120 13472 4126 13484
rect 4522 13472 4528 13484
rect 4580 13472 4586 13524
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6365 13515 6423 13521
rect 6365 13512 6377 13515
rect 6052 13484 6377 13512
rect 6052 13472 6058 13484
rect 6365 13481 6377 13484
rect 6411 13481 6423 13515
rect 7834 13512 7840 13524
rect 7795 13484 7840 13512
rect 6365 13475 6423 13481
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 8570 13472 8576 13524
rect 8628 13512 8634 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8628 13484 8953 13512
rect 8628 13472 8634 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 9306 13512 9312 13524
rect 9267 13484 9312 13512
rect 8941 13475 8999 13481
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 10468 13484 10517 13512
rect 10468 13472 10474 13484
rect 10505 13481 10517 13484
rect 10551 13512 10563 13515
rect 13170 13512 13176 13524
rect 10551 13484 11376 13512
rect 10551 13481 10563 13484
rect 10505 13475 10563 13481
rect 2041 13447 2099 13453
rect 2041 13413 2053 13447
rect 2087 13444 2099 13447
rect 4430 13444 4436 13456
rect 2087 13416 4436 13444
rect 2087 13413 2099 13416
rect 2041 13407 2099 13413
rect 4430 13404 4436 13416
rect 4488 13404 4494 13456
rect 5813 13447 5871 13453
rect 5813 13413 5825 13447
rect 5859 13444 5871 13447
rect 6546 13444 6552 13456
rect 5859 13416 6552 13444
rect 5859 13413 5871 13416
rect 5813 13407 5871 13413
rect 6546 13404 6552 13416
rect 6604 13404 6610 13456
rect 7190 13444 7196 13456
rect 6932 13416 7196 13444
rect 1394 13336 1400 13388
rect 1452 13376 1458 13388
rect 2317 13379 2375 13385
rect 2317 13376 2329 13379
rect 1452 13348 2329 13376
rect 1452 13336 1458 13348
rect 2317 13345 2329 13348
rect 2363 13376 2375 13379
rect 2406 13376 2412 13388
rect 2363 13348 2412 13376
rect 2363 13345 2375 13348
rect 2317 13339 2375 13345
rect 2406 13336 2412 13348
rect 2464 13336 2470 13388
rect 3326 13376 3332 13388
rect 3239 13348 3332 13376
rect 3326 13336 3332 13348
rect 3384 13376 3390 13388
rect 3510 13376 3516 13388
rect 3384 13348 3516 13376
rect 3384 13336 3390 13348
rect 3510 13336 3516 13348
rect 3568 13336 3574 13388
rect 4246 13336 4252 13388
rect 4304 13376 4310 13388
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 4304 13348 4537 13376
rect 4304 13336 4310 13348
rect 4525 13345 4537 13348
rect 4571 13345 4583 13379
rect 5166 13376 5172 13388
rect 5127 13348 5172 13376
rect 4525 13339 4583 13345
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 5350 13376 5356 13388
rect 5311 13348 5356 13376
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 3142 13308 3148 13320
rect 3099 13280 3148 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 4614 13268 4620 13320
rect 4672 13308 4678 13320
rect 5445 13311 5503 13317
rect 5445 13308 5457 13311
rect 4672 13280 5457 13308
rect 4672 13268 4678 13280
rect 5445 13277 5457 13280
rect 5491 13277 5503 13311
rect 5445 13271 5503 13277
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 6932 13308 6960 13416
rect 7190 13404 7196 13416
rect 7248 13404 7254 13456
rect 8588 13444 8616 13472
rect 8312 13416 8616 13444
rect 8312 13385 8340 13416
rect 7009 13379 7067 13385
rect 7009 13345 7021 13379
rect 7055 13345 7067 13379
rect 7009 13339 7067 13345
rect 8297 13379 8355 13385
rect 8297 13345 8309 13379
rect 8343 13345 8355 13379
rect 8297 13339 8355 13345
rect 6604 13280 6960 13308
rect 7024 13308 7052 13339
rect 8386 13336 8392 13388
rect 8444 13376 8450 13388
rect 8481 13379 8539 13385
rect 8481 13376 8493 13379
rect 8444 13348 8493 13376
rect 8444 13336 8450 13348
rect 8481 13345 8493 13348
rect 8527 13376 8539 13379
rect 9950 13376 9956 13388
rect 8527 13348 9956 13376
rect 8527 13345 8539 13348
rect 8481 13339 8539 13345
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10226 13376 10232 13388
rect 10187 13348 10232 13376
rect 10226 13336 10232 13348
rect 10284 13336 10290 13388
rect 11348 13385 11376 13484
rect 11532 13484 13176 13512
rect 11532 13385 11560 13484
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 14734 13512 14740 13524
rect 13964 13484 14740 13512
rect 13964 13472 13970 13484
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 15473 13515 15531 13521
rect 15473 13512 15485 13515
rect 15344 13484 15485 13512
rect 15344 13472 15350 13484
rect 15473 13481 15485 13484
rect 15519 13512 15531 13515
rect 17034 13512 17040 13524
rect 15519 13484 17040 13512
rect 15519 13481 15531 13484
rect 15473 13475 15531 13481
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 19518 13512 19524 13524
rect 19479 13484 19524 13512
rect 19518 13472 19524 13484
rect 19576 13512 19582 13524
rect 20162 13512 20168 13524
rect 19576 13484 20168 13512
rect 19576 13472 19582 13484
rect 20162 13472 20168 13484
rect 20220 13512 20226 13524
rect 21177 13515 21235 13521
rect 21177 13512 21189 13515
rect 20220 13484 21189 13512
rect 20220 13472 20226 13484
rect 21177 13481 21189 13484
rect 21223 13481 21235 13515
rect 21177 13475 21235 13481
rect 18874 13444 18880 13456
rect 18835 13416 18880 13444
rect 18874 13404 18880 13416
rect 18932 13404 18938 13456
rect 11333 13379 11391 13385
rect 11333 13345 11345 13379
rect 11379 13345 11391 13379
rect 11333 13339 11391 13345
rect 11517 13379 11575 13385
rect 11517 13345 11529 13379
rect 11563 13345 11575 13379
rect 11517 13339 11575 13345
rect 12158 13308 12164 13320
rect 7024 13280 11468 13308
rect 12119 13280 12164 13308
rect 6604 13268 6610 13280
rect 2406 13200 2412 13252
rect 2464 13240 2470 13252
rect 4433 13243 4491 13249
rect 4433 13240 4445 13243
rect 2464 13212 4445 13240
rect 2464 13200 2470 13212
rect 4433 13209 4445 13212
rect 4479 13240 4491 13243
rect 5258 13240 5264 13252
rect 4479 13212 5264 13240
rect 4479 13209 4491 13212
rect 4433 13203 4491 13209
rect 5258 13200 5264 13212
rect 5316 13200 5322 13252
rect 6733 13243 6791 13249
rect 6733 13209 6745 13243
rect 6779 13240 6791 13243
rect 7377 13243 7435 13249
rect 7377 13240 7389 13243
rect 6779 13212 7389 13240
rect 6779 13209 6791 13212
rect 6733 13203 6791 13209
rect 7377 13209 7389 13212
rect 7423 13209 7435 13243
rect 7377 13203 7435 13209
rect 10594 13200 10600 13252
rect 10652 13240 10658 13252
rect 10962 13240 10968 13252
rect 10652 13212 10968 13240
rect 10652 13200 10658 13212
rect 10962 13200 10968 13212
rect 11020 13240 11026 13252
rect 11241 13243 11299 13249
rect 11241 13240 11253 13243
rect 11020 13212 11253 13240
rect 11020 13200 11026 13212
rect 11241 13209 11253 13212
rect 11287 13209 11299 13243
rect 11241 13203 11299 13209
rect 1673 13175 1731 13181
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 1854 13172 1860 13184
rect 1719 13144 1860 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 3145 13175 3203 13181
rect 3145 13141 3157 13175
rect 3191 13172 3203 13175
rect 3970 13172 3976 13184
rect 3191 13144 3976 13172
rect 3191 13141 3203 13144
rect 3145 13135 3203 13141
rect 3970 13132 3976 13144
rect 4028 13132 4034 13184
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 4304 13144 4353 13172
rect 4304 13132 4310 13144
rect 4341 13141 4353 13144
rect 4387 13172 4399 13175
rect 4522 13172 4528 13184
rect 4387 13144 4528 13172
rect 4387 13141 4399 13144
rect 4341 13135 4399 13141
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 6880 13144 6925 13172
rect 6880 13132 6886 13144
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 8205 13175 8263 13181
rect 8205 13172 8217 13175
rect 7708 13144 8217 13172
rect 7708 13132 7714 13144
rect 8205 13141 8217 13144
rect 8251 13141 8263 13175
rect 10870 13172 10876 13184
rect 10831 13144 10876 13172
rect 8205 13135 8263 13141
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 11440 13172 11468 13280
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 13722 13268 13728 13320
rect 13780 13308 13786 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 13780 13280 14105 13308
rect 13780 13268 13786 13280
rect 14093 13277 14105 13280
rect 14139 13308 14151 13311
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 14139 13280 15761 13308
rect 14139 13277 14151 13280
rect 14093 13271 14151 13277
rect 15749 13277 15761 13280
rect 15795 13308 15807 13311
rect 17497 13311 17555 13317
rect 17497 13308 17509 13311
rect 15795 13280 17509 13308
rect 15795 13277 15807 13280
rect 15749 13271 15807 13277
rect 17497 13277 17509 13280
rect 17543 13308 17555 13311
rect 18046 13308 18052 13320
rect 17543 13280 18052 13308
rect 17543 13277 17555 13280
rect 17497 13271 17555 13277
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 20806 13268 20812 13320
rect 20864 13308 20870 13320
rect 20901 13311 20959 13317
rect 20901 13308 20913 13311
rect 20864 13280 20913 13308
rect 20864 13268 20870 13280
rect 20901 13277 20913 13280
rect 20947 13277 20959 13311
rect 20901 13271 20959 13277
rect 12250 13200 12256 13252
rect 12308 13240 12314 13252
rect 12406 13243 12464 13249
rect 12406 13240 12418 13243
rect 12308 13212 12418 13240
rect 12308 13200 12314 13212
rect 12406 13209 12418 13212
rect 12452 13209 12464 13243
rect 12406 13203 12464 13209
rect 13630 13200 13636 13252
rect 13688 13240 13694 13252
rect 14338 13243 14396 13249
rect 14338 13240 14350 13243
rect 13688 13212 14350 13240
rect 13688 13200 13694 13212
rect 14338 13209 14350 13212
rect 14384 13240 14396 13243
rect 14384 13209 14412 13240
rect 14338 13203 14412 13209
rect 13078 13172 13084 13184
rect 11440 13144 13084 13172
rect 13078 13132 13084 13144
rect 13136 13132 13142 13184
rect 13354 13132 13360 13184
rect 13412 13172 13418 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 13412 13144 13553 13172
rect 13412 13132 13418 13144
rect 13541 13141 13553 13144
rect 13587 13141 13599 13175
rect 14384 13172 14412 13203
rect 14458 13200 14464 13252
rect 14516 13240 14522 13252
rect 17742 13243 17800 13249
rect 17742 13240 17754 13243
rect 14516 13212 17754 13240
rect 14516 13200 14522 13212
rect 17742 13209 17754 13212
rect 17788 13240 17800 13243
rect 19334 13240 19340 13252
rect 17788 13212 19340 13240
rect 17788 13209 17800 13212
rect 17742 13203 17800 13209
rect 19334 13200 19340 13212
rect 19392 13240 19398 13252
rect 19978 13240 19984 13252
rect 19392 13212 19984 13240
rect 19392 13200 19398 13212
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 20070 13200 20076 13252
rect 20128 13240 20134 13252
rect 20656 13243 20714 13249
rect 20656 13240 20668 13243
rect 20128 13212 20668 13240
rect 20128 13200 20134 13212
rect 20656 13209 20668 13212
rect 20702 13240 20714 13243
rect 21082 13240 21088 13252
rect 20702 13212 21088 13240
rect 20702 13209 20714 13212
rect 20656 13203 20714 13209
rect 21082 13200 21088 13212
rect 21140 13200 21146 13252
rect 19610 13172 19616 13184
rect 14384 13144 19616 13172
rect 13541 13135 13599 13141
rect 19610 13132 19616 13144
rect 19668 13132 19674 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 1489 12971 1547 12977
rect 1489 12937 1501 12971
rect 1535 12968 1547 12971
rect 3142 12968 3148 12980
rect 1535 12940 3148 12968
rect 1535 12937 1547 12940
rect 1489 12931 1547 12937
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 5258 12968 5264 12980
rect 5219 12940 5264 12968
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 5350 12928 5356 12980
rect 5408 12928 5414 12980
rect 7101 12971 7159 12977
rect 7101 12937 7113 12971
rect 7147 12968 7159 12971
rect 7282 12968 7288 12980
rect 7147 12940 7288 12968
rect 7147 12937 7159 12940
rect 7101 12931 7159 12937
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 7653 12971 7711 12977
rect 7653 12937 7665 12971
rect 7699 12937 7711 12971
rect 7653 12931 7711 12937
rect 8113 12971 8171 12977
rect 8113 12937 8125 12971
rect 8159 12968 8171 12971
rect 8665 12971 8723 12977
rect 8665 12968 8677 12971
rect 8159 12940 8677 12968
rect 8159 12937 8171 12940
rect 8113 12931 8171 12937
rect 8665 12937 8677 12940
rect 8711 12937 8723 12971
rect 8665 12931 8723 12937
rect 9125 12971 9183 12977
rect 9125 12937 9137 12971
rect 9171 12968 9183 12971
rect 9214 12968 9220 12980
rect 9171 12940 9220 12968
rect 9171 12937 9183 12940
rect 9125 12931 9183 12937
rect 1949 12903 2007 12909
rect 1949 12869 1961 12903
rect 1995 12900 2007 12903
rect 2590 12900 2596 12912
rect 1995 12872 2596 12900
rect 1995 12869 2007 12872
rect 1949 12863 2007 12869
rect 2590 12860 2596 12872
rect 2648 12860 2654 12912
rect 3970 12860 3976 12912
rect 4028 12900 4034 12912
rect 4157 12903 4215 12909
rect 4157 12900 4169 12903
rect 4028 12872 4169 12900
rect 4028 12860 4034 12872
rect 4157 12869 4169 12872
rect 4203 12900 4215 12903
rect 5368 12900 5396 12928
rect 4203 12872 5396 12900
rect 4203 12869 4215 12872
rect 4157 12863 4215 12869
rect 6638 12860 6644 12912
rect 6696 12900 6702 12912
rect 7668 12900 7696 12931
rect 9214 12928 9220 12940
rect 9272 12968 9278 12980
rect 9677 12971 9735 12977
rect 9677 12968 9689 12971
rect 9272 12940 9689 12968
rect 9272 12928 9278 12940
rect 9677 12937 9689 12940
rect 9723 12937 9735 12971
rect 10594 12968 10600 12980
rect 10555 12940 10600 12968
rect 9677 12931 9735 12937
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 11146 12928 11152 12980
rect 11204 12968 11210 12980
rect 11974 12968 11980 12980
rect 11204 12940 11980 12968
rect 11204 12928 11210 12940
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 13446 12968 13452 12980
rect 12492 12940 13452 12968
rect 12492 12928 12498 12940
rect 13446 12928 13452 12940
rect 13504 12968 13510 12980
rect 16669 12971 16727 12977
rect 16669 12968 16681 12971
rect 13504 12940 16681 12968
rect 13504 12928 13510 12940
rect 16669 12937 16681 12940
rect 16715 12937 16727 12971
rect 19334 12968 19340 12980
rect 19295 12940 19340 12968
rect 16669 12931 16727 12937
rect 19334 12928 19340 12940
rect 19392 12928 19398 12980
rect 19794 12968 19800 12980
rect 19755 12940 19800 12968
rect 19794 12928 19800 12940
rect 19852 12928 19858 12980
rect 6696 12872 7696 12900
rect 6696 12860 6702 12872
rect 7834 12860 7840 12912
rect 7892 12900 7898 12912
rect 14458 12900 14464 12912
rect 7892 12872 14464 12900
rect 7892 12860 7898 12872
rect 14458 12860 14464 12872
rect 14516 12860 14522 12912
rect 14734 12860 14740 12912
rect 14792 12900 14798 12912
rect 17782 12903 17840 12909
rect 17782 12900 17794 12903
rect 14792 12872 17794 12900
rect 14792 12860 14798 12872
rect 17782 12869 17794 12872
rect 17828 12869 17840 12903
rect 17782 12863 17840 12869
rect 18874 12860 18880 12912
rect 18932 12900 18938 12912
rect 20910 12903 20968 12909
rect 20910 12900 20922 12903
rect 18932 12872 20922 12900
rect 18932 12860 18938 12872
rect 20910 12869 20922 12872
rect 20956 12869 20968 12903
rect 20910 12863 20968 12869
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12832 2283 12835
rect 2314 12832 2320 12844
rect 2271 12804 2320 12832
rect 2271 12801 2283 12804
rect 2225 12795 2283 12801
rect 2314 12792 2320 12804
rect 2372 12792 2378 12844
rect 2406 12792 2412 12844
rect 2464 12832 2470 12844
rect 2869 12835 2927 12841
rect 2869 12832 2881 12835
rect 2464 12804 2881 12832
rect 2464 12792 2470 12804
rect 2869 12801 2881 12804
rect 2915 12801 2927 12835
rect 3326 12832 3332 12844
rect 3239 12804 3332 12832
rect 2869 12795 2927 12801
rect 3326 12792 3332 12804
rect 3384 12832 3390 12844
rect 5353 12835 5411 12841
rect 5353 12832 5365 12835
rect 3384 12804 5365 12832
rect 3384 12792 3390 12804
rect 5353 12801 5365 12804
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6733 12835 6791 12841
rect 6733 12832 6745 12835
rect 6328 12804 6745 12832
rect 6328 12792 6334 12804
rect 6733 12801 6745 12804
rect 6779 12801 6791 12835
rect 8018 12832 8024 12844
rect 7979 12804 8024 12832
rect 6733 12795 6791 12801
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 9033 12835 9091 12841
rect 9033 12832 9045 12835
rect 8628 12804 9045 12832
rect 8628 12792 8634 12804
rect 9033 12801 9045 12804
rect 9079 12832 9091 12835
rect 9214 12832 9220 12844
rect 9079 12804 9220 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9214 12792 9220 12804
rect 9272 12792 9278 12844
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12832 11207 12835
rect 11885 12835 11943 12841
rect 11885 12832 11897 12835
rect 11195 12804 11897 12832
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 11885 12801 11897 12804
rect 11931 12801 11943 12835
rect 13906 12832 13912 12844
rect 11885 12795 11943 12801
rect 12636 12804 13912 12832
rect 3050 12724 3056 12776
rect 3108 12764 3114 12776
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 3108 12736 3617 12764
rect 3108 12724 3114 12736
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 4430 12764 4436 12776
rect 4391 12736 4436 12764
rect 3605 12727 3663 12733
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 5166 12764 5172 12776
rect 5127 12736 5172 12764
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 6454 12764 6460 12776
rect 6415 12736 6460 12764
rect 6454 12724 6460 12736
rect 6512 12724 6518 12776
rect 6638 12764 6644 12776
rect 6599 12736 6644 12764
rect 6638 12724 6644 12736
rect 6696 12724 6702 12776
rect 8202 12764 8208 12776
rect 8163 12736 8208 12764
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12764 9367 12767
rect 9582 12764 9588 12776
rect 9355 12736 9588 12764
rect 9355 12733 9367 12736
rect 9309 12727 9367 12733
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 11974 12764 11980 12776
rect 10008 12736 10916 12764
rect 11935 12736 11980 12764
rect 10008 12724 10014 12736
rect 2593 12699 2651 12705
rect 2593 12665 2605 12699
rect 2639 12696 2651 12699
rect 5721 12699 5779 12705
rect 2639 12668 3556 12696
rect 2639 12665 2651 12668
rect 2593 12659 2651 12665
rect 3528 12640 3556 12668
rect 5721 12665 5733 12699
rect 5767 12696 5779 12699
rect 10778 12696 10784 12708
rect 5767 12668 8248 12696
rect 5767 12665 5779 12668
rect 5721 12659 5779 12665
rect 1854 12588 1860 12640
rect 1912 12628 1918 12640
rect 3142 12628 3148 12640
rect 1912 12600 3148 12628
rect 1912 12588 1918 12600
rect 3142 12588 3148 12600
rect 3200 12588 3206 12640
rect 3510 12588 3516 12640
rect 3568 12628 3574 12640
rect 7834 12628 7840 12640
rect 3568 12600 7840 12628
rect 3568 12588 3574 12600
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 8220 12628 8248 12668
rect 9646 12668 10784 12696
rect 9646 12628 9674 12668
rect 10778 12656 10784 12668
rect 10836 12656 10842 12708
rect 10888 12696 10916 12736
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 12161 12767 12219 12773
rect 12161 12733 12173 12767
rect 12207 12764 12219 12767
rect 12250 12764 12256 12776
rect 12207 12736 12256 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 12250 12724 12256 12736
rect 12308 12724 12314 12776
rect 12636 12696 12664 12804
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 14205 12835 14263 12841
rect 14205 12801 14217 12835
rect 14251 12832 14263 12835
rect 14550 12832 14556 12844
rect 14251 12804 14556 12832
rect 14251 12801 14263 12804
rect 14205 12795 14263 12801
rect 14550 12792 14556 12804
rect 14608 12832 14614 12844
rect 16942 12832 16948 12844
rect 14608 12804 16948 12832
rect 14608 12792 14614 12804
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 18046 12832 18052 12844
rect 18007 12804 18052 12832
rect 18046 12792 18052 12804
rect 18104 12832 18110 12844
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 18104 12804 18337 12832
rect 18104 12792 18110 12804
rect 18325 12801 18337 12804
rect 18371 12832 18383 12835
rect 18969 12835 19027 12841
rect 18969 12832 18981 12835
rect 18371 12804 18981 12832
rect 18371 12801 18383 12804
rect 18325 12795 18383 12801
rect 18969 12801 18981 12804
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 14461 12767 14519 12773
rect 14461 12733 14473 12767
rect 14507 12764 14519 12767
rect 14737 12767 14795 12773
rect 14737 12764 14749 12767
rect 14507 12736 14749 12764
rect 14507 12733 14519 12736
rect 14461 12727 14519 12733
rect 14737 12733 14749 12736
rect 14783 12733 14795 12767
rect 14737 12727 14795 12733
rect 21177 12767 21235 12773
rect 21177 12733 21189 12767
rect 21223 12764 21235 12767
rect 21266 12764 21272 12776
rect 21223 12736 21272 12764
rect 21223 12733 21235 12736
rect 21177 12727 21235 12733
rect 10888 12668 12664 12696
rect 12728 12668 13584 12696
rect 11514 12628 11520 12640
rect 8220 12600 9674 12628
rect 11475 12600 11520 12628
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 12158 12588 12164 12640
rect 12216 12628 12222 12640
rect 12728 12637 12756 12668
rect 12713 12631 12771 12637
rect 12713 12628 12725 12631
rect 12216 12600 12725 12628
rect 12216 12588 12222 12600
rect 12713 12597 12725 12600
rect 12759 12597 12771 12631
rect 12713 12591 12771 12597
rect 12894 12588 12900 12640
rect 12952 12628 12958 12640
rect 13081 12631 13139 12637
rect 13081 12628 13093 12631
rect 12952 12600 13093 12628
rect 12952 12588 12958 12600
rect 13081 12597 13093 12600
rect 13127 12597 13139 12631
rect 13556 12628 13584 12668
rect 13722 12628 13728 12640
rect 13556 12600 13728 12628
rect 13081 12591 13139 12597
rect 13722 12588 13728 12600
rect 13780 12628 13786 12640
rect 14476 12628 14504 12727
rect 21266 12724 21272 12736
rect 21324 12724 21330 12776
rect 13780 12600 14504 12628
rect 13780 12588 13786 12600
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 1578 12424 1584 12436
rect 1539 12396 1584 12424
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 3421 12427 3479 12433
rect 3421 12393 3433 12427
rect 3467 12424 3479 12427
rect 4154 12424 4160 12436
rect 3467 12396 4160 12424
rect 3467 12393 3479 12396
rect 3421 12387 3479 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 4525 12427 4583 12433
rect 4525 12393 4537 12427
rect 4571 12424 4583 12427
rect 5626 12424 5632 12436
rect 4571 12396 5632 12424
rect 4571 12393 4583 12396
rect 4525 12387 4583 12393
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 9214 12424 9220 12436
rect 7208 12396 9220 12424
rect 1596 12152 1624 12384
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 5537 12359 5595 12365
rect 4120 12328 5120 12356
rect 4120 12316 4126 12328
rect 2222 12288 2228 12300
rect 2183 12260 2228 12288
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12288 2927 12291
rect 3142 12288 3148 12300
rect 2915 12260 3148 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 3142 12248 3148 12260
rect 3200 12288 3206 12300
rect 3786 12288 3792 12300
rect 3200 12260 3792 12288
rect 3200 12248 3206 12260
rect 3786 12248 3792 12260
rect 3844 12248 3850 12300
rect 3973 12291 4031 12297
rect 3973 12257 3985 12291
rect 4019 12288 4031 12291
rect 4614 12288 4620 12300
rect 4019 12260 4620 12288
rect 4019 12257 4031 12260
rect 3973 12251 4031 12257
rect 4614 12248 4620 12260
rect 4672 12288 4678 12300
rect 4798 12288 4804 12300
rect 4672 12260 4804 12288
rect 4672 12248 4678 12260
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 4982 12288 4988 12300
rect 4943 12260 4988 12288
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 2406 12220 2412 12232
rect 2367 12192 2412 12220
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 3050 12220 3056 12232
rect 3011 12192 3056 12220
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4430 12220 4436 12232
rect 4203 12192 4436 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 4430 12180 4436 12192
rect 4488 12180 4494 12232
rect 5092 12220 5120 12328
rect 5537 12325 5549 12359
rect 5583 12356 5595 12359
rect 7208 12356 7236 12396
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 9766 12424 9772 12436
rect 9723 12396 9772 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 11057 12427 11115 12433
rect 11057 12393 11069 12427
rect 11103 12424 11115 12427
rect 11790 12424 11796 12436
rect 11103 12396 11796 12424
rect 11103 12393 11115 12396
rect 11057 12387 11115 12393
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12069 12427 12127 12433
rect 12069 12424 12081 12427
rect 12032 12396 12081 12424
rect 12032 12384 12038 12396
rect 12069 12393 12081 12396
rect 12115 12393 12127 12427
rect 12069 12387 12127 12393
rect 16390 12384 16396 12436
rect 16448 12424 16454 12436
rect 19242 12424 19248 12436
rect 16448 12396 19248 12424
rect 16448 12384 16454 12396
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 5583 12328 7236 12356
rect 7285 12359 7343 12365
rect 5583 12325 5595 12328
rect 5537 12319 5595 12325
rect 7285 12325 7297 12359
rect 7331 12356 7343 12359
rect 10686 12356 10692 12368
rect 7331 12328 8800 12356
rect 7331 12325 7343 12328
rect 7285 12319 7343 12325
rect 6270 12288 6276 12300
rect 6231 12260 6276 12288
rect 6270 12248 6276 12260
rect 6328 12248 6334 12300
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12288 6791 12291
rect 6779 12260 7972 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 5092 12192 5181 12220
rect 5169 12189 5181 12192
rect 5215 12189 5227 12223
rect 5169 12183 5227 12189
rect 2961 12155 3019 12161
rect 2961 12152 2973 12155
rect 1596 12124 2973 12152
rect 2961 12121 2973 12124
rect 3007 12121 3019 12155
rect 2961 12115 3019 12121
rect 3878 12112 3884 12164
rect 3936 12152 3942 12164
rect 6638 12152 6644 12164
rect 3936 12124 6644 12152
rect 3936 12112 3942 12124
rect 6638 12112 6644 12124
rect 6696 12112 6702 12164
rect 6825 12155 6883 12161
rect 6825 12121 6837 12155
rect 6871 12152 6883 12155
rect 7006 12152 7012 12164
rect 6871 12124 7012 12152
rect 6871 12121 6883 12124
rect 6825 12115 6883 12121
rect 7006 12112 7012 12124
rect 7064 12152 7070 12164
rect 7944 12152 7972 12260
rect 8018 12248 8024 12300
rect 8076 12288 8082 12300
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 8076 12260 8401 12288
rect 8076 12248 8082 12260
rect 8389 12257 8401 12260
rect 8435 12257 8447 12291
rect 8389 12251 8447 12257
rect 8772 12220 8800 12328
rect 9140 12328 10692 12356
rect 9140 12297 9168 12328
rect 10686 12316 10692 12328
rect 10744 12316 10750 12368
rect 9125 12291 9183 12297
rect 9125 12257 9137 12291
rect 9171 12257 9183 12291
rect 9125 12251 9183 12257
rect 11517 12291 11575 12297
rect 11517 12257 11529 12291
rect 11563 12257 11575 12291
rect 11517 12251 11575 12257
rect 11609 12291 11667 12297
rect 11609 12257 11621 12291
rect 11655 12288 11667 12291
rect 11790 12288 11796 12300
rect 11655 12260 11796 12288
rect 11655 12257 11667 12260
rect 11609 12251 11667 12257
rect 10318 12220 10324 12232
rect 8772 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 11532 12220 11560 12251
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 14458 12248 14464 12300
rect 14516 12288 14522 12300
rect 14642 12288 14648 12300
rect 14516 12260 14648 12288
rect 14516 12248 14522 12260
rect 14642 12248 14648 12260
rect 14700 12248 14706 12300
rect 12434 12220 12440 12232
rect 11532 12192 12440 12220
rect 12434 12180 12440 12192
rect 12492 12180 12498 12232
rect 13078 12180 13084 12232
rect 13136 12220 13142 12232
rect 13136 12192 13584 12220
rect 13136 12180 13142 12192
rect 12710 12152 12716 12164
rect 7064 12124 7788 12152
rect 7944 12124 12716 12152
rect 7064 12112 7070 12124
rect 3142 12044 3148 12096
rect 3200 12084 3206 12096
rect 4065 12087 4123 12093
rect 4065 12084 4077 12087
rect 3200 12056 4077 12084
rect 3200 12044 3206 12056
rect 4065 12053 4077 12056
rect 4111 12053 4123 12087
rect 5074 12084 5080 12096
rect 5035 12056 5080 12084
rect 4065 12047 4123 12053
rect 5074 12044 5080 12056
rect 5132 12044 5138 12096
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 6788 12056 6929 12084
rect 6788 12044 6794 12056
rect 6917 12053 6929 12056
rect 6963 12053 6975 12087
rect 7650 12084 7656 12096
rect 7611 12056 7656 12084
rect 6917 12047 6975 12053
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 7760 12084 7788 12124
rect 12710 12112 12716 12124
rect 12768 12112 12774 12164
rect 13446 12152 13452 12164
rect 13504 12161 13510 12164
rect 13416 12124 13452 12152
rect 13446 12112 13452 12124
rect 13504 12115 13516 12161
rect 13556 12152 13584 12192
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 14185 12223 14243 12229
rect 14185 12220 14197 12223
rect 13780 12192 14197 12220
rect 13780 12180 13786 12192
rect 14185 12189 14197 12192
rect 14231 12220 14243 12223
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 14231 12192 15025 12220
rect 14231 12189 14243 12192
rect 14185 12183 14243 12189
rect 15013 12189 15025 12192
rect 15059 12220 15071 12223
rect 16114 12220 16120 12232
rect 15059 12192 16120 12220
rect 15059 12189 15071 12192
rect 15013 12183 15071 12189
rect 16114 12180 16120 12192
rect 16172 12220 16178 12232
rect 16669 12223 16727 12229
rect 16669 12220 16681 12223
rect 16172 12192 16681 12220
rect 16172 12180 16178 12192
rect 16669 12189 16681 12192
rect 16715 12220 16727 12223
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 16715 12192 17141 12220
rect 16715 12189 16727 12192
rect 16669 12183 16727 12189
rect 17129 12189 17141 12192
rect 17175 12220 17187 12223
rect 18785 12223 18843 12229
rect 18785 12220 18797 12223
rect 17175 12192 18797 12220
rect 17175 12189 17187 12192
rect 17129 12183 17187 12189
rect 18785 12189 18797 12192
rect 18831 12220 18843 12223
rect 19058 12220 19064 12232
rect 18831 12192 19064 12220
rect 18831 12189 18843 12192
rect 18785 12183 18843 12189
rect 19058 12180 19064 12192
rect 19116 12220 19122 12232
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 19116 12192 19257 12220
rect 19116 12180 19122 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 21361 12223 21419 12229
rect 21361 12220 21373 12223
rect 21324 12192 21373 12220
rect 21324 12180 21330 12192
rect 21361 12189 21373 12192
rect 21407 12189 21419 12223
rect 21361 12183 21419 12189
rect 15286 12161 15292 12164
rect 15280 12152 15292 12161
rect 13556 12124 14596 12152
rect 15247 12124 15292 12152
rect 13504 12112 13510 12115
rect 8021 12087 8079 12093
rect 8021 12084 8033 12087
rect 7760 12056 8033 12084
rect 8021 12053 8033 12056
rect 8067 12053 8079 12087
rect 8021 12047 8079 12053
rect 8110 12044 8116 12096
rect 8168 12084 8174 12096
rect 9217 12087 9275 12093
rect 9217 12084 9229 12087
rect 8168 12056 9229 12084
rect 8168 12044 8174 12056
rect 9217 12053 9229 12056
rect 9263 12053 9275 12087
rect 9217 12047 9275 12053
rect 9306 12044 9312 12096
rect 9364 12084 9370 12096
rect 9364 12056 9409 12084
rect 9364 12044 9370 12056
rect 9950 12044 9956 12096
rect 10008 12084 10014 12096
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 10008 12056 10609 12084
rect 10008 12044 10014 12056
rect 10597 12053 10609 12056
rect 10643 12084 10655 12087
rect 11698 12084 11704 12096
rect 10643 12056 11704 12084
rect 10643 12053 10655 12056
rect 10597 12047 10655 12053
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 12158 12044 12164 12096
rect 12216 12084 12222 12096
rect 12345 12087 12403 12093
rect 12345 12084 12357 12087
rect 12216 12056 12357 12084
rect 12216 12044 12222 12056
rect 12345 12053 12357 12056
rect 12391 12053 12403 12087
rect 13464 12084 13492 12112
rect 14458 12084 14464 12096
rect 13464 12056 14464 12084
rect 12345 12047 12403 12053
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 14568 12084 14596 12124
rect 15280 12115 15292 12124
rect 15286 12112 15292 12115
rect 15344 12112 15350 12164
rect 17374 12155 17432 12161
rect 17374 12152 17386 12155
rect 16546 12124 17386 12152
rect 16393 12087 16451 12093
rect 16393 12084 16405 12087
rect 14568 12056 16405 12084
rect 16393 12053 16405 12056
rect 16439 12084 16451 12087
rect 16546 12084 16574 12124
rect 17374 12121 17386 12124
rect 17420 12121 17432 12155
rect 21082 12152 21088 12164
rect 21140 12161 21146 12164
rect 17374 12115 17432 12121
rect 18524 12124 21088 12152
rect 18524 12096 18552 12124
rect 21082 12112 21088 12124
rect 21140 12115 21152 12161
rect 21140 12112 21146 12115
rect 18506 12084 18512 12096
rect 16439 12056 16574 12084
rect 18467 12056 18512 12084
rect 16439 12053 16451 12056
rect 16393 12047 16451 12053
rect 18506 12044 18512 12056
rect 18564 12044 18570 12096
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 18932 12056 19625 12084
rect 18932 12044 18938 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 19613 12047 19671 12053
rect 19981 12087 20039 12093
rect 19981 12053 19993 12087
rect 20027 12084 20039 12087
rect 20438 12084 20444 12096
rect 20027 12056 20444 12084
rect 20027 12053 20039 12056
rect 19981 12047 20039 12053
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 2041 11883 2099 11889
rect 2041 11849 2053 11883
rect 2087 11880 2099 11883
rect 2958 11880 2964 11892
rect 2087 11852 2964 11880
rect 2087 11849 2099 11852
rect 2041 11843 2099 11849
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 3142 11880 3148 11892
rect 3103 11852 3148 11880
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 3605 11883 3663 11889
rect 3605 11849 3617 11883
rect 3651 11880 3663 11883
rect 3970 11880 3976 11892
rect 3651 11852 3976 11880
rect 3651 11849 3663 11852
rect 3605 11843 3663 11849
rect 382 11772 388 11824
rect 440 11812 446 11824
rect 2593 11815 2651 11821
rect 2593 11812 2605 11815
rect 440 11784 2605 11812
rect 440 11772 446 11784
rect 2593 11781 2605 11784
rect 2639 11812 2651 11815
rect 3620 11812 3648 11843
rect 3970 11840 3976 11852
rect 4028 11880 4034 11892
rect 5074 11880 5080 11892
rect 4028 11852 5080 11880
rect 4028 11840 4034 11852
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 6638 11840 6644 11892
rect 6696 11880 6702 11892
rect 6917 11883 6975 11889
rect 6917 11880 6929 11883
rect 6696 11852 6929 11880
rect 6696 11840 6702 11852
rect 6917 11849 6929 11852
rect 6963 11849 6975 11883
rect 6917 11843 6975 11849
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 9217 11883 9275 11889
rect 7248 11852 9168 11880
rect 7248 11840 7254 11852
rect 7282 11812 7288 11824
rect 2639 11784 3648 11812
rect 4724 11784 7288 11812
rect 2639 11781 2651 11784
rect 2593 11775 2651 11781
rect 4724 11753 4752 11784
rect 7282 11772 7288 11784
rect 7340 11772 7346 11824
rect 9140 11812 9168 11852
rect 9217 11849 9229 11883
rect 9263 11880 9275 11883
rect 9306 11880 9312 11892
rect 9263 11852 9312 11880
rect 9263 11849 9275 11852
rect 9217 11843 9275 11849
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 10870 11880 10876 11892
rect 10831 11852 10876 11880
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 19610 11880 19616 11892
rect 13556 11852 14228 11880
rect 19571 11852 19616 11880
rect 9950 11812 9956 11824
rect 9140 11784 9956 11812
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 10042 11772 10048 11824
rect 10100 11812 10106 11824
rect 13556 11812 13584 11852
rect 13722 11812 13728 11824
rect 10100 11784 13584 11812
rect 13683 11784 13728 11812
rect 10100 11772 10106 11784
rect 13722 11772 13728 11784
rect 13780 11812 13786 11824
rect 14093 11815 14151 11821
rect 14093 11812 14105 11815
rect 13780 11784 14105 11812
rect 13780 11772 13786 11784
rect 14093 11781 14105 11784
rect 14139 11781 14151 11815
rect 14200 11812 14228 11852
rect 19610 11840 19616 11852
rect 19668 11840 19674 11892
rect 21082 11840 21088 11892
rect 21140 11880 21146 11892
rect 21269 11883 21327 11889
rect 21269 11880 21281 11883
rect 21140 11852 21281 11880
rect 21140 11840 21146 11852
rect 21269 11849 21281 11852
rect 21315 11849 21327 11883
rect 21269 11843 21327 11849
rect 14798 11815 14856 11821
rect 14798 11812 14810 11815
rect 14200 11784 14810 11812
rect 14093 11775 14151 11781
rect 14798 11781 14810 11784
rect 14844 11812 14856 11815
rect 15746 11812 15752 11824
rect 14844 11784 15752 11812
rect 14844 11781 14856 11784
rect 14798 11775 14856 11781
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 2271 11716 4445 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 4433 11713 4445 11716
rect 4479 11713 4491 11747
rect 4433 11707 4491 11713
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 5353 11747 5411 11753
rect 5353 11713 5365 11747
rect 5399 11744 5411 11747
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 5399 11716 6377 11744
rect 5399 11713 5411 11716
rect 5353 11707 5411 11713
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11744 7711 11747
rect 7834 11744 7840 11756
rect 7699 11716 7840 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 2314 11636 2320 11688
rect 2372 11676 2378 11688
rect 2372 11648 2774 11676
rect 2372 11636 2378 11648
rect 2746 11608 2774 11648
rect 3142 11636 3148 11688
rect 3200 11676 3206 11688
rect 4522 11676 4528 11688
rect 3200 11648 4528 11676
rect 3200 11636 3206 11648
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 5442 11676 5448 11688
rect 5403 11648 5448 11676
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11676 5687 11679
rect 7668 11676 7696 11707
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 10781 11747 10839 11753
rect 10781 11713 10793 11747
rect 10827 11744 10839 11747
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 10827 11716 11529 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 12710 11704 12716 11756
rect 12768 11744 12774 11756
rect 13182 11747 13240 11753
rect 13182 11744 13194 11747
rect 12768 11716 13194 11744
rect 12768 11704 12774 11716
rect 13182 11713 13194 11716
rect 13228 11744 13240 11747
rect 13354 11744 13360 11756
rect 13228 11716 13360 11744
rect 13228 11713 13240 11716
rect 13182 11707 13240 11713
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11744 13507 11747
rect 13740 11744 13768 11772
rect 13495 11716 13768 11744
rect 14108 11744 14136 11775
rect 15746 11772 15752 11784
rect 15804 11772 15810 11824
rect 17218 11772 17224 11824
rect 17276 11772 17282 11824
rect 18782 11772 18788 11824
rect 18840 11821 18846 11824
rect 18840 11812 18852 11821
rect 18840 11784 18885 11812
rect 19076 11784 21036 11812
rect 18840 11775 18852 11784
rect 18840 11772 18846 11775
rect 14553 11747 14611 11753
rect 14553 11744 14565 11747
rect 14108 11716 14565 11744
rect 13495 11713 13507 11716
rect 13449 11707 13507 11713
rect 14553 11713 14565 11716
rect 14599 11713 14611 11747
rect 14553 11707 14611 11713
rect 15102 11704 15108 11756
rect 15160 11744 15166 11756
rect 16298 11744 16304 11756
rect 15160 11716 16304 11744
rect 15160 11704 15166 11716
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 17236 11744 17264 11772
rect 19076 11756 19104 11784
rect 19058 11744 19064 11756
rect 17236 11716 17356 11744
rect 19019 11716 19064 11744
rect 10042 11676 10048 11688
rect 5675 11648 7696 11676
rect 10003 11648 10048 11676
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 12342 11676 12348 11688
rect 11103 11648 12348 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 12342 11636 12348 11648
rect 12400 11636 12406 11688
rect 16114 11636 16120 11688
rect 16172 11676 16178 11688
rect 16761 11679 16819 11685
rect 16761 11676 16773 11679
rect 16172 11648 16773 11676
rect 16172 11636 16178 11648
rect 16761 11645 16773 11648
rect 16807 11676 16819 11679
rect 17221 11679 17279 11685
rect 17221 11676 17233 11679
rect 16807 11648 17233 11676
rect 16807 11645 16819 11648
rect 16761 11639 16819 11645
rect 17221 11645 17233 11648
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 10413 11611 10471 11617
rect 10413 11608 10425 11611
rect 2746 11580 10425 11608
rect 10413 11577 10425 11580
rect 10459 11577 10471 11611
rect 10413 11571 10471 11577
rect 15933 11611 15991 11617
rect 15933 11577 15945 11611
rect 15979 11608 15991 11611
rect 17328 11608 17356 11716
rect 19058 11704 19064 11716
rect 19116 11704 19122 11756
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 21008 11753 21036 11784
rect 20726 11747 20784 11753
rect 20726 11744 20738 11747
rect 20496 11716 20738 11744
rect 20496 11704 20502 11716
rect 20726 11713 20738 11716
rect 20772 11713 20784 11747
rect 20726 11707 20784 11713
rect 20993 11747 21051 11753
rect 20993 11713 21005 11747
rect 21039 11744 21051 11747
rect 21266 11744 21272 11756
rect 21039 11716 21272 11744
rect 21039 11713 21051 11716
rect 20993 11707 21051 11713
rect 21266 11704 21272 11716
rect 21324 11704 21330 11756
rect 15979 11580 17356 11608
rect 15979 11577 15991 11580
rect 15933 11571 15991 11577
rect 3050 11500 3056 11552
rect 3108 11540 3114 11552
rect 3881 11543 3939 11549
rect 3881 11540 3893 11543
rect 3108 11512 3893 11540
rect 3108 11500 3114 11512
rect 3881 11509 3893 11512
rect 3927 11540 3939 11543
rect 4062 11540 4068 11552
rect 3927 11512 4068 11540
rect 3927 11509 3939 11512
rect 3881 11503 3939 11509
rect 4062 11500 4068 11512
rect 4120 11500 4126 11552
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4985 11543 5043 11549
rect 4985 11540 4997 11543
rect 4304 11512 4997 11540
rect 4304 11500 4310 11512
rect 4985 11509 4997 11512
rect 5031 11509 5043 11543
rect 4985 11503 5043 11509
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 6730 11540 6736 11552
rect 5960 11512 6736 11540
rect 5960 11500 5966 11512
rect 6730 11500 6736 11512
rect 6788 11540 6794 11552
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 6788 11512 7205 11540
rect 6788 11500 6794 11512
rect 7193 11509 7205 11512
rect 7239 11509 7251 11543
rect 12066 11540 12072 11552
rect 12027 11512 12072 11540
rect 7193 11503 7251 11509
rect 12066 11500 12072 11512
rect 12124 11540 12130 11552
rect 14734 11540 14740 11552
rect 12124 11512 14740 11540
rect 12124 11500 12130 11512
rect 14734 11500 14740 11512
rect 14792 11500 14798 11552
rect 16114 11500 16120 11552
rect 16172 11540 16178 11552
rect 16209 11543 16267 11549
rect 16209 11540 16221 11543
rect 16172 11512 16221 11540
rect 16172 11500 16178 11512
rect 16209 11509 16221 11512
rect 16255 11509 16267 11543
rect 16209 11503 16267 11509
rect 16298 11500 16304 11552
rect 16356 11540 16362 11552
rect 17681 11543 17739 11549
rect 17681 11540 17693 11543
rect 16356 11512 17693 11540
rect 16356 11500 16362 11512
rect 17681 11509 17693 11512
rect 17727 11540 17739 11543
rect 18414 11540 18420 11552
rect 17727 11512 18420 11540
rect 17727 11509 17739 11512
rect 17681 11503 17739 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 2041 11339 2099 11345
rect 2041 11305 2053 11339
rect 2087 11336 2099 11339
rect 2774 11336 2780 11348
rect 2087 11308 2780 11336
rect 2087 11305 2099 11308
rect 2041 11299 2099 11305
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 3053 11339 3111 11345
rect 3053 11305 3065 11339
rect 3099 11336 3111 11339
rect 4430 11336 4436 11348
rect 3099 11308 4436 11336
rect 3099 11305 3111 11308
rect 3053 11299 3111 11305
rect 4430 11296 4436 11308
rect 4488 11336 4494 11348
rect 5166 11336 5172 11348
rect 4488 11308 5172 11336
rect 4488 11296 4494 11308
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 5537 11339 5595 11345
rect 5537 11336 5549 11339
rect 5500 11308 5549 11336
rect 5500 11296 5506 11308
rect 5537 11305 5549 11308
rect 5583 11305 5595 11339
rect 5537 11299 5595 11305
rect 6733 11339 6791 11345
rect 6733 11305 6745 11339
rect 6779 11336 6791 11339
rect 8110 11336 8116 11348
rect 6779 11308 8116 11336
rect 6779 11305 6791 11308
rect 6733 11299 6791 11305
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8720 11308 8953 11336
rect 8720 11296 8726 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 13446 11336 13452 11348
rect 8941 11299 8999 11305
rect 9048 11308 13452 11336
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 9048 11268 9076 11308
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 14826 11296 14832 11348
rect 14884 11336 14890 11348
rect 14884 11308 15056 11336
rect 14884 11296 14890 11308
rect 11241 11271 11299 11277
rect 11241 11268 11253 11271
rect 4212 11240 6316 11268
rect 4212 11228 4218 11240
rect 1486 11160 1492 11212
rect 1544 11200 1550 11212
rect 3973 11203 4031 11209
rect 3973 11200 3985 11203
rect 1544 11172 3985 11200
rect 1544 11160 1550 11172
rect 3973 11169 3985 11172
rect 4019 11169 4031 11203
rect 3973 11163 4031 11169
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11200 5043 11203
rect 5626 11200 5632 11212
rect 5031 11172 5632 11200
rect 5031 11169 5043 11172
rect 4985 11163 5043 11169
rect 5626 11160 5632 11172
rect 5684 11200 5690 11212
rect 6178 11200 6184 11212
rect 5684 11172 6040 11200
rect 6139 11172 6184 11200
rect 5684 11160 5690 11172
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 4062 11132 4068 11144
rect 2271 11104 4068 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 4246 11132 4252 11144
rect 4207 11104 4252 11132
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 5077 11135 5135 11141
rect 5077 11132 5089 11135
rect 4396 11104 5089 11132
rect 4396 11092 4402 11104
rect 5077 11101 5089 11104
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5166 11092 5172 11144
rect 5224 11132 5230 11144
rect 6012 11132 6040 11172
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6288 11209 6316 11240
rect 6380 11240 9076 11268
rect 10704 11240 11253 11268
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11169 6331 11203
rect 6273 11163 6331 11169
rect 6380 11132 6408 11240
rect 6730 11160 6736 11212
rect 6788 11200 6794 11212
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 6788 11172 7757 11200
rect 6788 11160 6794 11172
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 9490 11200 9496 11212
rect 9451 11172 9496 11200
rect 7745 11163 7803 11169
rect 9490 11160 9496 11172
rect 9548 11160 9554 11212
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 10704 11209 10732 11240
rect 11241 11237 11253 11240
rect 11287 11237 11299 11271
rect 12342 11268 12348 11280
rect 12303 11240 12348 11268
rect 11241 11231 11299 11237
rect 12342 11228 12348 11240
rect 12400 11228 12406 11280
rect 15028 11268 15056 11308
rect 15194 11296 15200 11348
rect 15252 11336 15258 11348
rect 15470 11336 15476 11348
rect 15252 11308 15476 11336
rect 15252 11296 15258 11308
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 15580 11308 17417 11336
rect 15580 11268 15608 11308
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 17405 11299 17463 11305
rect 18782 11296 18788 11348
rect 18840 11336 18846 11348
rect 19610 11336 19616 11348
rect 18840 11308 19616 11336
rect 18840 11296 18846 11308
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 20806 11296 20812 11348
rect 20864 11336 20870 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20864 11308 21005 11336
rect 20864 11296 20870 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 21266 11336 21272 11348
rect 21227 11308 21272 11336
rect 20993 11299 21051 11305
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 15746 11268 15752 11280
rect 15028 11240 15608 11268
rect 15707 11240 15752 11268
rect 15746 11228 15752 11240
rect 15804 11228 15810 11280
rect 10689 11203 10747 11209
rect 10689 11200 10701 11203
rect 10192 11172 10701 11200
rect 10192 11160 10198 11172
rect 10689 11169 10701 11172
rect 10735 11169 10747 11203
rect 10689 11163 10747 11169
rect 10873 11203 10931 11209
rect 10873 11169 10885 11203
rect 10919 11200 10931 11203
rect 12710 11200 12716 11212
rect 10919 11172 12716 11200
rect 10919 11169 10931 11172
rect 10873 11163 10931 11169
rect 12710 11160 12716 11172
rect 12768 11160 12774 11212
rect 13722 11200 13728 11212
rect 13683 11172 13728 11200
rect 13722 11160 13728 11172
rect 13780 11200 13786 11212
rect 14093 11203 14151 11209
rect 14093 11200 14105 11203
rect 13780 11172 14105 11200
rect 13780 11160 13786 11172
rect 14093 11169 14105 11172
rect 14139 11169 14151 11203
rect 14093 11163 14151 11169
rect 19058 11160 19064 11212
rect 19116 11200 19122 11212
rect 19613 11203 19671 11209
rect 19613 11200 19625 11203
rect 19116 11172 19625 11200
rect 19116 11160 19122 11172
rect 19613 11169 19625 11172
rect 19659 11169 19671 11203
rect 19613 11163 19671 11169
rect 7466 11132 7472 11144
rect 5224 11104 5269 11132
rect 6012 11104 6408 11132
rect 7427 11104 7472 11132
rect 5224 11092 5230 11104
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9180 11104 9536 11132
rect 9180 11092 9186 11104
rect 9508 11076 9536 11104
rect 10042 11092 10048 11144
rect 10100 11132 10106 11144
rect 10597 11135 10655 11141
rect 10597 11132 10609 11135
rect 10100 11104 10609 11132
rect 10100 11092 10106 11104
rect 10597 11101 10609 11104
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 14366 11141 14372 11144
rect 13458 11135 13516 11141
rect 13458 11132 13470 11135
rect 13228 11104 13470 11132
rect 13228 11092 13234 11104
rect 13458 11101 13470 11104
rect 13504 11132 13516 11135
rect 13504 11104 14320 11132
rect 13504 11101 13516 11104
rect 13458 11095 13516 11101
rect 14292 11076 14320 11104
rect 14360 11095 14372 11141
rect 14424 11132 14430 11144
rect 14424 11104 14460 11132
rect 14366 11092 14372 11095
rect 14424 11092 14430 11104
rect 16114 11092 16120 11144
rect 16172 11132 16178 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 16172 11104 17141 11132
rect 16172 11092 16178 11104
rect 17129 11101 17141 11104
rect 17175 11132 17187 11135
rect 18785 11135 18843 11141
rect 18785 11132 18797 11135
rect 17175 11104 18797 11132
rect 17175 11101 17187 11104
rect 17129 11095 17187 11101
rect 18785 11101 18797 11104
rect 18831 11101 18843 11135
rect 18785 11095 18843 11101
rect 19518 11092 19524 11144
rect 19576 11132 19582 11144
rect 19869 11135 19927 11141
rect 19869 11132 19881 11135
rect 19576 11104 19881 11132
rect 19576 11092 19582 11104
rect 19869 11101 19881 11104
rect 19915 11101 19927 11135
rect 19869 11095 19927 11101
rect 3421 11067 3479 11073
rect 3421 11033 3433 11067
rect 3467 11064 3479 11067
rect 3510 11064 3516 11076
rect 3467 11036 3516 11064
rect 3467 11033 3479 11036
rect 3421 11027 3479 11033
rect 3510 11024 3516 11036
rect 3568 11024 3574 11076
rect 4982 11024 4988 11076
rect 5040 11064 5046 11076
rect 7193 11067 7251 11073
rect 7193 11064 7205 11067
rect 5040 11036 7205 11064
rect 5040 11024 5046 11036
rect 7193 11033 7205 11036
rect 7239 11033 7251 11067
rect 7193 11027 7251 11033
rect 8573 11067 8631 11073
rect 8573 11033 8585 11067
rect 8619 11064 8631 11067
rect 9309 11067 9367 11073
rect 9309 11064 9321 11067
rect 8619 11036 9321 11064
rect 8619 11033 8631 11036
rect 8573 11027 8631 11033
rect 9309 11033 9321 11036
rect 9355 11033 9367 11067
rect 9309 11027 9367 11033
rect 9490 11024 9496 11076
rect 9548 11024 9554 11076
rect 12268 11036 12480 11064
rect 5810 10956 5816 11008
rect 5868 10996 5874 11008
rect 6365 10999 6423 11005
rect 6365 10996 6377 10999
rect 5868 10968 6377 10996
rect 5868 10956 5874 10968
rect 6365 10965 6377 10968
rect 6411 10965 6423 10999
rect 6365 10959 6423 10965
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 9401 10999 9459 11005
rect 9401 10996 9413 10999
rect 9180 10968 9413 10996
rect 9180 10956 9186 10968
rect 9401 10965 9413 10968
rect 9447 10965 9459 10999
rect 10226 10996 10232 11008
rect 10187 10968 10232 10996
rect 9401 10959 9459 10965
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 10318 10956 10324 11008
rect 10376 10996 10382 11008
rect 12268 10996 12296 11036
rect 10376 10968 12296 10996
rect 12452 10996 12480 11036
rect 14274 11024 14280 11076
rect 14332 11024 14338 11076
rect 16884 11067 16942 11073
rect 15672 11036 15884 11064
rect 15672 10996 15700 11036
rect 12452 10968 15700 10996
rect 15856 10996 15884 11036
rect 16884 11033 16896 11067
rect 16930 11064 16942 11067
rect 17034 11064 17040 11076
rect 16930 11036 17040 11064
rect 16930 11033 16942 11036
rect 16884 11027 16942 11033
rect 17034 11024 17040 11036
rect 17092 11024 17098 11076
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 18540 11067 18598 11073
rect 18540 11064 18552 11067
rect 17368 11036 18552 11064
rect 17368 11024 17374 11036
rect 18540 11033 18552 11036
rect 18586 11064 18598 11067
rect 19245 11067 19303 11073
rect 19245 11064 19257 11067
rect 18586 11036 19257 11064
rect 18586 11033 18598 11036
rect 18540 11027 18598 11033
rect 19245 11033 19257 11036
rect 19291 11033 19303 11067
rect 19245 11027 19303 11033
rect 18322 10996 18328 11008
rect 15856 10968 18328 10996
rect 10376 10956 10382 10968
rect 18322 10956 18328 10968
rect 18380 10956 18386 11008
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 2041 10795 2099 10801
rect 2041 10792 2053 10795
rect 1820 10764 2053 10792
rect 1820 10752 1826 10764
rect 2041 10761 2053 10764
rect 2087 10761 2099 10795
rect 2041 10755 2099 10761
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4338 10792 4344 10804
rect 4019 10764 4344 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 4614 10792 4620 10804
rect 4575 10764 4620 10792
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 6730 10792 6736 10804
rect 6691 10764 6736 10792
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 7101 10795 7159 10801
rect 7101 10761 7113 10795
rect 7147 10792 7159 10795
rect 7745 10795 7803 10801
rect 7745 10792 7757 10795
rect 7147 10764 7757 10792
rect 7147 10761 7159 10764
rect 7101 10755 7159 10761
rect 7745 10761 7757 10764
rect 7791 10761 7803 10795
rect 7745 10755 7803 10761
rect 7837 10795 7895 10801
rect 7837 10761 7849 10795
rect 7883 10792 7895 10795
rect 9766 10792 9772 10804
rect 7883 10764 9772 10792
rect 7883 10761 7895 10764
rect 7837 10755 7895 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 10284 10764 10333 10792
rect 10284 10752 10290 10764
rect 10321 10761 10333 10764
rect 10367 10761 10379 10795
rect 12986 10792 12992 10804
rect 12947 10764 12992 10792
rect 10321 10755 10379 10761
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 15378 10792 15384 10804
rect 13188 10764 15384 10792
rect 2593 10727 2651 10733
rect 2593 10693 2605 10727
rect 2639 10724 2651 10727
rect 2682 10724 2688 10736
rect 2639 10696 2688 10724
rect 2639 10693 2651 10696
rect 2593 10687 2651 10693
rect 2682 10684 2688 10696
rect 2740 10684 2746 10736
rect 4062 10684 4068 10736
rect 4120 10724 4126 10736
rect 5721 10727 5779 10733
rect 5721 10724 5733 10727
rect 4120 10696 5733 10724
rect 4120 10684 4126 10696
rect 5721 10693 5733 10696
rect 5767 10693 5779 10727
rect 6641 10727 6699 10733
rect 6641 10724 6653 10727
rect 5721 10687 5779 10693
rect 5828 10696 6653 10724
rect 1486 10616 1492 10668
rect 1544 10656 1550 10668
rect 1857 10659 1915 10665
rect 1857 10656 1869 10659
rect 1544 10628 1869 10656
rect 1544 10616 1550 10628
rect 1857 10625 1869 10628
rect 1903 10625 1915 10659
rect 2866 10656 2872 10668
rect 2827 10628 2872 10656
rect 1857 10619 1915 10625
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 3602 10656 3608 10668
rect 3563 10628 3608 10656
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4249 10659 4307 10665
rect 4249 10656 4261 10659
rect 4212 10628 4261 10656
rect 4212 10616 4218 10628
rect 4249 10625 4261 10628
rect 4295 10625 4307 10659
rect 4249 10619 4307 10625
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10656 5319 10659
rect 5828 10656 5856 10696
rect 6641 10693 6653 10696
rect 6687 10724 6699 10727
rect 7006 10724 7012 10736
rect 6687 10696 7012 10724
rect 6687 10693 6699 10696
rect 6641 10687 6699 10693
rect 7006 10684 7012 10696
rect 7064 10684 7070 10736
rect 8478 10684 8484 10736
rect 8536 10724 8542 10736
rect 8665 10727 8723 10733
rect 8665 10724 8677 10727
rect 8536 10696 8677 10724
rect 8536 10684 8542 10696
rect 8665 10693 8677 10696
rect 8711 10724 8723 10727
rect 13188 10724 13216 10764
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 19702 10792 19708 10804
rect 19663 10764 19708 10792
rect 19702 10752 19708 10764
rect 19760 10752 19766 10804
rect 19981 10795 20039 10801
rect 19981 10761 19993 10795
rect 20027 10792 20039 10795
rect 20070 10792 20076 10804
rect 20027 10764 20076 10792
rect 20027 10761 20039 10764
rect 19981 10755 20039 10761
rect 20070 10752 20076 10764
rect 20128 10752 20134 10804
rect 8711 10696 13216 10724
rect 13740 10696 14412 10724
rect 8711 10693 8723 10696
rect 8665 10687 8723 10693
rect 5307 10628 5856 10656
rect 5997 10659 6055 10665
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 5997 10625 6009 10659
rect 6043 10656 6055 10659
rect 8386 10656 8392 10668
rect 6043 10628 8392 10656
rect 6043 10625 6055 10628
rect 5997 10619 6055 10625
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10656 10287 10659
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10275 10628 10885 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 12621 10659 12679 10665
rect 12621 10625 12633 10659
rect 12667 10656 12679 10659
rect 13740 10656 13768 10696
rect 12667 10628 13768 10656
rect 12667 10625 12679 10628
rect 12621 10619 12679 10625
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 14102 10659 14160 10665
rect 14102 10656 14114 10659
rect 13872 10628 14114 10656
rect 13872 10616 13878 10628
rect 14102 10625 14114 10628
rect 14148 10625 14160 10659
rect 14102 10619 14160 10625
rect 14274 10616 14280 10668
rect 14332 10616 14338 10668
rect 14384 10665 14412 10696
rect 14734 10684 14740 10736
rect 14792 10724 14798 10736
rect 15758 10727 15816 10733
rect 15758 10724 15770 10727
rect 14792 10696 15770 10724
rect 14792 10684 14798 10696
rect 15758 10693 15770 10696
rect 15804 10693 15816 10727
rect 15758 10687 15816 10693
rect 16684 10696 18368 10724
rect 16684 10665 16712 10696
rect 14369 10659 14427 10665
rect 14369 10625 14381 10659
rect 14415 10656 14427 10659
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 14415 10628 16068 10656
rect 14415 10625 14427 10628
rect 14369 10619 14427 10625
rect 2498 10548 2504 10600
rect 2556 10588 2562 10600
rect 3329 10591 3387 10597
rect 3329 10588 3341 10591
rect 2556 10560 3341 10588
rect 2556 10548 2562 10560
rect 3329 10557 3341 10560
rect 3375 10557 3387 10591
rect 3329 10551 3387 10557
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 8018 10588 8024 10600
rect 6604 10560 6649 10588
rect 7979 10560 8024 10588
rect 6604 10548 6610 10560
rect 8018 10548 8024 10560
rect 8076 10548 8082 10600
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 9306 10588 9312 10600
rect 9171 10560 9312 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10588 10563 10591
rect 12066 10588 12072 10600
rect 10551 10560 12072 10588
rect 10551 10557 10563 10560
rect 10505 10551 10563 10557
rect 12066 10548 12072 10560
rect 12124 10548 12130 10600
rect 14292 10588 14320 10616
rect 16040 10597 16068 10628
rect 16546 10628 16681 10656
rect 16025 10591 16083 10597
rect 14292 10560 14688 10588
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 14660 10529 14688 10560
rect 16025 10557 16037 10591
rect 16071 10588 16083 10591
rect 16114 10588 16120 10600
rect 16071 10560 16120 10588
rect 16071 10557 16083 10560
rect 16025 10551 16083 10557
rect 16114 10548 16120 10560
rect 16172 10588 16178 10600
rect 16546 10588 16574 10628
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 16936 10659 16994 10665
rect 16936 10625 16948 10659
rect 16982 10656 16994 10659
rect 17218 10656 17224 10668
rect 16982 10628 17224 10656
rect 16982 10625 16994 10628
rect 16936 10619 16994 10625
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 18340 10665 18368 10696
rect 18414 10684 18420 10736
rect 18472 10724 18478 10736
rect 18570 10727 18628 10733
rect 18570 10724 18582 10727
rect 18472 10696 18582 10724
rect 18472 10684 18478 10696
rect 18570 10693 18582 10696
rect 18616 10693 18628 10727
rect 18570 10687 18628 10693
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10625 18383 10659
rect 18325 10619 18383 10625
rect 21082 10616 21088 10668
rect 21140 10665 21146 10668
rect 21140 10656 21152 10665
rect 21140 10628 21185 10656
rect 21140 10619 21152 10628
rect 21140 10616 21146 10619
rect 21266 10616 21272 10668
rect 21324 10656 21330 10668
rect 21361 10659 21419 10665
rect 21361 10656 21373 10659
rect 21324 10628 21373 10656
rect 21324 10616 21330 10628
rect 21361 10625 21373 10628
rect 21407 10625 21419 10659
rect 21361 10619 21419 10625
rect 16172 10560 16574 10588
rect 16172 10548 16178 10560
rect 9861 10523 9919 10529
rect 9861 10520 9873 10523
rect 6788 10492 9873 10520
rect 6788 10480 6794 10492
rect 9861 10489 9873 10492
rect 9907 10489 9919 10523
rect 9861 10483 9919 10489
rect 14645 10523 14703 10529
rect 14645 10489 14657 10523
rect 14691 10489 14703 10523
rect 14645 10483 14703 10489
rect 1486 10452 1492 10464
rect 1447 10424 1492 10452
rect 1486 10412 1492 10424
rect 1544 10412 1550 10464
rect 7282 10412 7288 10464
rect 7340 10452 7346 10464
rect 7377 10455 7435 10461
rect 7377 10452 7389 10455
rect 7340 10424 7389 10452
rect 7340 10412 7346 10424
rect 7377 10421 7389 10424
rect 7423 10421 7435 10455
rect 7377 10415 7435 10421
rect 9122 10412 9128 10464
rect 9180 10452 9186 10464
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9180 10424 9413 10452
rect 9180 10412 9186 10424
rect 9401 10421 9413 10424
rect 9447 10421 9459 10455
rect 9401 10415 9459 10421
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 15286 10452 15292 10464
rect 10008 10424 15292 10452
rect 10008 10412 10014 10424
rect 15286 10412 15292 10424
rect 15344 10452 15350 10464
rect 15746 10452 15752 10464
rect 15344 10424 15752 10452
rect 15344 10412 15350 10424
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 18049 10455 18107 10461
rect 18049 10452 18061 10455
rect 17920 10424 18061 10452
rect 17920 10412 17926 10424
rect 18049 10421 18061 10424
rect 18095 10421 18107 10455
rect 18049 10415 18107 10421
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 2038 10248 2044 10260
rect 1999 10220 2044 10248
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 2924 10220 4169 10248
rect 2924 10208 2930 10220
rect 4157 10217 4169 10220
rect 4203 10217 4215 10251
rect 4157 10211 4215 10217
rect 5537 10251 5595 10257
rect 5537 10217 5549 10251
rect 5583 10248 5595 10251
rect 5626 10248 5632 10260
rect 5583 10220 5632 10248
rect 5583 10217 5595 10220
rect 5537 10211 5595 10217
rect 5626 10208 5632 10220
rect 5684 10208 5690 10260
rect 6822 10248 6828 10260
rect 6783 10220 6828 10248
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7466 10208 7472 10260
rect 7524 10248 7530 10260
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 7524 10220 7849 10248
rect 7524 10208 7530 10220
rect 7837 10217 7849 10220
rect 7883 10217 7895 10251
rect 7837 10211 7895 10217
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 9490 10248 9496 10260
rect 8260 10220 9496 10248
rect 8260 10208 8266 10220
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 9674 10248 9680 10260
rect 9635 10220 9680 10248
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 12345 10251 12403 10257
rect 12345 10217 12357 10251
rect 12391 10248 12403 10251
rect 14366 10248 14372 10260
rect 12391 10220 14372 10248
rect 12391 10217 12403 10220
rect 12345 10211 12403 10217
rect 3418 10140 3424 10192
rect 3476 10180 3482 10192
rect 5718 10180 5724 10192
rect 3476 10152 5724 10180
rect 3476 10140 3482 10152
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 6546 10140 6552 10192
rect 6604 10180 6610 10192
rect 7190 10180 7196 10192
rect 6604 10152 7196 10180
rect 6604 10140 6610 10152
rect 7190 10140 7196 10152
rect 7248 10140 7254 10192
rect 9950 10180 9956 10192
rect 7484 10152 9956 10180
rect 3881 10115 3939 10121
rect 3881 10081 3893 10115
rect 3927 10112 3939 10115
rect 4801 10115 4859 10121
rect 4801 10112 4813 10115
rect 3927 10084 4813 10112
rect 3927 10081 3939 10084
rect 3881 10075 3939 10081
rect 4801 10081 4813 10084
rect 4847 10112 4859 10115
rect 5534 10112 5540 10124
rect 4847 10084 5540 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 7484 10121 7512 10152
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 7469 10115 7527 10121
rect 7469 10081 7481 10115
rect 7515 10081 7527 10115
rect 8478 10112 8484 10124
rect 8439 10084 8484 10112
rect 7469 10075 7527 10081
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 9125 10115 9183 10121
rect 9125 10081 9137 10115
rect 9171 10112 9183 10115
rect 9398 10112 9404 10124
rect 9171 10084 9404 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 12360 10112 12388 10211
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 15746 10248 15752 10260
rect 15707 10220 15752 10248
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 18785 10251 18843 10257
rect 18785 10248 18797 10251
rect 18656 10220 18797 10248
rect 18656 10208 18662 10220
rect 18785 10217 18797 10220
rect 18831 10217 18843 10251
rect 18785 10211 18843 10217
rect 19429 10251 19487 10257
rect 19429 10217 19441 10251
rect 19475 10248 19487 10251
rect 19610 10248 19616 10260
rect 19475 10220 19616 10248
rect 19475 10217 19487 10220
rect 19429 10211 19487 10217
rect 13814 10140 13820 10192
rect 13872 10180 13878 10192
rect 14093 10183 14151 10189
rect 14093 10180 14105 10183
rect 13872 10152 14105 10180
rect 13872 10140 13878 10152
rect 14093 10149 14105 10152
rect 14139 10149 14151 10183
rect 14093 10143 14151 10149
rect 9640 10084 12388 10112
rect 9640 10072 9646 10084
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 4982 10044 4988 10056
rect 2271 10016 4988 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 9306 10044 9312 10056
rect 9267 10016 9312 10044
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 12342 10004 12348 10056
rect 12400 10044 12406 10056
rect 13458 10047 13516 10053
rect 13458 10044 13470 10047
rect 12400 10016 13470 10044
rect 12400 10004 12406 10016
rect 13458 10013 13470 10016
rect 13504 10013 13516 10047
rect 13458 10007 13516 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 13906 10044 13912 10056
rect 13771 10016 13912 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 13906 10004 13912 10016
rect 13964 10044 13970 10056
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 13964 10016 15485 10044
rect 13964 10004 13970 10016
rect 15473 10013 15485 10016
rect 15519 10044 15531 10047
rect 16114 10044 16120 10056
rect 15519 10016 16120 10044
rect 15519 10013 15531 10016
rect 15473 10007 15531 10013
rect 16114 10004 16120 10016
rect 16172 10044 16178 10056
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16172 10016 17141 10044
rect 16172 10004 16178 10016
rect 17129 10013 17141 10016
rect 17175 10044 17187 10047
rect 17402 10044 17408 10056
rect 17175 10016 17408 10044
rect 17175 10013 17187 10016
rect 17129 10007 17187 10013
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 18800 10044 18828 10211
rect 19610 10208 19616 10220
rect 19668 10208 19674 10260
rect 19058 10044 19064 10056
rect 18800 10016 19064 10044
rect 19058 10004 19064 10016
rect 19116 10044 19122 10056
rect 19981 10047 20039 10053
rect 19116 10016 19932 10044
rect 19116 10004 19122 10016
rect 4525 9979 4583 9985
rect 4525 9945 4537 9979
rect 4571 9976 4583 9979
rect 5994 9976 6000 9988
rect 4571 9948 6000 9976
rect 4571 9945 4583 9948
rect 4525 9939 4583 9945
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 6549 9979 6607 9985
rect 6549 9945 6561 9979
rect 6595 9976 6607 9979
rect 7098 9976 7104 9988
rect 6595 9948 7104 9976
rect 6595 9945 6607 9948
rect 6549 9939 6607 9945
rect 7098 9936 7104 9948
rect 7156 9936 7162 9988
rect 8205 9979 8263 9985
rect 8205 9945 8217 9979
rect 8251 9976 8263 9979
rect 9214 9976 9220 9988
rect 8251 9948 8616 9976
rect 9175 9948 9220 9976
rect 8251 9945 8263 9948
rect 8205 9939 8263 9945
rect 8588 9920 8616 9948
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 10042 9936 10048 9988
rect 10100 9976 10106 9988
rect 10689 9979 10747 9985
rect 10689 9976 10701 9979
rect 10100 9948 10701 9976
rect 10100 9936 10106 9948
rect 10689 9945 10701 9948
rect 10735 9976 10747 9979
rect 15194 9976 15200 9988
rect 15252 9985 15258 9988
rect 10735 9948 14228 9976
rect 15164 9948 15200 9976
rect 10735 9945 10747 9948
rect 10689 9939 10747 9945
rect 4614 9908 4620 9920
rect 4575 9880 4620 9908
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 5810 9908 5816 9920
rect 5771 9880 5816 9908
rect 5810 9868 5816 9880
rect 5868 9868 5874 9920
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7193 9911 7251 9917
rect 7193 9908 7205 9911
rect 6972 9880 7205 9908
rect 6972 9868 6978 9880
rect 7193 9877 7205 9880
rect 7239 9877 7251 9911
rect 7193 9871 7251 9877
rect 7285 9911 7343 9917
rect 7285 9877 7297 9911
rect 7331 9908 7343 9911
rect 7834 9908 7840 9920
rect 7331 9880 7840 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 8352 9880 8397 9908
rect 8352 9868 8358 9880
rect 8570 9868 8576 9920
rect 8628 9868 8634 9920
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 10229 9911 10287 9917
rect 10229 9908 10241 9911
rect 9548 9880 10241 9908
rect 9548 9868 9554 9880
rect 10229 9877 10241 9880
rect 10275 9908 10287 9911
rect 10778 9908 10784 9920
rect 10275 9880 10784 9908
rect 10275 9877 10287 9880
rect 10229 9871 10287 9877
rect 10778 9868 10784 9880
rect 10836 9868 10842 9920
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 14090 9908 14096 9920
rect 10928 9880 14096 9908
rect 10928 9868 10934 9880
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 14200 9908 14228 9948
rect 15194 9936 15200 9948
rect 15252 9939 15264 9985
rect 16862 9979 16920 9985
rect 15304 9948 16574 9976
rect 15252 9936 15258 9939
rect 15304 9908 15332 9948
rect 14200 9880 15332 9908
rect 16546 9908 16574 9948
rect 16862 9945 16874 9979
rect 16908 9945 16920 9979
rect 16862 9939 16920 9945
rect 17672 9979 17730 9985
rect 17672 9945 17684 9979
rect 17718 9976 17730 9979
rect 17862 9976 17868 9988
rect 17718 9948 17868 9976
rect 17718 9945 17730 9948
rect 17672 9939 17730 9945
rect 16758 9908 16764 9920
rect 16546 9880 16764 9908
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 16868 9908 16896 9939
rect 17862 9936 17868 9948
rect 17920 9976 17926 9988
rect 19794 9976 19800 9988
rect 17920 9948 19800 9976
rect 17920 9936 17926 9948
rect 19794 9936 19800 9948
rect 19852 9936 19858 9988
rect 19904 9976 19932 10016
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 20714 10044 20720 10056
rect 20027 10016 20720 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 20714 10004 20720 10016
rect 20772 10044 20778 10056
rect 21266 10044 21272 10056
rect 20772 10016 21272 10044
rect 20772 10004 20778 10016
rect 21266 10004 21272 10016
rect 21324 10004 21330 10056
rect 20226 9979 20284 9985
rect 20226 9976 20238 9979
rect 19904 9948 20238 9976
rect 20226 9945 20238 9948
rect 20272 9945 20284 9979
rect 20226 9939 20284 9945
rect 16942 9908 16948 9920
rect 16868 9880 16948 9908
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 21358 9908 21364 9920
rect 21319 9880 21364 9908
rect 21358 9868 21364 9880
rect 21416 9868 21422 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 6052 9676 6745 9704
rect 6052 9664 6058 9676
rect 6733 9673 6745 9676
rect 6779 9673 6791 9707
rect 7834 9704 7840 9716
rect 7795 9676 7840 9704
rect 6733 9667 6791 9673
rect 7834 9664 7840 9676
rect 7892 9664 7898 9716
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 9401 9707 9459 9713
rect 9401 9704 9413 9707
rect 8352 9676 9413 9704
rect 8352 9664 8358 9676
rect 9401 9673 9413 9676
rect 9447 9673 9459 9707
rect 9401 9667 9459 9673
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 10413 9707 10471 9713
rect 10413 9704 10425 9707
rect 9815 9676 10425 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 10413 9673 10425 9676
rect 10459 9673 10471 9707
rect 10778 9704 10784 9716
rect 10739 9676 10784 9704
rect 10413 9667 10471 9673
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 13906 9704 13912 9716
rect 13867 9676 13912 9704
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 16114 9664 16120 9716
rect 16172 9704 16178 9716
rect 16669 9707 16727 9713
rect 16669 9704 16681 9707
rect 16172 9676 16681 9704
rect 16172 9664 16178 9676
rect 16669 9673 16681 9676
rect 16715 9673 16727 9707
rect 16669 9667 16727 9673
rect 17129 9707 17187 9713
rect 17129 9673 17141 9707
rect 17175 9704 17187 9707
rect 17218 9704 17224 9716
rect 17175 9676 17224 9704
rect 17175 9673 17187 9676
rect 17129 9667 17187 9673
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 17402 9664 17408 9716
rect 17460 9704 17466 9716
rect 17497 9707 17555 9713
rect 17497 9704 17509 9707
rect 17460 9676 17509 9704
rect 17460 9664 17466 9676
rect 17497 9673 17509 9676
rect 17543 9704 17555 9707
rect 18233 9707 18291 9713
rect 18233 9704 18245 9707
rect 17543 9676 18245 9704
rect 17543 9673 17555 9676
rect 17497 9667 17555 9673
rect 18233 9673 18245 9676
rect 18279 9704 18291 9707
rect 18877 9707 18935 9713
rect 18877 9704 18889 9707
rect 18279 9676 18889 9704
rect 18279 9673 18291 9676
rect 18233 9667 18291 9673
rect 18877 9673 18889 9676
rect 18923 9673 18935 9707
rect 19794 9704 19800 9716
rect 19755 9676 19800 9704
rect 18877 9667 18935 9673
rect 19794 9664 19800 9676
rect 19852 9664 19858 9716
rect 20257 9707 20315 9713
rect 20257 9673 20269 9707
rect 20303 9704 20315 9707
rect 20714 9704 20720 9716
rect 20303 9676 20720 9704
rect 20303 9673 20315 9676
rect 20257 9667 20315 9673
rect 20714 9664 20720 9676
rect 20772 9704 20778 9716
rect 20901 9707 20959 9713
rect 20901 9704 20913 9707
rect 20772 9676 20913 9704
rect 20772 9664 20778 9676
rect 20901 9673 20913 9676
rect 20947 9704 20959 9707
rect 21269 9707 21327 9713
rect 21269 9704 21281 9707
rect 20947 9676 21281 9704
rect 20947 9673 20959 9676
rect 20901 9667 20959 9673
rect 21269 9673 21281 9676
rect 21315 9673 21327 9707
rect 21269 9667 21327 9673
rect 5721 9639 5779 9645
rect 5721 9636 5733 9639
rect 2240 9608 5733 9636
rect 2240 9577 2268 9608
rect 5721 9605 5733 9608
rect 5767 9605 5779 9639
rect 7098 9636 7104 9648
rect 7059 9608 7104 9636
rect 5721 9599 5779 9605
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 8018 9596 8024 9648
rect 8076 9636 8082 9648
rect 9861 9639 9919 9645
rect 8076 9608 9720 9636
rect 8076 9596 8082 9608
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2774 9568 2780 9580
rect 2547 9540 2780 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2774 9528 2780 9540
rect 2832 9568 2838 9580
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 2832 9540 3065 9568
rect 2832 9528 2838 9540
rect 3053 9537 3065 9540
rect 3099 9537 3111 9571
rect 4522 9568 4528 9580
rect 4483 9540 4528 9568
rect 3053 9531 3111 9537
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9568 6055 9571
rect 7374 9568 7380 9580
rect 6043 9540 7380 9568
rect 6043 9537 6055 9540
rect 5997 9531 6055 9537
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9568 8815 9571
rect 9582 9568 9588 9580
rect 8803 9540 9588 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 2314 9460 2320 9512
rect 2372 9500 2378 9512
rect 4709 9503 4767 9509
rect 4709 9500 4721 9503
rect 2372 9472 4721 9500
rect 2372 9460 2378 9472
rect 4709 9469 4721 9472
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 5166 9460 5172 9512
rect 5224 9500 5230 9512
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 5224 9472 6377 9500
rect 5224 9460 5230 9472
rect 6365 9469 6377 9472
rect 6411 9500 6423 9503
rect 6914 9500 6920 9512
rect 6411 9472 6920 9500
rect 6411 9469 6423 9472
rect 6365 9463 6423 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7098 9460 7104 9512
rect 7156 9500 7162 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 7156 9472 7205 9500
rect 7156 9460 7162 9472
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 7282 9460 7288 9512
rect 7340 9500 7346 9512
rect 8849 9503 8907 9509
rect 7340 9472 7385 9500
rect 7340 9460 7346 9472
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 8849 9463 8907 9469
rect 2041 9435 2099 9441
rect 2041 9401 2053 9435
rect 2087 9432 2099 9435
rect 2958 9432 2964 9444
rect 2087 9404 2964 9432
rect 2087 9401 2099 9404
rect 2041 9395 2099 9401
rect 2958 9392 2964 9404
rect 3016 9392 3022 9444
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 5810 9432 5816 9444
rect 4120 9404 5816 9432
rect 4120 9392 4126 9404
rect 5810 9392 5816 9404
rect 5868 9392 5874 9444
rect 8386 9432 8392 9444
rect 8347 9404 8392 9432
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 8864 9432 8892 9463
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9692 9500 9720 9608
rect 9861 9605 9873 9639
rect 9907 9636 9919 9639
rect 12434 9636 12440 9648
rect 9907 9608 12440 9636
rect 9907 9605 9919 9608
rect 9861 9599 9919 9605
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 12986 9596 12992 9648
rect 13044 9636 13050 9648
rect 13274 9639 13332 9645
rect 13274 9636 13286 9639
rect 13044 9608 13286 9636
rect 13044 9596 13050 9608
rect 13274 9605 13286 9608
rect 13320 9605 13332 9639
rect 13274 9599 13332 9605
rect 10778 9528 10784 9580
rect 10836 9568 10842 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 10836 9540 11529 9568
rect 10836 9528 10842 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13924 9568 13952 9664
rect 18414 9596 18420 9648
rect 18472 9636 18478 9648
rect 18509 9639 18567 9645
rect 18509 9636 18521 9639
rect 18472 9608 18521 9636
rect 18472 9596 18478 9608
rect 18509 9605 18521 9608
rect 18555 9605 18567 9639
rect 19518 9636 19524 9648
rect 19479 9608 19524 9636
rect 18509 9599 18567 9605
rect 19518 9596 19524 9608
rect 19576 9596 19582 9648
rect 20530 9636 20536 9648
rect 20491 9608 20536 9636
rect 20530 9596 20536 9608
rect 20588 9596 20594 9648
rect 14461 9571 14519 9577
rect 14461 9568 14473 9571
rect 13587 9540 14473 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 14461 9537 14473 9540
rect 14507 9537 14519 9571
rect 14717 9571 14775 9577
rect 14717 9568 14729 9571
rect 14461 9531 14519 9537
rect 14568 9540 14729 9568
rect 10042 9500 10048 9512
rect 9692 9472 9904 9500
rect 10003 9472 10048 9500
rect 9674 9432 9680 9444
rect 8864 9404 9680 9432
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 9876 9432 9904 9472
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 10744 9472 10885 9500
rect 10744 9460 10750 9472
rect 10873 9469 10885 9472
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 14568 9500 14596 9540
rect 14717 9537 14729 9540
rect 14763 9537 14775 9571
rect 14717 9531 14775 9537
rect 11020 9472 11065 9500
rect 14476 9472 14596 9500
rect 11020 9460 11026 9472
rect 12161 9435 12219 9441
rect 12161 9432 12173 9435
rect 9876 9404 12173 9432
rect 12161 9401 12173 9404
rect 12207 9432 12219 9435
rect 12207 9404 12434 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 2685 9367 2743 9373
rect 2685 9364 2697 9367
rect 1728 9336 2697 9364
rect 1728 9324 1734 9336
rect 2685 9333 2697 9336
rect 2731 9333 2743 9367
rect 2685 9327 2743 9333
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 5902 9364 5908 9376
rect 4028 9336 5908 9364
rect 4028 9324 4034 9336
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 10870 9364 10876 9376
rect 7248 9336 10876 9364
rect 7248 9324 7254 9336
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 12406 9364 12434 9404
rect 14476 9364 14504 9472
rect 15838 9432 15844 9444
rect 15799 9404 15844 9432
rect 15838 9392 15844 9404
rect 15896 9432 15902 9444
rect 16942 9432 16948 9444
rect 15896 9404 16948 9432
rect 15896 9392 15902 9404
rect 16942 9392 16948 9404
rect 17000 9392 17006 9444
rect 16114 9364 16120 9376
rect 12406 9336 14504 9364
rect 16075 9336 16120 9364
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 2130 9160 2136 9172
rect 2091 9132 2136 9160
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 4522 9160 4528 9172
rect 4483 9132 4528 9160
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 8018 9160 8024 9172
rect 6972 9132 8024 9160
rect 6972 9120 6978 9132
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 9582 9160 9588 9172
rect 9543 9132 9588 9160
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 9732 9132 10609 9160
rect 9732 9120 9738 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 13262 9160 13268 9172
rect 11020 9132 13268 9160
rect 11020 9120 11026 9132
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 19058 9120 19064 9172
rect 19116 9160 19122 9172
rect 19797 9163 19855 9169
rect 19797 9160 19809 9163
rect 19116 9132 19809 9160
rect 19116 9120 19122 9132
rect 19797 9129 19809 9132
rect 19843 9129 19855 9163
rect 19797 9123 19855 9129
rect 3970 9052 3976 9104
rect 4028 9092 4034 9104
rect 9122 9092 9128 9104
rect 4028 9064 9128 9092
rect 4028 9052 4034 9064
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 14918 9092 14924 9104
rect 11348 9064 14924 9092
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 5166 9024 5172 9036
rect 4295 8996 5172 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 6181 9027 6239 9033
rect 6181 9024 6193 9027
rect 5684 8996 6193 9024
rect 5684 8984 5690 8996
rect 6181 8993 6193 8996
rect 6227 9024 6239 9027
rect 6638 9024 6644 9036
rect 6227 8996 6644 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6638 8984 6644 8996
rect 6696 9024 6702 9036
rect 9858 9024 9864 9036
rect 6696 8996 9864 9024
rect 6696 8984 6702 8996
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 10229 9027 10287 9033
rect 10229 8993 10241 9027
rect 10275 9024 10287 9027
rect 11241 9027 11299 9033
rect 11241 9024 11253 9027
rect 10275 8996 11253 9024
rect 10275 8993 10287 8996
rect 10229 8987 10287 8993
rect 11241 8993 11253 8996
rect 11287 9024 11299 9027
rect 11348 9024 11376 9064
rect 14918 9052 14924 9064
rect 14976 9052 14982 9104
rect 11287 8996 11376 9024
rect 12253 9027 12311 9033
rect 11287 8993 11299 8996
rect 11241 8987 11299 8993
rect 12253 8993 12265 9027
rect 12299 9024 12311 9027
rect 12526 9024 12532 9036
rect 12299 8996 12532 9024
rect 12299 8993 12311 8996
rect 12253 8987 12311 8993
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 2314 8956 2320 8968
rect 2275 8928 2320 8956
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5994 8956 6000 8968
rect 5031 8928 6000 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 8076 8928 10057 8956
rect 8076 8916 8082 8928
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 10778 8916 10784 8968
rect 10836 8956 10842 8968
rect 11977 8959 12035 8965
rect 11977 8956 11989 8959
rect 10836 8928 11989 8956
rect 10836 8916 10842 8928
rect 11977 8925 11989 8928
rect 12023 8925 12035 8959
rect 12621 8959 12679 8965
rect 12621 8956 12633 8959
rect 11977 8919 12035 8925
rect 12406 8928 12633 8956
rect 4893 8891 4951 8897
rect 4893 8857 4905 8891
rect 4939 8888 4951 8891
rect 5905 8891 5963 8897
rect 4939 8860 5580 8888
rect 4939 8857 4951 8860
rect 4893 8851 4951 8857
rect 5552 8829 5580 8860
rect 5905 8857 5917 8891
rect 5951 8888 5963 8891
rect 6549 8891 6607 8897
rect 6549 8888 6561 8891
rect 5951 8860 6561 8888
rect 5951 8857 5963 8860
rect 5905 8851 5963 8857
rect 6549 8857 6561 8860
rect 6595 8857 6607 8891
rect 6549 8851 6607 8857
rect 7282 8848 7288 8900
rect 7340 8888 7346 8900
rect 7653 8891 7711 8897
rect 7653 8888 7665 8891
rect 7340 8860 7665 8888
rect 7340 8848 7346 8860
rect 7653 8857 7665 8860
rect 7699 8888 7711 8891
rect 8202 8888 8208 8900
rect 7699 8860 8208 8888
rect 7699 8857 7711 8860
rect 7653 8851 7711 8857
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 9309 8891 9367 8897
rect 9309 8857 9321 8891
rect 9355 8888 9367 8891
rect 9953 8891 10011 8897
rect 9953 8888 9965 8891
rect 9355 8860 9965 8888
rect 9355 8857 9367 8860
rect 9309 8851 9367 8857
rect 9953 8857 9965 8860
rect 9999 8857 10011 8891
rect 9953 8851 10011 8857
rect 10965 8891 11023 8897
rect 10965 8857 10977 8891
rect 11011 8888 11023 8891
rect 11011 8860 11652 8888
rect 11011 8857 11023 8860
rect 10965 8851 11023 8857
rect 5537 8823 5595 8829
rect 5537 8789 5549 8823
rect 5583 8789 5595 8823
rect 5537 8783 5595 8789
rect 5997 8823 6055 8829
rect 5997 8789 6009 8823
rect 6043 8820 6055 8823
rect 6914 8820 6920 8832
rect 6043 8792 6920 8820
rect 6043 8789 6055 8792
rect 5997 8783 6055 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 7101 8823 7159 8829
rect 7101 8789 7113 8823
rect 7147 8820 7159 8823
rect 7190 8820 7196 8832
rect 7147 8792 7196 8820
rect 7147 8789 7159 8792
rect 7101 8783 7159 8789
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 9398 8820 9404 8832
rect 8619 8792 9404 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 11054 8820 11060 8832
rect 11015 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11624 8829 11652 8860
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8789 11667 8823
rect 12066 8820 12072 8832
rect 12027 8792 12072 8820
rect 11609 8783 11667 8789
rect 12066 8780 12072 8792
rect 12124 8820 12130 8832
rect 12406 8820 12434 8928
rect 12621 8925 12633 8928
rect 12667 8925 12679 8959
rect 12621 8919 12679 8925
rect 20349 8891 20407 8897
rect 20349 8888 20361 8891
rect 19260 8860 20361 8888
rect 12124 8792 12434 8820
rect 13725 8823 13783 8829
rect 12124 8780 12130 8792
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 16025 8823 16083 8829
rect 16025 8820 16037 8823
rect 13771 8792 16037 8820
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 16025 8789 16037 8792
rect 16071 8820 16083 8823
rect 16114 8820 16120 8832
rect 16071 8792 16120 8820
rect 16071 8789 16083 8792
rect 16025 8783 16083 8789
rect 16114 8780 16120 8792
rect 16172 8820 16178 8832
rect 19260 8829 19288 8860
rect 20349 8857 20361 8860
rect 20395 8888 20407 8891
rect 20717 8891 20775 8897
rect 20717 8888 20729 8891
rect 20395 8860 20729 8888
rect 20395 8857 20407 8860
rect 20349 8851 20407 8857
rect 20717 8857 20729 8860
rect 20763 8888 20775 8891
rect 21085 8891 21143 8897
rect 21085 8888 21097 8891
rect 20763 8860 21097 8888
rect 20763 8857 20775 8860
rect 20717 8851 20775 8857
rect 21085 8857 21097 8860
rect 21131 8888 21143 8891
rect 21266 8888 21272 8900
rect 21131 8860 21272 8888
rect 21131 8857 21143 8860
rect 21085 8851 21143 8857
rect 21266 8848 21272 8860
rect 21324 8848 21330 8900
rect 19245 8823 19303 8829
rect 19245 8820 19257 8823
rect 16172 8792 19257 8820
rect 16172 8780 16178 8792
rect 19245 8789 19257 8792
rect 19291 8789 19303 8823
rect 19245 8783 19303 8789
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 4706 8576 4712 8628
rect 4764 8616 4770 8628
rect 5169 8619 5227 8625
rect 5169 8616 5181 8619
rect 4764 8588 5181 8616
rect 4764 8576 4770 8588
rect 5169 8585 5181 8588
rect 5215 8616 5227 8619
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 5215 8588 6837 8616
rect 5215 8585 5227 8588
rect 5169 8579 5227 8585
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 7374 8616 7380 8628
rect 7335 8588 7380 8616
rect 6825 8579 6883 8585
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 8570 8576 8576 8628
rect 8628 8616 8634 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8628 8588 9045 8616
rect 8628 8576 8634 8588
rect 9033 8585 9045 8588
rect 9079 8585 9091 8619
rect 9398 8616 9404 8628
rect 9359 8588 9404 8616
rect 9033 8579 9091 8585
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 9824 8588 10425 8616
rect 9824 8576 9830 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 10413 8579 10471 8585
rect 10873 8619 10931 8625
rect 10873 8585 10885 8619
rect 10919 8616 10931 8619
rect 10962 8616 10968 8628
rect 10919 8588 10968 8616
rect 10919 8585 10931 8588
rect 10873 8579 10931 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11698 8616 11704 8628
rect 11659 8588 11704 8616
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 12434 8616 12440 8628
rect 12395 8588 12440 8616
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 20993 8619 21051 8625
rect 20993 8585 21005 8619
rect 21039 8616 21051 8619
rect 21082 8616 21088 8628
rect 21039 8588 21088 8616
rect 21039 8585 21051 8588
rect 20993 8579 21051 8585
rect 21082 8576 21088 8588
rect 21140 8576 21146 8628
rect 21266 8616 21272 8628
rect 21227 8588 21272 8616
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 5626 8548 5632 8560
rect 5587 8520 5632 8548
rect 5626 8508 5632 8520
rect 5684 8508 5690 8560
rect 7745 8551 7803 8557
rect 7745 8517 7757 8551
rect 7791 8548 7803 8551
rect 8662 8548 8668 8560
rect 7791 8520 8668 8548
rect 7791 8517 7803 8520
rect 7745 8511 7803 8517
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 12161 8551 12219 8557
rect 8772 8520 11100 8548
rect 6730 8480 6736 8492
rect 5552 8452 6736 8480
rect 5552 8424 5580 8452
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8480 7895 8483
rect 8386 8480 8392 8492
rect 7883 8452 8392 8480
rect 7883 8449 7895 8452
rect 7837 8443 7895 8449
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 4893 8415 4951 8421
rect 4893 8381 4905 8415
rect 4939 8412 4951 8415
rect 5534 8412 5540 8424
rect 4939 8384 5540 8412
rect 4939 8381 4951 8384
rect 4893 8375 4951 8381
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 7098 8412 7104 8424
rect 7055 8384 7104 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 5997 8347 6055 8353
rect 5997 8313 6009 8347
rect 6043 8344 6055 8347
rect 7024 8344 7052 8375
rect 7098 8372 7104 8384
rect 7156 8412 7162 8424
rect 7926 8412 7932 8424
rect 7156 8384 7932 8412
rect 7156 8372 7162 8384
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8412 8079 8415
rect 8110 8412 8116 8424
rect 8067 8384 8116 8412
rect 8067 8381 8079 8384
rect 8021 8375 8079 8381
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 8772 8412 8800 8520
rect 10134 8440 10140 8492
rect 10192 8480 10198 8492
rect 10781 8483 10839 8489
rect 10781 8480 10793 8483
rect 10192 8452 10793 8480
rect 10192 8440 10198 8452
rect 10781 8449 10793 8452
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 8260 8384 8800 8412
rect 9493 8415 9551 8421
rect 8260 8372 8266 8384
rect 9493 8381 9505 8415
rect 9539 8381 9551 8415
rect 9493 8375 9551 8381
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 10042 8412 10048 8424
rect 9723 8384 10048 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 9508 8344 9536 8375
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 10870 8372 10876 8424
rect 10928 8412 10934 8424
rect 10965 8415 11023 8421
rect 10965 8412 10977 8415
rect 10928 8384 10977 8412
rect 10928 8372 10934 8384
rect 10965 8381 10977 8384
rect 11011 8381 11023 8415
rect 11072 8412 11100 8520
rect 12161 8517 12173 8551
rect 12207 8548 12219 8551
rect 12250 8548 12256 8560
rect 12207 8520 12256 8548
rect 12207 8517 12219 8520
rect 12161 8511 12219 8517
rect 12250 8508 12256 8520
rect 12308 8548 12314 8560
rect 12897 8551 12955 8557
rect 12897 8548 12909 8551
rect 12308 8520 12909 8548
rect 12308 8508 12314 8520
rect 12897 8517 12909 8520
rect 12943 8517 12955 8551
rect 18506 8548 18512 8560
rect 12897 8511 12955 8517
rect 16546 8520 18512 8548
rect 11698 8440 11704 8492
rect 11756 8480 11762 8492
rect 12805 8483 12863 8489
rect 12805 8480 12817 8483
rect 11756 8452 12817 8480
rect 11756 8440 11762 8452
rect 12805 8449 12817 8452
rect 12851 8449 12863 8483
rect 12805 8443 12863 8449
rect 13081 8415 13139 8421
rect 11072 8384 12434 8412
rect 10965 8375 11023 8381
rect 6043 8316 7052 8344
rect 8680 8316 9536 8344
rect 6043 8313 6055 8316
rect 5997 8307 6055 8313
rect 6362 8276 6368 8288
rect 6323 8248 6368 8276
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 8018 8236 8024 8288
rect 8076 8276 8082 8288
rect 8680 8285 8708 8316
rect 9950 8304 9956 8356
rect 10008 8344 10014 8356
rect 10686 8344 10692 8356
rect 10008 8316 10692 8344
rect 10008 8304 10014 8316
rect 10060 8285 10088 8316
rect 10686 8304 10692 8316
rect 10744 8344 10750 8356
rect 12066 8344 12072 8356
rect 10744 8316 12072 8344
rect 10744 8304 10750 8316
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 12406 8344 12434 8384
rect 13081 8381 13093 8415
rect 13127 8412 13139 8415
rect 13262 8412 13268 8424
rect 13127 8384 13268 8412
rect 13127 8381 13139 8384
rect 13081 8375 13139 8381
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 16546 8344 16574 8520
rect 18506 8508 18512 8520
rect 18564 8508 18570 8560
rect 12406 8316 16574 8344
rect 8665 8279 8723 8285
rect 8665 8276 8677 8279
rect 8076 8248 8677 8276
rect 8076 8236 8082 8248
rect 8665 8245 8677 8248
rect 8711 8245 8723 8279
rect 8665 8239 8723 8245
rect 10045 8279 10103 8285
rect 10045 8245 10057 8279
rect 10091 8245 10103 8279
rect 10045 8239 10103 8245
rect 10318 8236 10324 8288
rect 10376 8276 10382 8288
rect 15010 8276 15016 8288
rect 10376 8248 15016 8276
rect 10376 8236 10382 8248
rect 15010 8236 15016 8248
rect 15068 8236 15074 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 5994 8072 6000 8084
rect 5955 8044 6000 8072
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8720 8044 8953 8072
rect 8720 8032 8726 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10597 8075 10655 8081
rect 10597 8072 10609 8075
rect 10100 8044 10609 8072
rect 10100 8032 10106 8044
rect 10597 8041 10609 8044
rect 10643 8041 10655 8075
rect 10597 8035 10655 8041
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 11112 8044 12265 8072
rect 11112 8032 11118 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 13262 8072 13268 8084
rect 12253 8035 12311 8041
rect 12728 8044 13268 8072
rect 4614 7964 4620 8016
rect 4672 8004 4678 8016
rect 7285 8007 7343 8013
rect 7285 8004 7297 8007
rect 4672 7976 7297 8004
rect 4672 7964 4678 7976
rect 7285 7973 7297 7976
rect 7331 7973 7343 8007
rect 7285 7967 7343 7973
rect 8110 7964 8116 8016
rect 8168 8004 8174 8016
rect 10318 8004 10324 8016
rect 8168 7976 10324 8004
rect 8168 7964 8174 7976
rect 10318 7964 10324 7976
rect 10376 7964 10382 8016
rect 11146 7964 11152 8016
rect 11204 8004 11210 8016
rect 11241 8007 11299 8013
rect 11241 8004 11253 8007
rect 11204 7976 11253 8004
rect 11204 7964 11210 7976
rect 11241 7973 11253 7976
rect 11287 7973 11299 8007
rect 11241 7967 11299 7973
rect 11698 7964 11704 8016
rect 11756 8004 11762 8016
rect 11882 8004 11888 8016
rect 11756 7976 11888 8004
rect 11756 7964 11762 7976
rect 11882 7964 11888 7976
rect 11940 8004 11946 8016
rect 11940 7976 12434 8004
rect 11940 7964 11946 7976
rect 6362 7896 6368 7948
rect 6420 7936 6426 7948
rect 6457 7939 6515 7945
rect 6457 7936 6469 7939
rect 6420 7908 6469 7936
rect 6420 7896 6426 7908
rect 6457 7905 6469 7908
rect 6503 7905 6515 7939
rect 6638 7936 6644 7948
rect 6599 7908 6644 7936
rect 6457 7899 6515 7905
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 7742 7936 7748 7948
rect 7703 7908 7748 7936
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7936 7987 7939
rect 8202 7936 8208 7948
rect 7975 7908 8208 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 9582 7936 9588 7948
rect 9543 7908 9588 7936
rect 9582 7896 9588 7908
rect 9640 7896 9646 7948
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 6788 7840 7665 7868
rect 6788 7828 6794 7840
rect 7653 7837 7665 7840
rect 7699 7868 7711 7871
rect 10134 7868 10140 7880
rect 7699 7840 10140 7868
rect 7699 7837 7711 7840
rect 7653 7831 7711 7837
rect 10134 7828 10140 7840
rect 10192 7868 10198 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 10192 7840 10241 7868
rect 10192 7828 10198 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 8573 7803 8631 7809
rect 8573 7769 8585 7803
rect 8619 7800 8631 7803
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 8619 7772 9321 7800
rect 8619 7769 8631 7772
rect 8573 7763 8631 7769
rect 9309 7769 9321 7772
rect 9355 7769 9367 7803
rect 12406 7800 12434 7976
rect 12728 7945 12756 8044
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 12713 7939 12771 7945
rect 12713 7905 12725 7939
rect 12759 7905 12771 7939
rect 12713 7899 12771 7905
rect 12805 7939 12863 7945
rect 12805 7905 12817 7939
rect 12851 7905 12863 7939
rect 12805 7899 12863 7905
rect 12526 7828 12532 7880
rect 12584 7868 12590 7880
rect 12820 7868 12848 7899
rect 12584 7840 12848 7868
rect 12584 7828 12590 7840
rect 12621 7803 12679 7809
rect 12621 7800 12633 7803
rect 12406 7772 12633 7800
rect 9309 7763 9367 7769
rect 12621 7769 12633 7772
rect 12667 7769 12679 7803
rect 12621 7763 12679 7769
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 5629 7735 5687 7741
rect 5629 7732 5641 7735
rect 5592 7704 5641 7732
rect 5592 7692 5598 7704
rect 5629 7701 5641 7704
rect 5675 7701 5687 7735
rect 5629 7695 5687 7701
rect 6365 7735 6423 7741
rect 6365 7701 6377 7735
rect 6411 7732 6423 7735
rect 7006 7732 7012 7744
rect 6411 7704 7012 7732
rect 6411 7701 6423 7704
rect 6365 7695 6423 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 9398 7732 9404 7744
rect 9359 7704 9404 7732
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 6638 7528 6644 7540
rect 6043 7500 6644 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7006 7528 7012 7540
rect 6967 7500 7012 7528
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 8110 7528 8116 7540
rect 8071 7500 8116 7528
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8386 7528 8392 7540
rect 8347 7500 8392 7528
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 9493 7531 9551 7537
rect 9493 7497 9505 7531
rect 9539 7528 9551 7531
rect 9582 7528 9588 7540
rect 9539 7500 9588 7528
rect 9539 7497 9551 7500
rect 9493 7491 9551 7497
rect 9582 7488 9588 7500
rect 9640 7528 9646 7540
rect 9861 7531 9919 7537
rect 9861 7528 9873 7531
rect 9640 7500 9873 7528
rect 9640 7488 9646 7500
rect 9861 7497 9873 7500
rect 9907 7528 9919 7531
rect 18690 7528 18696 7540
rect 9907 7500 18696 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 6733 7463 6791 7469
rect 6733 7429 6745 7463
rect 6779 7460 6791 7463
rect 7098 7460 7104 7472
rect 6779 7432 7104 7460
rect 6779 7429 6791 7432
rect 6733 7423 6791 7429
rect 7098 7420 7104 7432
rect 7156 7460 7162 7472
rect 8849 7463 8907 7469
rect 7156 7432 7512 7460
rect 7156 7420 7162 7432
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 5776 7364 7389 7392
rect 5776 7352 5782 7364
rect 6748 7256 6776 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7484 7392 7512 7432
rect 8849 7429 8861 7463
rect 8895 7460 8907 7463
rect 10318 7460 10324 7472
rect 8895 7432 10324 7460
rect 8895 7429 8907 7432
rect 8849 7423 8907 7429
rect 10318 7420 10324 7432
rect 10376 7420 10382 7472
rect 8757 7395 8815 7401
rect 7484 7364 7604 7392
rect 7377 7355 7435 7361
rect 7576 7336 7604 7364
rect 8757 7361 8769 7395
rect 8803 7392 8815 7395
rect 9122 7392 9128 7404
rect 8803 7364 9128 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 7469 7327 7527 7333
rect 7469 7324 7481 7327
rect 6880 7296 7481 7324
rect 6880 7284 6886 7296
rect 7469 7293 7481 7296
rect 7515 7293 7527 7327
rect 7469 7287 7527 7293
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 9033 7327 9091 7333
rect 7616 7296 7709 7324
rect 7616 7284 7622 7296
rect 9033 7293 9045 7327
rect 9079 7324 9091 7327
rect 9582 7324 9588 7336
rect 9079 7296 9588 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9582 7284 9588 7296
rect 9640 7284 9646 7336
rect 8478 7256 8484 7268
rect 6748 7228 8484 7256
rect 8478 7216 8484 7228
rect 8536 7216 8542 7268
rect 5629 7191 5687 7197
rect 5629 7157 5641 7191
rect 5675 7188 5687 7191
rect 5718 7188 5724 7200
rect 5675 7160 5724 7188
rect 5675 7157 5687 7160
rect 5629 7151 5687 7157
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 10229 7191 10287 7197
rect 10229 7157 10241 7191
rect 10275 7188 10287 7191
rect 10962 7188 10968 7200
rect 10275 7160 10968 7188
rect 10275 7157 10287 7160
rect 10229 7151 10287 7157
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 3418 6944 3424 6996
rect 3476 6984 3482 6996
rect 4709 6987 4767 6993
rect 4709 6984 4721 6987
rect 3476 6956 4721 6984
rect 3476 6944 3482 6956
rect 4709 6953 4721 6956
rect 4755 6953 4767 6987
rect 4709 6947 4767 6953
rect 9033 6987 9091 6993
rect 9033 6953 9045 6987
rect 9079 6984 9091 6987
rect 9398 6984 9404 6996
rect 9079 6956 9404 6984
rect 9079 6953 9091 6956
rect 9033 6947 9091 6953
rect 4724 6780 4752 6947
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 10318 6984 10324 6996
rect 10279 6956 10324 6984
rect 10318 6944 10324 6956
rect 10376 6944 10382 6996
rect 5261 6919 5319 6925
rect 5261 6885 5273 6919
rect 5307 6885 5319 6919
rect 5261 6879 5319 6885
rect 5276 6848 5304 6879
rect 10870 6876 10876 6928
rect 10928 6916 10934 6928
rect 10928 6888 11100 6916
rect 10928 6876 10934 6888
rect 5276 6820 7512 6848
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4724 6752 5089 6780
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5626 6780 5632 6792
rect 5587 6752 5632 6780
rect 5077 6743 5135 6749
rect 5626 6740 5632 6752
rect 5684 6740 5690 6792
rect 5902 6740 5908 6792
rect 5960 6780 5966 6792
rect 6181 6783 6239 6789
rect 6181 6780 6193 6783
rect 5960 6752 6193 6780
rect 5960 6740 5966 6752
rect 6181 6749 6193 6752
rect 6227 6749 6239 6783
rect 7484 6780 7512 6820
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 7616 6820 7661 6848
rect 7616 6808 7622 6820
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 8297 6851 8355 6857
rect 8297 6848 8309 6851
rect 8260 6820 8309 6848
rect 8260 6808 8266 6820
rect 8297 6817 8309 6820
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 9766 6848 9772 6860
rect 9723 6820 9772 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 9766 6808 9772 6820
rect 9824 6848 9830 6860
rect 10962 6848 10968 6860
rect 9824 6820 10968 6848
rect 9824 6808 9830 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11072 6848 11100 6888
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 11072 6820 11805 6848
rect 11793 6817 11805 6820
rect 11839 6848 11851 6851
rect 11974 6848 11980 6860
rect 11839 6820 11980 6848
rect 11839 6817 11851 6820
rect 11793 6811 11851 6817
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 19886 6780 19892 6792
rect 7484 6752 19892 6780
rect 6181 6743 6239 6749
rect 19886 6740 19892 6752
rect 19944 6740 19950 6792
rect 21542 6712 21548 6724
rect 5828 6684 21548 6712
rect 5828 6653 5856 6684
rect 21542 6672 21548 6684
rect 21600 6672 21606 6724
rect 5813 6647 5871 6653
rect 5813 6613 5825 6647
rect 5859 6613 5871 6647
rect 5813 6607 5871 6613
rect 6365 6647 6423 6653
rect 6365 6613 6377 6647
rect 6411 6644 6423 6647
rect 6914 6644 6920 6656
rect 6411 6616 6920 6644
rect 6411 6613 6423 6616
rect 6365 6607 6423 6613
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 7374 6644 7380 6656
rect 7064 6616 7109 6644
rect 7335 6616 7380 6644
rect 7064 6604 7070 6616
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 7524 6616 7569 6644
rect 7524 6604 7530 6616
rect 8202 6604 8208 6656
rect 8260 6644 8266 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 8260 6616 9413 6644
rect 8260 6604 8266 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9401 6607 9459 6613
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 9548 6616 9593 6644
rect 9548 6604 9554 6616
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 10192 6616 10701 6644
rect 10192 6604 10198 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10689 6607 10747 6613
rect 10781 6647 10839 6653
rect 10781 6613 10793 6647
rect 10827 6644 10839 6647
rect 10870 6644 10876 6656
rect 10827 6616 10876 6644
rect 10827 6613 10839 6616
rect 10781 6607 10839 6613
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 11020 6616 11437 6644
rect 11020 6604 11026 6616
rect 11425 6613 11437 6616
rect 11471 6644 11483 6647
rect 18966 6644 18972 6656
rect 11471 6616 18972 6644
rect 11471 6613 11483 6616
rect 11425 6607 11483 6613
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 5537 6443 5595 6449
rect 5537 6440 5549 6443
rect 4120 6412 5549 6440
rect 4120 6400 4126 6412
rect 5537 6409 5549 6412
rect 5583 6440 5595 6443
rect 5626 6440 5632 6452
rect 5583 6412 5632 6440
rect 5583 6409 5595 6412
rect 5537 6403 5595 6409
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 7800 6412 8125 6440
rect 7800 6400 7806 6412
rect 8113 6409 8125 6412
rect 8159 6409 8171 6443
rect 9122 6440 9128 6452
rect 9083 6412 9128 6440
rect 8113 6403 8171 6409
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 10134 6440 10140 6452
rect 10095 6412 10140 6440
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 10962 6440 10968 6452
rect 10643 6412 10968 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 21450 6440 21456 6452
rect 16546 6412 21456 6440
rect 6914 6332 6920 6384
rect 6972 6372 6978 6384
rect 16546 6372 16574 6412
rect 21450 6400 21456 6412
rect 21508 6400 21514 6452
rect 6972 6344 16574 6372
rect 6972 6332 6978 6344
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 7616 6276 7757 6304
rect 7616 6264 7622 6276
rect 7745 6273 7757 6276
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 8536 6276 9505 6304
rect 8536 6264 8542 6276
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 4062 6196 4068 6248
rect 4120 6236 4126 6248
rect 5902 6236 5908 6248
rect 4120 6208 5908 6236
rect 4120 6196 4126 6208
rect 5902 6196 5908 6208
rect 5960 6196 5966 6248
rect 6822 6236 6828 6248
rect 6380 6208 6828 6236
rect 5626 6128 5632 6180
rect 5684 6168 5690 6180
rect 6380 6168 6408 6208
rect 6822 6196 6828 6208
rect 6880 6236 6886 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6880 6208 6929 6236
rect 6880 6196 6886 6208
rect 6917 6205 6929 6208
rect 6963 6236 6975 6239
rect 9306 6236 9312 6248
rect 6963 6208 9312 6236
rect 6963 6205 6975 6208
rect 6917 6199 6975 6205
rect 9306 6196 9312 6208
rect 9364 6236 9370 6248
rect 9585 6239 9643 6245
rect 9585 6236 9597 6239
rect 9364 6208 9597 6236
rect 9364 6196 9370 6208
rect 9585 6205 9597 6208
rect 9631 6205 9643 6239
rect 9766 6236 9772 6248
rect 9727 6208 9772 6236
rect 9585 6199 9643 6205
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 7374 6168 7380 6180
rect 5684 6140 6408 6168
rect 6472 6140 7380 6168
rect 5684 6128 5690 6140
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 6472 6109 6500 6140
rect 7374 6128 7380 6140
rect 7432 6128 7438 6180
rect 6457 6103 6515 6109
rect 6457 6100 6469 6103
rect 4212 6072 6469 6100
rect 4212 6060 4218 6072
rect 6457 6069 6469 6072
rect 6503 6069 6515 6103
rect 7190 6100 7196 6112
rect 7151 6072 7196 6100
rect 6457 6063 6515 6069
rect 7190 6060 7196 6072
rect 7248 6100 7254 6112
rect 7466 6100 7472 6112
rect 7248 6072 7472 6100
rect 7248 6060 7254 6072
rect 7466 6060 7472 6072
rect 7524 6100 7530 6112
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 7524 6072 8769 6100
rect 7524 6060 7530 6072
rect 8757 6069 8769 6072
rect 8803 6100 8815 6103
rect 9490 6100 9496 6112
rect 8803 6072 9496 6100
rect 8803 6069 8815 6072
rect 8757 6063 8815 6069
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 8202 5896 8208 5908
rect 7432 5868 8208 5896
rect 7432 5856 7438 5868
rect 8202 5856 8208 5868
rect 8260 5896 8266 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8260 5868 8953 5896
rect 8260 5856 8266 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 9306 5896 9312 5908
rect 9267 5868 9312 5896
rect 8941 5859 8999 5865
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 8478 5828 8484 5840
rect 8439 5800 8484 5828
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 10870 5624 10876 5636
rect 4120 5596 10876 5624
rect 4120 5584 4126 5596
rect 10870 5584 10876 5596
rect 10928 5584 10934 5636
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 7650 5352 7656 5364
rect 4120 5324 7656 5352
rect 4120 5312 4126 5324
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 3970 5244 3976 5296
rect 4028 5284 4034 5296
rect 7190 5284 7196 5296
rect 4028 5256 7196 5284
rect 4028 5244 4034 5256
rect 7190 5244 7196 5256
rect 7248 5244 7254 5296
rect 10870 5216 10876 5228
rect 10831 5188 10876 5216
rect 10870 5176 10876 5188
rect 10928 5216 10934 5228
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 10928 5188 11529 5216
rect 10928 5176 10934 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 11057 5083 11115 5089
rect 11057 5049 11069 5083
rect 11103 5080 11115 5083
rect 21174 5080 21180 5092
rect 11103 5052 21180 5080
rect 11103 5049 11115 5052
rect 11057 5043 11115 5049
rect 21174 5040 21180 5052
rect 21232 5040 21238 5092
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 5718 4128 5724 4140
rect 4120 4100 5724 4128
rect 4120 4088 4126 4100
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 8294 4060 8300 4072
rect 3476 4032 8300 4060
rect 3476 4020 3482 4032
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 3970 3952 3976 4004
rect 4028 3992 4034 4004
rect 9950 3992 9956 4004
rect 4028 3964 9956 3992
rect 4028 3952 4034 3964
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 3510 2592 3516 2644
rect 3568 2632 3574 2644
rect 11882 2632 11888 2644
rect 3568 2604 11888 2632
rect 3568 2592 3574 2604
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 4062 2524 4068 2576
rect 4120 2564 4126 2576
rect 5626 2564 5632 2576
rect 4120 2536 5632 2564
rect 4120 2524 4126 2536
rect 5626 2524 5632 2536
rect 5684 2524 5690 2576
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 2866 1776 2872 1828
rect 2924 1816 2930 1828
rect 5534 1816 5540 1828
rect 2924 1788 5540 1816
rect 2924 1776 2930 1788
rect 5534 1776 5540 1788
rect 5592 1776 5598 1828
<< via1 >>
rect 21180 20748 21232 20800
rect 21824 20748 21876 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 5264 20544 5316 20596
rect 5356 20544 5408 20596
rect 12532 20544 12584 20596
rect 6000 20408 6052 20460
rect 13084 20476 13136 20528
rect 5540 20340 5592 20392
rect 5816 20272 5868 20324
rect 6184 20340 6236 20392
rect 7012 20408 7064 20460
rect 8300 20451 8352 20460
rect 8300 20417 8309 20451
rect 8309 20417 8343 20451
rect 8343 20417 8352 20451
rect 8300 20408 8352 20417
rect 9496 20451 9548 20460
rect 9496 20417 9505 20451
rect 9505 20417 9539 20451
rect 9539 20417 9548 20451
rect 9496 20408 9548 20417
rect 10140 20451 10192 20460
rect 10140 20417 10149 20451
rect 10149 20417 10183 20451
rect 10183 20417 10192 20451
rect 10140 20408 10192 20417
rect 22284 20408 22336 20460
rect 6736 20272 6788 20324
rect 10048 20340 10100 20392
rect 21364 20340 21416 20392
rect 5632 20247 5684 20256
rect 5632 20213 5641 20247
rect 5641 20213 5675 20247
rect 5675 20213 5684 20247
rect 5632 20204 5684 20213
rect 6828 20204 6880 20256
rect 7932 20247 7984 20256
rect 7932 20213 7941 20247
rect 7941 20213 7975 20247
rect 7975 20213 7984 20247
rect 7932 20204 7984 20213
rect 9312 20204 9364 20256
rect 14924 20272 14976 20324
rect 13544 20204 13596 20256
rect 19064 20204 19116 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 1492 20043 1544 20052
rect 1492 20009 1501 20043
rect 1501 20009 1535 20043
rect 1535 20009 1544 20043
rect 1492 20000 1544 20009
rect 2044 20043 2096 20052
rect 2044 20009 2053 20043
rect 2053 20009 2087 20043
rect 2087 20009 2096 20043
rect 2044 20000 2096 20009
rect 2780 20000 2832 20052
rect 5172 20000 5224 20052
rect 1400 19932 1452 19984
rect 2504 19932 2556 19984
rect 4160 19932 4212 19984
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 2504 19839 2556 19848
rect 2504 19805 2513 19839
rect 2513 19805 2547 19839
rect 2547 19805 2556 19839
rect 2504 19796 2556 19805
rect 5356 19796 5408 19848
rect 5816 19796 5868 19848
rect 18972 20000 19024 20052
rect 9404 19975 9456 19984
rect 9404 19941 9413 19975
rect 9413 19941 9447 19975
rect 9447 19941 9456 19975
rect 9404 19932 9456 19941
rect 9864 19932 9916 19984
rect 10416 19932 10468 19984
rect 15844 19932 15896 19984
rect 6736 19796 6788 19848
rect 9404 19796 9456 19848
rect 11980 19864 12032 19916
rect 12716 19864 12768 19916
rect 16304 19864 16356 19916
rect 9864 19839 9916 19848
rect 9864 19805 9873 19839
rect 9873 19805 9907 19839
rect 9907 19805 9916 19839
rect 9864 19796 9916 19805
rect 10692 19839 10744 19848
rect 10692 19805 10701 19839
rect 10701 19805 10735 19839
rect 10735 19805 10744 19839
rect 10692 19796 10744 19805
rect 11244 19839 11296 19848
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 12808 19796 12860 19848
rect 15292 19796 15344 19848
rect 18512 19796 18564 19848
rect 5264 19728 5316 19780
rect 6828 19728 6880 19780
rect 5448 19660 5500 19712
rect 6184 19660 6236 19712
rect 6552 19660 6604 19712
rect 7472 19660 7524 19712
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 15384 19728 15436 19780
rect 19064 19796 19116 19848
rect 21364 19839 21416 19848
rect 21364 19805 21373 19839
rect 21373 19805 21407 19839
rect 21407 19805 21416 19839
rect 21364 19796 21416 19805
rect 20168 19728 20220 19780
rect 20996 19728 21048 19780
rect 7564 19660 7616 19669
rect 13728 19660 13780 19712
rect 14648 19660 14700 19712
rect 18328 19660 18380 19712
rect 19432 19660 19484 19712
rect 20720 19660 20772 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 5172 19456 5224 19508
rect 6000 19499 6052 19508
rect 6000 19465 6009 19499
rect 6009 19465 6043 19499
rect 6043 19465 6052 19499
rect 6000 19456 6052 19465
rect 6552 19456 6604 19508
rect 7472 19499 7524 19508
rect 1584 19388 1636 19440
rect 1676 19388 1728 19440
rect 4528 19388 4580 19440
rect 3424 19320 3476 19372
rect 3884 19363 3936 19372
rect 3884 19329 3893 19363
rect 3893 19329 3927 19363
rect 3927 19329 3936 19363
rect 3884 19320 3936 19329
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 7472 19465 7481 19499
rect 7481 19465 7515 19499
rect 7515 19465 7524 19499
rect 7472 19456 7524 19465
rect 7564 19388 7616 19440
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 3056 19252 3108 19304
rect 7564 19252 7616 19304
rect 7932 19252 7984 19304
rect 9588 19363 9640 19372
rect 9588 19329 9597 19363
rect 9597 19329 9631 19363
rect 9631 19329 9640 19363
rect 9588 19320 9640 19329
rect 9956 19320 10008 19372
rect 13636 19456 13688 19508
rect 13728 19456 13780 19508
rect 12716 19320 12768 19372
rect 12992 19320 13044 19372
rect 10232 19252 10284 19304
rect 14280 19456 14332 19508
rect 17500 19456 17552 19508
rect 16764 19388 16816 19440
rect 15200 19363 15252 19372
rect 15200 19329 15218 19363
rect 15218 19329 15252 19363
rect 15200 19320 15252 19329
rect 16580 19320 16632 19372
rect 20812 19363 20864 19372
rect 20812 19329 20830 19363
rect 20830 19329 20864 19363
rect 20812 19320 20864 19329
rect 15752 19295 15804 19304
rect 15752 19261 15761 19295
rect 15761 19261 15795 19295
rect 15795 19261 15804 19295
rect 15752 19252 15804 19261
rect 18236 19252 18288 19304
rect 19892 19252 19944 19304
rect 21088 19295 21140 19304
rect 21088 19261 21097 19295
rect 21097 19261 21131 19295
rect 21131 19261 21140 19295
rect 21088 19252 21140 19261
rect 21364 19252 21416 19304
rect 1124 19116 1176 19168
rect 5632 19184 5684 19236
rect 3516 19116 3568 19168
rect 4252 19116 4304 19168
rect 4528 19159 4580 19168
rect 4528 19125 4537 19159
rect 4537 19125 4571 19159
rect 4571 19125 4580 19159
rect 4528 19116 4580 19125
rect 5264 19116 5316 19168
rect 7840 19159 7892 19168
rect 7840 19125 7849 19159
rect 7849 19125 7883 19159
rect 7883 19125 7892 19159
rect 7840 19116 7892 19125
rect 7932 19116 7984 19168
rect 12808 19116 12860 19168
rect 17960 19184 18012 19236
rect 19340 19184 19392 19236
rect 16948 19116 17000 19168
rect 18328 19159 18380 19168
rect 18328 19125 18337 19159
rect 18337 19125 18371 19159
rect 18371 19125 18380 19159
rect 18328 19116 18380 19125
rect 19616 19116 19668 19168
rect 19708 19159 19760 19168
rect 19708 19125 19717 19159
rect 19717 19125 19751 19159
rect 19751 19125 19760 19159
rect 19708 19116 19760 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 2136 18912 2188 18964
rect 4160 18912 4212 18964
rect 4988 18912 5040 18964
rect 5724 18912 5776 18964
rect 12440 18912 12492 18964
rect 12532 18912 12584 18964
rect 18604 18912 18656 18964
rect 18696 18912 18748 18964
rect 22744 18912 22796 18964
rect 2320 18887 2372 18896
rect 2320 18853 2329 18887
rect 2329 18853 2363 18887
rect 2363 18853 2372 18887
rect 2320 18844 2372 18853
rect 2964 18844 3016 18896
rect 4528 18844 4580 18896
rect 3148 18776 3200 18828
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 15568 18844 15620 18896
rect 16488 18844 16540 18896
rect 12532 18776 12584 18828
rect 204 18572 256 18624
rect 5540 18640 5592 18692
rect 5080 18615 5132 18624
rect 5080 18581 5089 18615
rect 5089 18581 5123 18615
rect 5123 18581 5132 18615
rect 5080 18572 5132 18581
rect 5724 18572 5776 18624
rect 6828 18640 6880 18692
rect 6276 18572 6328 18624
rect 7380 18615 7432 18624
rect 7380 18581 7389 18615
rect 7389 18581 7423 18615
rect 7423 18581 7432 18615
rect 7380 18572 7432 18581
rect 9772 18751 9824 18760
rect 8116 18640 8168 18692
rect 9772 18717 9781 18751
rect 9781 18717 9815 18751
rect 9815 18717 9824 18751
rect 9772 18708 9824 18717
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 10232 18708 10284 18760
rect 13728 18751 13780 18760
rect 9680 18640 9732 18692
rect 12532 18640 12584 18692
rect 13268 18640 13320 18692
rect 13452 18683 13504 18692
rect 13452 18649 13470 18683
rect 13470 18649 13504 18683
rect 13452 18640 13504 18649
rect 13728 18717 13737 18751
rect 13737 18717 13771 18751
rect 13771 18717 13780 18751
rect 13728 18708 13780 18717
rect 15752 18751 15804 18760
rect 14464 18640 14516 18692
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 18328 18708 18380 18760
rect 21088 18708 21140 18760
rect 15292 18640 15344 18692
rect 16120 18640 16172 18692
rect 8208 18615 8260 18624
rect 8208 18581 8217 18615
rect 8217 18581 8251 18615
rect 8251 18581 8260 18615
rect 8208 18572 8260 18581
rect 11796 18572 11848 18624
rect 12072 18572 12124 18624
rect 12716 18572 12768 18624
rect 14188 18572 14240 18624
rect 19340 18640 19392 18692
rect 18420 18615 18472 18624
rect 18420 18581 18429 18615
rect 18429 18581 18463 18615
rect 18463 18581 18472 18615
rect 19708 18640 19760 18692
rect 18420 18572 18472 18581
rect 20260 18572 20312 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 4160 18368 4212 18420
rect 5356 18368 5408 18420
rect 5908 18368 5960 18420
rect 6828 18368 6880 18420
rect 7840 18368 7892 18420
rect 8208 18368 8260 18420
rect 2504 18343 2556 18352
rect 2504 18309 2513 18343
rect 2513 18309 2547 18343
rect 2547 18309 2556 18343
rect 2504 18300 2556 18309
rect 3424 18300 3476 18352
rect 7380 18300 7432 18352
rect 10140 18300 10192 18352
rect 2780 18275 2832 18284
rect 2780 18241 2789 18275
rect 2789 18241 2823 18275
rect 2823 18241 2832 18275
rect 2780 18232 2832 18241
rect 5448 18232 5500 18284
rect 7656 18275 7708 18284
rect 7656 18241 7665 18275
rect 7665 18241 7699 18275
rect 7699 18241 7708 18275
rect 7656 18232 7708 18241
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 10784 18275 10836 18284
rect 10784 18241 10793 18275
rect 10793 18241 10827 18275
rect 10827 18241 10836 18275
rect 10784 18232 10836 18241
rect 4436 18164 4488 18216
rect 4712 18164 4764 18216
rect 3240 18139 3292 18148
rect 3240 18105 3249 18139
rect 3249 18105 3283 18139
rect 3283 18105 3292 18139
rect 3240 18096 3292 18105
rect 3424 18096 3476 18148
rect 4804 18096 4856 18148
rect 7840 18164 7892 18216
rect 12440 18368 12492 18420
rect 12532 18368 12584 18420
rect 15200 18368 15252 18420
rect 15384 18368 15436 18420
rect 20996 18368 21048 18420
rect 11796 18300 11848 18352
rect 12716 18300 12768 18352
rect 17684 18300 17736 18352
rect 13452 18232 13504 18284
rect 4896 18028 4948 18080
rect 5632 18071 5684 18080
rect 5632 18037 5641 18071
rect 5641 18037 5675 18071
rect 5675 18037 5684 18071
rect 5632 18028 5684 18037
rect 6092 18028 6144 18080
rect 6920 18071 6972 18080
rect 6920 18037 6929 18071
rect 6929 18037 6963 18071
rect 6963 18037 6972 18071
rect 6920 18028 6972 18037
rect 8576 18096 8628 18148
rect 8668 18028 8720 18080
rect 10508 18028 10560 18080
rect 10876 18028 10928 18080
rect 11796 18028 11848 18080
rect 15476 18275 15528 18284
rect 15476 18241 15494 18275
rect 15494 18241 15528 18275
rect 15476 18232 15528 18241
rect 17500 18232 17552 18284
rect 17776 18275 17828 18284
rect 17776 18241 17794 18275
rect 17794 18241 17828 18275
rect 17776 18232 17828 18241
rect 19616 18232 19668 18284
rect 20260 18275 20312 18284
rect 20260 18241 20294 18275
rect 20294 18241 20312 18275
rect 20260 18232 20312 18241
rect 18052 18207 18104 18216
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 16948 18096 17000 18148
rect 13728 18028 13780 18080
rect 13820 18028 13872 18080
rect 15568 18028 15620 18080
rect 15752 18028 15804 18080
rect 16120 18028 16172 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 2872 17824 2924 17876
rect 3884 17824 3936 17876
rect 4528 17824 4580 17876
rect 4712 17824 4764 17876
rect 5448 17867 5500 17876
rect 5448 17833 5457 17867
rect 5457 17833 5491 17867
rect 5491 17833 5500 17867
rect 5448 17824 5500 17833
rect 7104 17867 7156 17876
rect 7104 17833 7113 17867
rect 7113 17833 7147 17867
rect 7147 17833 7156 17867
rect 7104 17824 7156 17833
rect 12256 17824 12308 17876
rect 12532 17824 12584 17876
rect 5080 17756 5132 17808
rect 5264 17688 5316 17740
rect 6092 17731 6144 17740
rect 6092 17697 6101 17731
rect 6101 17697 6135 17731
rect 6135 17697 6144 17731
rect 6092 17688 6144 17697
rect 9036 17688 9088 17740
rect 9312 17688 9364 17740
rect 2688 17663 2740 17672
rect 2688 17629 2697 17663
rect 2697 17629 2731 17663
rect 2731 17629 2740 17663
rect 2688 17620 2740 17629
rect 4436 17663 4488 17672
rect 4436 17629 4445 17663
rect 4445 17629 4479 17663
rect 4479 17629 4488 17663
rect 4436 17620 4488 17629
rect 4896 17620 4948 17672
rect 8668 17620 8720 17672
rect 8760 17620 8812 17672
rect 4068 17552 4120 17604
rect 7288 17552 7340 17604
rect 8852 17552 8904 17604
rect 3608 17484 3660 17536
rect 4528 17527 4580 17536
rect 4528 17493 4537 17527
rect 4537 17493 4571 17527
rect 4571 17493 4580 17527
rect 5172 17527 5224 17536
rect 4528 17484 4580 17493
rect 5172 17493 5181 17527
rect 5181 17493 5215 17527
rect 5215 17493 5224 17527
rect 5172 17484 5224 17493
rect 5908 17527 5960 17536
rect 5908 17493 5917 17527
rect 5917 17493 5951 17527
rect 5951 17493 5960 17527
rect 5908 17484 5960 17493
rect 7932 17484 7984 17536
rect 8024 17484 8076 17536
rect 8576 17527 8628 17536
rect 8576 17493 8585 17527
rect 8585 17493 8619 17527
rect 8619 17493 8628 17527
rect 8576 17484 8628 17493
rect 8944 17527 8996 17536
rect 8944 17493 8953 17527
rect 8953 17493 8987 17527
rect 8987 17493 8996 17527
rect 8944 17484 8996 17493
rect 11244 17688 11296 17740
rect 12440 17756 12492 17808
rect 20260 17824 20312 17876
rect 10784 17620 10836 17672
rect 13728 17663 13780 17672
rect 11152 17552 11204 17604
rect 11244 17552 11296 17604
rect 12072 17552 12124 17604
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 14464 17688 14516 17740
rect 17132 17688 17184 17740
rect 19616 17731 19668 17740
rect 19616 17697 19625 17731
rect 19625 17697 19659 17731
rect 19659 17697 19668 17731
rect 19616 17688 19668 17697
rect 11888 17484 11940 17536
rect 12624 17484 12676 17536
rect 13268 17484 13320 17536
rect 14740 17552 14792 17604
rect 20720 17620 20772 17672
rect 21364 17663 21416 17672
rect 21364 17629 21373 17663
rect 21373 17629 21407 17663
rect 21407 17629 21416 17663
rect 21364 17620 21416 17629
rect 15844 17552 15896 17604
rect 14556 17484 14608 17536
rect 15292 17484 15344 17536
rect 15752 17527 15804 17536
rect 15752 17493 15761 17527
rect 15761 17493 15795 17527
rect 15795 17493 15804 17527
rect 15752 17484 15804 17493
rect 17408 17484 17460 17536
rect 20812 17552 20864 17604
rect 18052 17484 18104 17536
rect 19064 17484 19116 17536
rect 19708 17484 19760 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 2780 17280 2832 17332
rect 3608 17323 3660 17332
rect 3608 17289 3617 17323
rect 3617 17289 3651 17323
rect 3651 17289 3660 17323
rect 3608 17280 3660 17289
rect 4528 17323 4580 17332
rect 4528 17289 4537 17323
rect 4537 17289 4571 17323
rect 4571 17289 4580 17323
rect 4528 17280 4580 17289
rect 4988 17323 5040 17332
rect 4988 17289 4997 17323
rect 4997 17289 5031 17323
rect 5031 17289 5040 17323
rect 4988 17280 5040 17289
rect 5908 17280 5960 17332
rect 6828 17323 6880 17332
rect 6828 17289 6837 17323
rect 6837 17289 6871 17323
rect 6871 17289 6880 17323
rect 6828 17280 6880 17289
rect 7656 17280 7708 17332
rect 7932 17323 7984 17332
rect 7932 17289 7941 17323
rect 7941 17289 7975 17323
rect 7975 17289 7984 17323
rect 7932 17280 7984 17289
rect 8944 17280 8996 17332
rect 9036 17280 9088 17332
rect 17408 17280 17460 17332
rect 20904 17280 20956 17332
rect 21548 17280 21600 17332
rect 2688 17255 2740 17264
rect 2688 17221 2697 17255
rect 2697 17221 2731 17255
rect 2731 17221 2740 17255
rect 2688 17212 2740 17221
rect 4896 17255 4948 17264
rect 4896 17221 4905 17255
rect 4905 17221 4939 17255
rect 4939 17221 4948 17255
rect 4896 17212 4948 17221
rect 5172 17212 5224 17264
rect 2872 17144 2924 17196
rect 4160 17144 4212 17196
rect 5540 17187 5592 17196
rect 5540 17153 5549 17187
rect 5549 17153 5583 17187
rect 5583 17153 5592 17187
rect 5540 17144 5592 17153
rect 7012 17212 7064 17264
rect 8852 17212 8904 17264
rect 3332 17076 3384 17128
rect 5172 17119 5224 17128
rect 3240 17008 3292 17060
rect 5172 17085 5181 17119
rect 5181 17085 5215 17119
rect 5215 17085 5224 17119
rect 5172 17076 5224 17085
rect 5632 17076 5684 17128
rect 5908 17076 5960 17128
rect 6920 17119 6972 17128
rect 6920 17085 6929 17119
rect 6929 17085 6963 17119
rect 6963 17085 6972 17119
rect 6920 17076 6972 17085
rect 7564 17076 7616 17128
rect 8576 17144 8628 17196
rect 9496 17212 9548 17264
rect 9312 17144 9364 17196
rect 10600 17212 10652 17264
rect 11704 17212 11756 17264
rect 12348 17212 12400 17264
rect 14464 17212 14516 17264
rect 17224 17212 17276 17264
rect 19616 17212 19668 17264
rect 13360 17187 13412 17196
rect 13360 17153 13378 17187
rect 13378 17153 13412 17187
rect 13360 17144 13412 17153
rect 14280 17144 14332 17196
rect 18144 17144 18196 17196
rect 10600 17076 10652 17128
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 13728 17076 13780 17128
rect 8208 17008 8260 17060
rect 10784 17008 10836 17060
rect 11704 16940 11756 16992
rect 14372 17008 14424 17060
rect 13728 16940 13780 16992
rect 15752 17008 15804 17060
rect 21364 17119 21416 17128
rect 21364 17085 21373 17119
rect 21373 17085 21407 17119
rect 21407 17085 21416 17119
rect 21364 17076 21416 17085
rect 18696 17008 18748 17060
rect 18236 16940 18288 16992
rect 18972 16983 19024 16992
rect 18972 16949 18981 16983
rect 18981 16949 19015 16983
rect 19015 16949 19024 16983
rect 18972 16940 19024 16949
rect 19064 16940 19116 16992
rect 19524 16940 19576 16992
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1952 16779 2004 16788
rect 1952 16745 1961 16779
rect 1961 16745 1995 16779
rect 1995 16745 2004 16779
rect 1952 16736 2004 16745
rect 3056 16736 3108 16788
rect 4160 16779 4212 16788
rect 4160 16745 4169 16779
rect 4169 16745 4203 16779
rect 4203 16745 4212 16779
rect 4160 16736 4212 16745
rect 3700 16668 3752 16720
rect 4712 16736 4764 16788
rect 5172 16736 5224 16788
rect 6644 16736 6696 16788
rect 6000 16668 6052 16720
rect 7104 16668 7156 16720
rect 5080 16600 5132 16652
rect 7196 16643 7248 16652
rect 7196 16609 7205 16643
rect 7205 16609 7239 16643
rect 7239 16609 7248 16643
rect 7196 16600 7248 16609
rect 2780 16532 2832 16584
rect 2872 16532 2924 16584
rect 5816 16575 5868 16584
rect 5816 16541 5825 16575
rect 5825 16541 5859 16575
rect 5859 16541 5868 16575
rect 5816 16532 5868 16541
rect 6552 16532 6604 16584
rect 6920 16439 6972 16448
rect 6920 16405 6929 16439
rect 6929 16405 6963 16439
rect 6963 16405 6972 16439
rect 6920 16396 6972 16405
rect 7564 16396 7616 16448
rect 8024 16643 8076 16652
rect 8024 16609 8033 16643
rect 8033 16609 8067 16643
rect 8067 16609 8076 16643
rect 8024 16600 8076 16609
rect 8392 16600 8444 16652
rect 13728 16736 13780 16788
rect 8116 16532 8168 16584
rect 9680 16532 9732 16584
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 10048 16532 10100 16541
rect 10876 16575 10928 16584
rect 10876 16541 10885 16575
rect 10885 16541 10919 16575
rect 10919 16541 10928 16575
rect 10876 16532 10928 16541
rect 14004 16736 14056 16788
rect 17776 16736 17828 16788
rect 15476 16711 15528 16720
rect 15476 16677 15485 16711
rect 15485 16677 15519 16711
rect 15519 16677 15528 16711
rect 15476 16668 15528 16677
rect 19064 16600 19116 16652
rect 8208 16439 8260 16448
rect 8208 16405 8217 16439
rect 8217 16405 8251 16439
rect 8251 16405 8260 16439
rect 13820 16532 13872 16584
rect 18880 16575 18932 16584
rect 12624 16507 12676 16516
rect 12624 16473 12658 16507
rect 12658 16473 12676 16507
rect 12624 16464 12676 16473
rect 13268 16464 13320 16516
rect 14372 16507 14424 16516
rect 8208 16396 8260 16405
rect 10232 16396 10284 16448
rect 11888 16396 11940 16448
rect 12440 16396 12492 16448
rect 13728 16439 13780 16448
rect 13728 16405 13737 16439
rect 13737 16405 13771 16439
rect 13771 16405 13780 16439
rect 13728 16396 13780 16405
rect 14372 16473 14406 16507
rect 14406 16473 14424 16507
rect 14372 16464 14424 16473
rect 14464 16464 14516 16516
rect 17132 16439 17184 16448
rect 17132 16405 17141 16439
rect 17141 16405 17175 16439
rect 17175 16405 17184 16439
rect 17132 16396 17184 16405
rect 18880 16541 18889 16575
rect 18889 16541 18923 16575
rect 18923 16541 18932 16575
rect 18880 16532 18932 16541
rect 19524 16532 19576 16584
rect 20812 16532 20864 16584
rect 21364 16532 21416 16584
rect 18236 16464 18288 16516
rect 20628 16396 20680 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 2044 16192 2096 16244
rect 3332 16235 3384 16244
rect 3332 16201 3341 16235
rect 3341 16201 3375 16235
rect 3375 16201 3384 16235
rect 3332 16192 3384 16201
rect 3424 16192 3476 16244
rect 5356 16192 5408 16244
rect 6000 16192 6052 16244
rect 6920 16192 6972 16244
rect 7932 16235 7984 16244
rect 7932 16201 7941 16235
rect 7941 16201 7975 16235
rect 7975 16201 7984 16235
rect 7932 16192 7984 16201
rect 8576 16192 8628 16244
rect 9312 16192 9364 16244
rect 11888 16235 11940 16244
rect 11888 16201 11897 16235
rect 11897 16201 11931 16235
rect 11931 16201 11940 16235
rect 11888 16192 11940 16201
rect 13728 16192 13780 16244
rect 19524 16192 19576 16244
rect 2780 16167 2832 16176
rect 2780 16133 2789 16167
rect 2789 16133 2823 16167
rect 2823 16133 2832 16167
rect 3700 16167 3752 16176
rect 2780 16124 2832 16133
rect 3700 16133 3709 16167
rect 3709 16133 3743 16167
rect 3743 16133 3752 16167
rect 3700 16124 3752 16133
rect 4068 16124 4120 16176
rect 6828 16124 6880 16176
rect 1492 16056 1544 16108
rect 3332 16056 3384 16108
rect 3148 15988 3200 16040
rect 4068 15988 4120 16040
rect 5172 16056 5224 16108
rect 6276 15988 6328 16040
rect 6644 15988 6696 16040
rect 9680 16124 9732 16176
rect 9864 16124 9916 16176
rect 10692 16124 10744 16176
rect 13820 16124 13872 16176
rect 9036 16056 9088 16108
rect 10232 16099 10284 16108
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 10508 16099 10560 16108
rect 10508 16065 10517 16099
rect 10517 16065 10551 16099
rect 10551 16065 10560 16099
rect 10508 16056 10560 16065
rect 6000 15920 6052 15972
rect 7196 15920 7248 15972
rect 11336 15988 11388 16040
rect 14004 16056 14056 16108
rect 16488 16124 16540 16176
rect 18696 16167 18748 16176
rect 18696 16133 18705 16167
rect 18705 16133 18739 16167
rect 18739 16133 18748 16167
rect 18696 16124 18748 16133
rect 18972 16124 19024 16176
rect 18328 16056 18380 16108
rect 18880 16056 18932 16108
rect 3056 15852 3108 15904
rect 4988 15852 5040 15904
rect 7380 15852 7432 15904
rect 15384 15920 15436 15972
rect 16488 15920 16540 15972
rect 21088 15920 21140 15972
rect 10508 15852 10560 15904
rect 13268 15852 13320 15904
rect 14924 15895 14976 15904
rect 14924 15861 14933 15895
rect 14933 15861 14967 15895
rect 14967 15861 14976 15895
rect 14924 15852 14976 15861
rect 15108 15852 15160 15904
rect 16948 15852 17000 15904
rect 18328 15895 18380 15904
rect 18328 15861 18337 15895
rect 18337 15861 18371 15895
rect 18371 15861 18380 15895
rect 18328 15852 18380 15861
rect 20444 15895 20496 15904
rect 20444 15861 20453 15895
rect 20453 15861 20487 15895
rect 20487 15861 20496 15895
rect 20444 15852 20496 15861
rect 20812 15895 20864 15904
rect 20812 15861 20821 15895
rect 20821 15861 20855 15895
rect 20855 15861 20864 15895
rect 20812 15852 20864 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1860 15648 1912 15700
rect 2412 15648 2464 15700
rect 2964 15648 3016 15700
rect 3148 15648 3200 15700
rect 6736 15648 6788 15700
rect 7380 15691 7432 15700
rect 7380 15657 7389 15691
rect 7389 15657 7423 15691
rect 7423 15657 7432 15691
rect 7380 15648 7432 15657
rect 9404 15648 9456 15700
rect 9496 15648 9548 15700
rect 13728 15648 13780 15700
rect 14096 15648 14148 15700
rect 15844 15648 15896 15700
rect 3424 15580 3476 15632
rect 5080 15512 5132 15564
rect 2136 15487 2188 15496
rect 2136 15453 2145 15487
rect 2145 15453 2179 15487
rect 2179 15453 2188 15487
rect 2136 15444 2188 15453
rect 2688 15487 2740 15496
rect 2688 15453 2697 15487
rect 2697 15453 2731 15487
rect 2731 15453 2740 15487
rect 2688 15444 2740 15453
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 7104 15580 7156 15632
rect 6276 15555 6328 15564
rect 6276 15521 6285 15555
rect 6285 15521 6319 15555
rect 6319 15521 6328 15555
rect 6276 15512 6328 15521
rect 8024 15555 8076 15564
rect 8024 15521 8033 15555
rect 8033 15521 8067 15555
rect 8067 15521 8076 15555
rect 8668 15580 8720 15632
rect 13452 15580 13504 15632
rect 8024 15512 8076 15521
rect 5724 15444 5776 15496
rect 3424 15376 3476 15428
rect 5356 15376 5408 15428
rect 8208 15444 8260 15496
rect 5724 15308 5776 15360
rect 6644 15376 6696 15428
rect 6736 15376 6788 15428
rect 7380 15376 7432 15428
rect 8484 15444 8536 15496
rect 9588 15444 9640 15496
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 13544 15444 13596 15496
rect 13820 15444 13872 15496
rect 18328 15444 18380 15496
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 20812 15444 20864 15496
rect 6276 15308 6328 15360
rect 6920 15308 6972 15360
rect 7564 15308 7616 15360
rect 7932 15308 7984 15360
rect 8116 15351 8168 15360
rect 8116 15317 8125 15351
rect 8125 15317 8159 15351
rect 8159 15317 8168 15351
rect 8116 15308 8168 15317
rect 8668 15308 8720 15360
rect 10784 15351 10836 15360
rect 10784 15317 10793 15351
rect 10793 15317 10827 15351
rect 10827 15317 10836 15351
rect 10784 15308 10836 15317
rect 10876 15308 10928 15360
rect 11336 15308 11388 15360
rect 14096 15308 14148 15360
rect 14464 15376 14516 15428
rect 17040 15419 17092 15428
rect 17040 15385 17074 15419
rect 17074 15385 17092 15419
rect 17040 15376 17092 15385
rect 20628 15376 20680 15428
rect 16120 15308 16172 15360
rect 16396 15351 16448 15360
rect 16396 15317 16405 15351
rect 16405 15317 16439 15351
rect 16439 15317 16448 15351
rect 16396 15308 16448 15317
rect 18144 15351 18196 15360
rect 18144 15317 18153 15351
rect 18153 15317 18187 15351
rect 18187 15317 18196 15351
rect 18144 15308 18196 15317
rect 18972 15308 19024 15360
rect 19800 15308 19852 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 2872 15104 2924 15156
rect 5816 15104 5868 15156
rect 2136 15036 2188 15088
rect 3424 15036 3476 15088
rect 7104 15079 7156 15088
rect 7104 15045 7113 15079
rect 7113 15045 7147 15079
rect 7147 15045 7156 15079
rect 7104 15036 7156 15045
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 3884 14968 3936 15020
rect 5632 15011 5684 15020
rect 3332 14943 3384 14952
rect 3332 14909 3341 14943
rect 3341 14909 3375 14943
rect 3375 14909 3384 14943
rect 3332 14900 3384 14909
rect 3976 14900 4028 14952
rect 4436 14943 4488 14952
rect 4436 14909 4445 14943
rect 4445 14909 4479 14943
rect 4479 14909 4488 14943
rect 4436 14900 4488 14909
rect 5632 14977 5641 15011
rect 5641 14977 5675 15011
rect 5675 14977 5684 15011
rect 5632 14968 5684 14977
rect 6092 14900 6144 14952
rect 7012 14943 7064 14952
rect 7012 14909 7021 14943
rect 7021 14909 7055 14943
rect 7055 14909 7064 14943
rect 7012 14900 7064 14909
rect 4620 14832 4672 14884
rect 2320 14764 2372 14816
rect 6644 14832 6696 14884
rect 4988 14807 5040 14816
rect 4988 14773 4997 14807
rect 4997 14773 5031 14807
rect 5031 14773 5040 14807
rect 4988 14764 5040 14773
rect 5724 14764 5776 14816
rect 6736 14764 6788 14816
rect 7104 14764 7156 14816
rect 8024 15104 8076 15156
rect 8392 15104 8444 15156
rect 14464 15104 14516 15156
rect 8484 15036 8536 15088
rect 9956 15036 10008 15088
rect 11980 15036 12032 15088
rect 7564 14968 7616 15020
rect 8024 14968 8076 15020
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 11520 15011 11572 15020
rect 11520 14977 11529 15011
rect 11529 14977 11563 15011
rect 11563 14977 11572 15011
rect 11520 14968 11572 14977
rect 11704 14968 11756 15020
rect 13728 15036 13780 15088
rect 14280 15036 14332 15088
rect 9312 14943 9364 14952
rect 8208 14832 8260 14884
rect 9312 14909 9321 14943
rect 9321 14909 9355 14943
rect 9355 14909 9364 14943
rect 9312 14900 9364 14909
rect 8852 14875 8904 14884
rect 8852 14841 8861 14875
rect 8861 14841 8895 14875
rect 8895 14841 8904 14875
rect 8852 14832 8904 14841
rect 12992 14900 13044 14952
rect 14924 14968 14976 15020
rect 16396 15036 16448 15088
rect 17960 15011 18012 15020
rect 20812 15036 20864 15088
rect 17960 14977 17978 15011
rect 17978 14977 18012 15011
rect 17960 14968 18012 14977
rect 18328 14968 18380 15020
rect 19708 14968 19760 15020
rect 16580 14900 16632 14952
rect 14464 14832 14516 14884
rect 10692 14764 10744 14816
rect 12808 14764 12860 14816
rect 14280 14764 14332 14816
rect 14740 14764 14792 14816
rect 17960 14764 18012 14816
rect 18328 14764 18380 14816
rect 19800 14764 19852 14816
rect 19984 14807 20036 14816
rect 19984 14773 19993 14807
rect 19993 14773 20027 14807
rect 20027 14773 20036 14807
rect 19984 14764 20036 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 2504 14560 2556 14612
rect 3976 14603 4028 14612
rect 3976 14569 3985 14603
rect 3985 14569 4019 14603
rect 4019 14569 4028 14603
rect 3976 14560 4028 14569
rect 4160 14560 4212 14612
rect 5448 14603 5500 14612
rect 3516 14492 3568 14544
rect 4252 14492 4304 14544
rect 4436 14492 4488 14544
rect 2228 14356 2280 14408
rect 3332 14356 3384 14408
rect 3700 14356 3752 14408
rect 2504 14288 2556 14340
rect 3148 14288 3200 14340
rect 3332 14263 3384 14272
rect 3332 14229 3341 14263
rect 3341 14229 3375 14263
rect 3375 14229 3384 14263
rect 3332 14220 3384 14229
rect 4252 14288 4304 14340
rect 5448 14569 5457 14603
rect 5457 14569 5491 14603
rect 5491 14569 5500 14603
rect 5448 14560 5500 14569
rect 5816 14560 5868 14612
rect 7656 14560 7708 14612
rect 8392 14560 8444 14612
rect 9312 14560 9364 14612
rect 4988 14492 5040 14544
rect 10876 14560 10928 14612
rect 11520 14560 11572 14612
rect 15844 14603 15896 14612
rect 15844 14569 15853 14603
rect 15853 14569 15887 14603
rect 15887 14569 15896 14603
rect 15844 14560 15896 14569
rect 19708 14560 19760 14612
rect 7656 14424 7708 14476
rect 8024 14424 8076 14476
rect 8300 14467 8352 14476
rect 8300 14433 8309 14467
rect 8309 14433 8343 14467
rect 8343 14433 8352 14467
rect 8300 14424 8352 14433
rect 9128 14424 9180 14476
rect 13820 14492 13872 14544
rect 16580 14535 16632 14544
rect 16580 14501 16589 14535
rect 16589 14501 16623 14535
rect 16623 14501 16632 14535
rect 16580 14492 16632 14501
rect 17960 14492 18012 14544
rect 10692 14467 10744 14476
rect 5356 14356 5408 14408
rect 7564 14356 7616 14408
rect 8484 14356 8536 14408
rect 9312 14399 9364 14408
rect 9312 14365 9321 14399
rect 9321 14365 9355 14399
rect 9355 14365 9364 14399
rect 9312 14356 9364 14365
rect 10692 14433 10701 14467
rect 10701 14433 10735 14467
rect 10735 14433 10744 14467
rect 10692 14424 10744 14433
rect 19708 14424 19760 14476
rect 20168 14424 20220 14476
rect 13544 14356 13596 14408
rect 13728 14356 13780 14408
rect 15016 14356 15068 14408
rect 4620 14220 4672 14272
rect 6828 14220 6880 14272
rect 7012 14220 7064 14272
rect 10784 14263 10836 14272
rect 10784 14229 10793 14263
rect 10793 14229 10827 14263
rect 10827 14229 10836 14263
rect 10784 14220 10836 14229
rect 10876 14263 10928 14272
rect 10876 14229 10885 14263
rect 10885 14229 10919 14263
rect 10919 14229 10928 14263
rect 13728 14263 13780 14272
rect 10876 14220 10928 14229
rect 13728 14229 13737 14263
rect 13737 14229 13771 14263
rect 13771 14229 13780 14263
rect 13728 14220 13780 14229
rect 14556 14288 14608 14340
rect 17408 14288 17460 14340
rect 17684 14331 17736 14340
rect 17684 14297 17702 14331
rect 17702 14297 17736 14331
rect 17684 14288 17736 14297
rect 16580 14220 16632 14272
rect 17316 14220 17368 14272
rect 18236 14220 18288 14272
rect 18696 14220 18748 14272
rect 20444 14288 20496 14340
rect 20812 14288 20864 14340
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 1400 14016 1452 14068
rect 3516 14016 3568 14068
rect 4252 14059 4304 14068
rect 4252 14025 4261 14059
rect 4261 14025 4295 14059
rect 4295 14025 4304 14059
rect 4252 14016 4304 14025
rect 4804 14016 4856 14068
rect 5540 14016 5592 14068
rect 7012 14016 7064 14068
rect 7104 14016 7156 14068
rect 8116 14016 8168 14068
rect 8576 14016 8628 14068
rect 9128 14016 9180 14068
rect 9312 14016 9364 14068
rect 10048 14016 10100 14068
rect 10876 14059 10928 14068
rect 10876 14025 10885 14059
rect 10885 14025 10919 14059
rect 10919 14025 10928 14059
rect 10876 14016 10928 14025
rect 13544 14016 13596 14068
rect 2320 13855 2372 13864
rect 1860 13744 1912 13796
rect 2320 13821 2329 13855
rect 2329 13821 2363 13855
rect 2363 13821 2372 13855
rect 2320 13812 2372 13821
rect 4160 13880 4212 13932
rect 2412 13676 2464 13728
rect 3332 13744 3384 13796
rect 3700 13812 3752 13864
rect 4804 13812 4856 13864
rect 4068 13744 4120 13796
rect 4712 13744 4764 13796
rect 5172 13812 5224 13864
rect 10968 13948 11020 14000
rect 12532 13948 12584 14000
rect 8392 13880 8444 13932
rect 9680 13880 9732 13932
rect 10048 13880 10100 13932
rect 10232 13923 10284 13932
rect 10232 13889 10241 13923
rect 10241 13889 10275 13923
rect 10275 13889 10284 13923
rect 10232 13880 10284 13889
rect 13452 13880 13504 13932
rect 14464 13880 14516 13932
rect 14924 14016 14976 14068
rect 17040 14016 17092 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 17684 14016 17736 14068
rect 19800 14016 19852 14068
rect 20720 14059 20772 14068
rect 15016 13948 15068 14000
rect 20720 14025 20729 14059
rect 20729 14025 20763 14059
rect 20763 14025 20772 14059
rect 20720 14016 20772 14025
rect 20168 13923 20220 13932
rect 20168 13889 20186 13923
rect 20186 13889 20220 13923
rect 20168 13880 20220 13889
rect 20812 13880 20864 13932
rect 5448 13744 5500 13796
rect 7840 13812 7892 13864
rect 10324 13855 10376 13864
rect 4620 13719 4672 13728
rect 4620 13685 4629 13719
rect 4629 13685 4663 13719
rect 4663 13685 4672 13719
rect 4620 13676 4672 13685
rect 5080 13676 5132 13728
rect 7104 13744 7156 13796
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 12256 13812 12308 13864
rect 13728 13812 13780 13864
rect 9496 13744 9548 13796
rect 6920 13676 6972 13728
rect 8392 13676 8444 13728
rect 12256 13676 12308 13728
rect 15476 13676 15528 13728
rect 18052 13676 18104 13728
rect 19064 13719 19116 13728
rect 19064 13685 19073 13719
rect 19073 13685 19107 13719
rect 19107 13685 19116 13719
rect 19064 13676 19116 13685
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 2320 13472 2372 13524
rect 3884 13472 3936 13524
rect 4068 13472 4120 13524
rect 4528 13472 4580 13524
rect 6000 13472 6052 13524
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 8576 13472 8628 13524
rect 9312 13515 9364 13524
rect 9312 13481 9321 13515
rect 9321 13481 9355 13515
rect 9355 13481 9364 13515
rect 9312 13472 9364 13481
rect 10416 13472 10468 13524
rect 4436 13404 4488 13456
rect 6552 13404 6604 13456
rect 1400 13336 1452 13388
rect 2412 13336 2464 13388
rect 3332 13379 3384 13388
rect 3332 13345 3341 13379
rect 3341 13345 3375 13379
rect 3375 13345 3384 13379
rect 3332 13336 3384 13345
rect 3516 13336 3568 13388
rect 4252 13336 4304 13388
rect 5172 13379 5224 13388
rect 5172 13345 5181 13379
rect 5181 13345 5215 13379
rect 5215 13345 5224 13379
rect 5172 13336 5224 13345
rect 5356 13379 5408 13388
rect 5356 13345 5365 13379
rect 5365 13345 5399 13379
rect 5399 13345 5408 13379
rect 5356 13336 5408 13345
rect 3148 13268 3200 13320
rect 4620 13268 4672 13320
rect 6552 13268 6604 13320
rect 7196 13404 7248 13456
rect 8392 13336 8444 13388
rect 9956 13336 10008 13388
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 13176 13472 13228 13524
rect 13912 13472 13964 13524
rect 14740 13472 14792 13524
rect 15292 13472 15344 13524
rect 17040 13472 17092 13524
rect 19524 13515 19576 13524
rect 19524 13481 19533 13515
rect 19533 13481 19567 13515
rect 19567 13481 19576 13515
rect 19524 13472 19576 13481
rect 20168 13472 20220 13524
rect 18880 13447 18932 13456
rect 18880 13413 18889 13447
rect 18889 13413 18923 13447
rect 18923 13413 18932 13447
rect 18880 13404 18932 13413
rect 12164 13311 12216 13320
rect 2412 13200 2464 13252
rect 5264 13200 5316 13252
rect 10600 13200 10652 13252
rect 10968 13200 11020 13252
rect 1860 13132 1912 13184
rect 3976 13132 4028 13184
rect 4252 13132 4304 13184
rect 4528 13132 4580 13184
rect 6828 13175 6880 13184
rect 6828 13141 6837 13175
rect 6837 13141 6871 13175
rect 6871 13141 6880 13175
rect 6828 13132 6880 13141
rect 7656 13132 7708 13184
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 12164 13268 12216 13277
rect 13728 13268 13780 13320
rect 18052 13268 18104 13320
rect 20812 13268 20864 13320
rect 12256 13200 12308 13252
rect 13636 13200 13688 13252
rect 13084 13132 13136 13184
rect 13360 13132 13412 13184
rect 14464 13200 14516 13252
rect 19340 13200 19392 13252
rect 19984 13200 20036 13252
rect 20076 13200 20128 13252
rect 21088 13200 21140 13252
rect 19616 13132 19668 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 3148 12928 3200 12980
rect 5264 12971 5316 12980
rect 5264 12937 5273 12971
rect 5273 12937 5307 12971
rect 5307 12937 5316 12971
rect 5264 12928 5316 12937
rect 5356 12928 5408 12980
rect 7288 12928 7340 12980
rect 2596 12860 2648 12912
rect 3976 12860 4028 12912
rect 6644 12860 6696 12912
rect 9220 12928 9272 12980
rect 10600 12971 10652 12980
rect 10600 12937 10609 12971
rect 10609 12937 10643 12971
rect 10643 12937 10652 12971
rect 10600 12928 10652 12937
rect 11152 12928 11204 12980
rect 11980 12928 12032 12980
rect 12440 12928 12492 12980
rect 13452 12928 13504 12980
rect 19340 12971 19392 12980
rect 19340 12937 19349 12971
rect 19349 12937 19383 12971
rect 19383 12937 19392 12971
rect 19340 12928 19392 12937
rect 19800 12971 19852 12980
rect 19800 12937 19809 12971
rect 19809 12937 19843 12971
rect 19843 12937 19852 12971
rect 19800 12928 19852 12937
rect 7840 12860 7892 12912
rect 14464 12860 14516 12912
rect 14740 12860 14792 12912
rect 18880 12860 18932 12912
rect 2320 12792 2372 12844
rect 2412 12792 2464 12844
rect 3332 12835 3384 12844
rect 3332 12801 3341 12835
rect 3341 12801 3375 12835
rect 3375 12801 3384 12835
rect 3332 12792 3384 12801
rect 6276 12792 6328 12844
rect 8024 12835 8076 12844
rect 8024 12801 8033 12835
rect 8033 12801 8067 12835
rect 8067 12801 8076 12835
rect 8024 12792 8076 12801
rect 8576 12792 8628 12844
rect 9220 12792 9272 12844
rect 3056 12724 3108 12776
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4436 12724 4488 12733
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 6460 12767 6512 12776
rect 6460 12733 6469 12767
rect 6469 12733 6503 12767
rect 6503 12733 6512 12767
rect 6460 12724 6512 12733
rect 6644 12767 6696 12776
rect 6644 12733 6653 12767
rect 6653 12733 6687 12767
rect 6687 12733 6696 12767
rect 6644 12724 6696 12733
rect 8208 12767 8260 12776
rect 8208 12733 8217 12767
rect 8217 12733 8251 12767
rect 8251 12733 8260 12767
rect 8208 12724 8260 12733
rect 9588 12724 9640 12776
rect 9956 12724 10008 12776
rect 11980 12767 12032 12776
rect 1860 12588 1912 12640
rect 3148 12588 3200 12640
rect 3516 12588 3568 12640
rect 7840 12588 7892 12640
rect 10784 12656 10836 12708
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 12256 12724 12308 12776
rect 13912 12792 13964 12844
rect 14556 12792 14608 12844
rect 16948 12792 17000 12844
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 12164 12588 12216 12640
rect 12900 12588 12952 12640
rect 13728 12588 13780 12640
rect 21272 12724 21324 12776
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 4160 12384 4212 12436
rect 5632 12384 5684 12436
rect 4068 12316 4120 12368
rect 2228 12291 2280 12300
rect 2228 12257 2237 12291
rect 2237 12257 2271 12291
rect 2271 12257 2280 12291
rect 2228 12248 2280 12257
rect 3148 12248 3200 12300
rect 3792 12248 3844 12300
rect 4620 12248 4672 12300
rect 4804 12248 4856 12300
rect 4988 12291 5040 12300
rect 4988 12257 4997 12291
rect 4997 12257 5031 12291
rect 5031 12257 5040 12291
rect 4988 12248 5040 12257
rect 2412 12223 2464 12232
rect 2412 12189 2421 12223
rect 2421 12189 2455 12223
rect 2455 12189 2464 12223
rect 2412 12180 2464 12189
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 4436 12180 4488 12232
rect 9220 12384 9272 12436
rect 9772 12384 9824 12436
rect 11796 12384 11848 12436
rect 11980 12384 12032 12436
rect 16396 12384 16448 12436
rect 19248 12384 19300 12436
rect 6276 12291 6328 12300
rect 6276 12257 6285 12291
rect 6285 12257 6319 12291
rect 6319 12257 6328 12291
rect 6276 12248 6328 12257
rect 3884 12112 3936 12164
rect 6644 12112 6696 12164
rect 7012 12112 7064 12164
rect 8024 12248 8076 12300
rect 10692 12316 10744 12368
rect 10324 12180 10376 12232
rect 11796 12248 11848 12300
rect 14464 12248 14516 12300
rect 14648 12248 14700 12300
rect 12440 12180 12492 12232
rect 13084 12180 13136 12232
rect 3148 12044 3200 12096
rect 5080 12087 5132 12096
rect 5080 12053 5089 12087
rect 5089 12053 5123 12087
rect 5123 12053 5132 12087
rect 5080 12044 5132 12053
rect 6736 12044 6788 12096
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 12716 12112 12768 12164
rect 13452 12155 13504 12164
rect 13452 12121 13470 12155
rect 13470 12121 13504 12155
rect 13452 12112 13504 12121
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 16120 12180 16172 12232
rect 19064 12180 19116 12232
rect 21272 12180 21324 12232
rect 15292 12155 15344 12164
rect 8116 12044 8168 12096
rect 9312 12087 9364 12096
rect 9312 12053 9321 12087
rect 9321 12053 9355 12087
rect 9355 12053 9364 12087
rect 9312 12044 9364 12053
rect 9956 12044 10008 12096
rect 11704 12087 11756 12096
rect 11704 12053 11713 12087
rect 11713 12053 11747 12087
rect 11747 12053 11756 12087
rect 11704 12044 11756 12053
rect 12164 12044 12216 12096
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 15292 12121 15326 12155
rect 15326 12121 15344 12155
rect 15292 12112 15344 12121
rect 21088 12155 21140 12164
rect 21088 12121 21106 12155
rect 21106 12121 21140 12155
rect 21088 12112 21140 12121
rect 18512 12087 18564 12096
rect 18512 12053 18521 12087
rect 18521 12053 18555 12087
rect 18555 12053 18564 12087
rect 18512 12044 18564 12053
rect 18880 12044 18932 12096
rect 20444 12044 20496 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 2964 11840 3016 11892
rect 3148 11883 3200 11892
rect 3148 11849 3157 11883
rect 3157 11849 3191 11883
rect 3191 11849 3200 11883
rect 3148 11840 3200 11849
rect 388 11772 440 11824
rect 3976 11840 4028 11892
rect 5080 11840 5132 11892
rect 6644 11840 6696 11892
rect 7196 11840 7248 11892
rect 7288 11772 7340 11824
rect 9312 11840 9364 11892
rect 10876 11883 10928 11892
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 19616 11883 19668 11892
rect 9956 11772 10008 11824
rect 10048 11772 10100 11824
rect 13728 11815 13780 11824
rect 13728 11781 13737 11815
rect 13737 11781 13771 11815
rect 13771 11781 13780 11815
rect 13728 11772 13780 11781
rect 19616 11849 19625 11883
rect 19625 11849 19659 11883
rect 19659 11849 19668 11883
rect 19616 11840 19668 11849
rect 21088 11840 21140 11892
rect 2320 11636 2372 11688
rect 3148 11636 3200 11688
rect 4528 11636 4580 11688
rect 5448 11679 5500 11688
rect 5448 11645 5457 11679
rect 5457 11645 5491 11679
rect 5491 11645 5500 11679
rect 5448 11636 5500 11645
rect 7840 11704 7892 11756
rect 12716 11704 12768 11756
rect 13360 11704 13412 11756
rect 15752 11772 15804 11824
rect 17224 11772 17276 11824
rect 18788 11815 18840 11824
rect 18788 11781 18806 11815
rect 18806 11781 18840 11815
rect 18788 11772 18840 11781
rect 15108 11704 15160 11756
rect 16304 11704 16356 11756
rect 19064 11747 19116 11756
rect 10048 11679 10100 11688
rect 10048 11645 10057 11679
rect 10057 11645 10091 11679
rect 10091 11645 10100 11679
rect 10048 11636 10100 11645
rect 12348 11636 12400 11688
rect 16120 11636 16172 11688
rect 19064 11713 19073 11747
rect 19073 11713 19107 11747
rect 19107 11713 19116 11747
rect 19064 11704 19116 11713
rect 20444 11704 20496 11756
rect 21272 11704 21324 11756
rect 3056 11500 3108 11552
rect 4068 11500 4120 11552
rect 4252 11500 4304 11552
rect 5908 11500 5960 11552
rect 6736 11500 6788 11552
rect 12072 11543 12124 11552
rect 12072 11509 12081 11543
rect 12081 11509 12115 11543
rect 12115 11509 12124 11543
rect 12072 11500 12124 11509
rect 14740 11500 14792 11552
rect 16120 11500 16172 11552
rect 16304 11500 16356 11552
rect 18420 11500 18472 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 2780 11296 2832 11348
rect 4436 11296 4488 11348
rect 5172 11296 5224 11348
rect 5448 11296 5500 11348
rect 8116 11296 8168 11348
rect 8668 11296 8720 11348
rect 4160 11228 4212 11280
rect 13452 11296 13504 11348
rect 14832 11296 14884 11348
rect 1492 11160 1544 11212
rect 5632 11160 5684 11212
rect 6184 11203 6236 11212
rect 4068 11092 4120 11144
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 4344 11092 4396 11144
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 6736 11160 6788 11212
rect 9496 11203 9548 11212
rect 9496 11169 9505 11203
rect 9505 11169 9539 11203
rect 9539 11169 9548 11203
rect 9496 11160 9548 11169
rect 10140 11160 10192 11212
rect 12348 11271 12400 11280
rect 12348 11237 12357 11271
rect 12357 11237 12391 11271
rect 12391 11237 12400 11271
rect 12348 11228 12400 11237
rect 15200 11296 15252 11348
rect 15476 11339 15528 11348
rect 15476 11305 15485 11339
rect 15485 11305 15519 11339
rect 15519 11305 15528 11339
rect 15476 11296 15528 11305
rect 18788 11296 18840 11348
rect 19616 11296 19668 11348
rect 20812 11296 20864 11348
rect 21272 11339 21324 11348
rect 21272 11305 21281 11339
rect 21281 11305 21315 11339
rect 21315 11305 21324 11339
rect 21272 11296 21324 11305
rect 15752 11271 15804 11280
rect 15752 11237 15761 11271
rect 15761 11237 15795 11271
rect 15795 11237 15804 11271
rect 15752 11228 15804 11237
rect 12716 11160 12768 11212
rect 13728 11203 13780 11212
rect 13728 11169 13737 11203
rect 13737 11169 13771 11203
rect 13771 11169 13780 11203
rect 13728 11160 13780 11169
rect 19064 11160 19116 11212
rect 7472 11135 7524 11144
rect 5172 11092 5224 11101
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 9128 11092 9180 11144
rect 10048 11092 10100 11144
rect 13176 11092 13228 11144
rect 14372 11135 14424 11144
rect 14372 11101 14406 11135
rect 14406 11101 14424 11135
rect 14372 11092 14424 11101
rect 16120 11092 16172 11144
rect 19524 11092 19576 11144
rect 3516 11024 3568 11076
rect 4988 11024 5040 11076
rect 9496 11024 9548 11076
rect 5816 10956 5868 11008
rect 9128 10956 9180 11008
rect 10232 10999 10284 11008
rect 10232 10965 10241 10999
rect 10241 10965 10275 10999
rect 10275 10965 10284 10999
rect 10232 10956 10284 10965
rect 10324 10956 10376 11008
rect 14280 11024 14332 11076
rect 17040 11024 17092 11076
rect 17316 11024 17368 11076
rect 18328 10956 18380 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 1768 10752 1820 10804
rect 4344 10752 4396 10804
rect 4620 10795 4672 10804
rect 4620 10761 4629 10795
rect 4629 10761 4663 10795
rect 4663 10761 4672 10795
rect 4620 10752 4672 10761
rect 6736 10795 6788 10804
rect 6736 10761 6745 10795
rect 6745 10761 6779 10795
rect 6779 10761 6788 10795
rect 6736 10752 6788 10761
rect 9772 10752 9824 10804
rect 10232 10752 10284 10804
rect 12992 10795 13044 10804
rect 12992 10761 13001 10795
rect 13001 10761 13035 10795
rect 13035 10761 13044 10795
rect 12992 10752 13044 10761
rect 2688 10684 2740 10736
rect 4068 10684 4120 10736
rect 1492 10616 1544 10668
rect 2872 10659 2924 10668
rect 2872 10625 2881 10659
rect 2881 10625 2915 10659
rect 2915 10625 2924 10659
rect 2872 10616 2924 10625
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 4160 10616 4212 10668
rect 7012 10684 7064 10736
rect 8484 10684 8536 10736
rect 15384 10752 15436 10804
rect 19708 10795 19760 10804
rect 19708 10761 19717 10795
rect 19717 10761 19751 10795
rect 19751 10761 19760 10795
rect 19708 10752 19760 10761
rect 20076 10752 20128 10804
rect 8392 10616 8444 10668
rect 13820 10616 13872 10668
rect 14280 10616 14332 10668
rect 14740 10684 14792 10736
rect 2504 10548 2556 10600
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 8024 10591 8076 10600
rect 6552 10548 6604 10557
rect 8024 10557 8033 10591
rect 8033 10557 8067 10591
rect 8067 10557 8076 10591
rect 8024 10548 8076 10557
rect 9312 10548 9364 10600
rect 12072 10548 12124 10600
rect 6736 10480 6788 10532
rect 16120 10548 16172 10600
rect 17224 10616 17276 10668
rect 18420 10684 18472 10736
rect 21088 10659 21140 10668
rect 21088 10625 21106 10659
rect 21106 10625 21140 10659
rect 21088 10616 21140 10625
rect 21272 10616 21324 10668
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 7288 10412 7340 10464
rect 9128 10412 9180 10464
rect 9956 10412 10008 10464
rect 15292 10412 15344 10464
rect 15752 10412 15804 10464
rect 17868 10412 17920 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 2044 10251 2096 10260
rect 2044 10217 2053 10251
rect 2053 10217 2087 10251
rect 2087 10217 2096 10251
rect 2044 10208 2096 10217
rect 2872 10208 2924 10260
rect 5632 10208 5684 10260
rect 6828 10251 6880 10260
rect 6828 10217 6837 10251
rect 6837 10217 6871 10251
rect 6871 10217 6880 10251
rect 6828 10208 6880 10217
rect 7472 10208 7524 10260
rect 8208 10208 8260 10260
rect 9496 10208 9548 10260
rect 9680 10251 9732 10260
rect 9680 10217 9689 10251
rect 9689 10217 9723 10251
rect 9723 10217 9732 10251
rect 9680 10208 9732 10217
rect 3424 10140 3476 10192
rect 5724 10140 5776 10192
rect 6552 10140 6604 10192
rect 7196 10140 7248 10192
rect 5540 10072 5592 10124
rect 9956 10140 10008 10192
rect 8484 10115 8536 10124
rect 8484 10081 8493 10115
rect 8493 10081 8527 10115
rect 8527 10081 8536 10115
rect 8484 10072 8536 10081
rect 9404 10072 9456 10124
rect 9588 10072 9640 10124
rect 14372 10208 14424 10260
rect 15752 10251 15804 10260
rect 15752 10217 15761 10251
rect 15761 10217 15795 10251
rect 15795 10217 15804 10251
rect 15752 10208 15804 10217
rect 18604 10208 18656 10260
rect 13820 10140 13872 10192
rect 4988 10004 5040 10056
rect 9312 10047 9364 10056
rect 9312 10013 9321 10047
rect 9321 10013 9355 10047
rect 9355 10013 9364 10047
rect 9312 10004 9364 10013
rect 12348 10004 12400 10056
rect 13912 10004 13964 10056
rect 16120 10004 16172 10056
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 19616 10208 19668 10260
rect 19064 10004 19116 10056
rect 6000 9936 6052 9988
rect 7104 9936 7156 9988
rect 9220 9979 9272 9988
rect 9220 9945 9229 9979
rect 9229 9945 9263 9979
rect 9263 9945 9272 9979
rect 9220 9936 9272 9945
rect 10048 9936 10100 9988
rect 15200 9979 15252 9988
rect 4620 9911 4672 9920
rect 4620 9877 4629 9911
rect 4629 9877 4663 9911
rect 4663 9877 4672 9911
rect 4620 9868 4672 9877
rect 5816 9911 5868 9920
rect 5816 9877 5825 9911
rect 5825 9877 5859 9911
rect 5859 9877 5868 9911
rect 5816 9868 5868 9877
rect 6920 9868 6972 9920
rect 7840 9868 7892 9920
rect 8300 9911 8352 9920
rect 8300 9877 8309 9911
rect 8309 9877 8343 9911
rect 8343 9877 8352 9911
rect 8300 9868 8352 9877
rect 8576 9868 8628 9920
rect 9496 9868 9548 9920
rect 10784 9868 10836 9920
rect 10876 9868 10928 9920
rect 14096 9868 14148 9920
rect 15200 9945 15218 9979
rect 15218 9945 15252 9979
rect 15200 9936 15252 9945
rect 16764 9868 16816 9920
rect 17868 9936 17920 9988
rect 19800 9936 19852 9988
rect 20720 10004 20772 10056
rect 21272 10004 21324 10056
rect 16948 9868 17000 9920
rect 21364 9911 21416 9920
rect 21364 9877 21373 9911
rect 21373 9877 21407 9911
rect 21407 9877 21416 9911
rect 21364 9868 21416 9877
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 6000 9664 6052 9716
rect 7840 9707 7892 9716
rect 7840 9673 7849 9707
rect 7849 9673 7883 9707
rect 7883 9673 7892 9707
rect 7840 9664 7892 9673
rect 8300 9664 8352 9716
rect 10784 9707 10836 9716
rect 10784 9673 10793 9707
rect 10793 9673 10827 9707
rect 10827 9673 10836 9707
rect 10784 9664 10836 9673
rect 13912 9707 13964 9716
rect 13912 9673 13921 9707
rect 13921 9673 13955 9707
rect 13955 9673 13964 9707
rect 13912 9664 13964 9673
rect 16120 9664 16172 9716
rect 17224 9664 17276 9716
rect 17408 9664 17460 9716
rect 19800 9707 19852 9716
rect 19800 9673 19809 9707
rect 19809 9673 19843 9707
rect 19843 9673 19852 9707
rect 19800 9664 19852 9673
rect 20720 9664 20772 9716
rect 7104 9639 7156 9648
rect 7104 9605 7113 9639
rect 7113 9605 7147 9639
rect 7147 9605 7156 9639
rect 7104 9596 7156 9605
rect 8024 9596 8076 9648
rect 2780 9528 2832 9580
rect 4528 9571 4580 9580
rect 4528 9537 4537 9571
rect 4537 9537 4571 9571
rect 4571 9537 4580 9571
rect 4528 9528 4580 9537
rect 7380 9528 7432 9580
rect 9588 9528 9640 9580
rect 2320 9460 2372 9512
rect 5172 9460 5224 9512
rect 6920 9460 6972 9512
rect 7104 9460 7156 9512
rect 7288 9503 7340 9512
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 9036 9503 9088 9512
rect 2964 9392 3016 9444
rect 4068 9392 4120 9444
rect 5816 9392 5868 9444
rect 8392 9435 8444 9444
rect 8392 9401 8401 9435
rect 8401 9401 8435 9435
rect 8435 9401 8444 9435
rect 8392 9392 8444 9401
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 12440 9596 12492 9648
rect 12992 9596 13044 9648
rect 10784 9528 10836 9580
rect 18420 9596 18472 9648
rect 19524 9639 19576 9648
rect 19524 9605 19533 9639
rect 19533 9605 19567 9639
rect 19567 9605 19576 9639
rect 19524 9596 19576 9605
rect 20536 9639 20588 9648
rect 20536 9605 20545 9639
rect 20545 9605 20579 9639
rect 20579 9605 20588 9639
rect 20536 9596 20588 9605
rect 10048 9503 10100 9512
rect 9680 9392 9732 9444
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 10048 9460 10100 9469
rect 10692 9460 10744 9512
rect 10968 9503 11020 9512
rect 10968 9469 10977 9503
rect 10977 9469 11011 9503
rect 11011 9469 11020 9503
rect 10968 9460 11020 9469
rect 1676 9324 1728 9376
rect 3976 9324 4028 9376
rect 5908 9324 5960 9376
rect 7196 9324 7248 9376
rect 10876 9324 10928 9376
rect 15844 9435 15896 9444
rect 15844 9401 15853 9435
rect 15853 9401 15887 9435
rect 15887 9401 15896 9435
rect 15844 9392 15896 9401
rect 16948 9392 17000 9444
rect 16120 9367 16172 9376
rect 16120 9333 16129 9367
rect 16129 9333 16163 9367
rect 16163 9333 16172 9367
rect 16120 9324 16172 9333
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 2136 9163 2188 9172
rect 2136 9129 2145 9163
rect 2145 9129 2179 9163
rect 2179 9129 2188 9163
rect 2136 9120 2188 9129
rect 4528 9163 4580 9172
rect 4528 9129 4537 9163
rect 4537 9129 4571 9163
rect 4571 9129 4580 9163
rect 4528 9120 4580 9129
rect 6920 9120 6972 9172
rect 8024 9163 8076 9172
rect 8024 9129 8033 9163
rect 8033 9129 8067 9163
rect 8067 9129 8076 9163
rect 8024 9120 8076 9129
rect 9588 9163 9640 9172
rect 9588 9129 9597 9163
rect 9597 9129 9631 9163
rect 9631 9129 9640 9163
rect 9588 9120 9640 9129
rect 9680 9120 9732 9172
rect 10968 9120 11020 9172
rect 13268 9120 13320 9172
rect 19064 9120 19116 9172
rect 3976 9052 4028 9104
rect 9128 9052 9180 9104
rect 5172 9027 5224 9036
rect 5172 8993 5181 9027
rect 5181 8993 5215 9027
rect 5215 8993 5224 9027
rect 5172 8984 5224 8993
rect 5632 8984 5684 9036
rect 6644 8984 6696 9036
rect 9864 8984 9916 9036
rect 14924 9052 14976 9104
rect 12532 8984 12584 9036
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 6000 8916 6052 8968
rect 8024 8916 8076 8968
rect 10784 8916 10836 8968
rect 7288 8848 7340 8900
rect 8208 8848 8260 8900
rect 6920 8780 6972 8832
rect 7196 8780 7248 8832
rect 9404 8780 9456 8832
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 12072 8823 12124 8832
rect 12072 8789 12081 8823
rect 12081 8789 12115 8823
rect 12115 8789 12124 8823
rect 12072 8780 12124 8789
rect 16120 8780 16172 8832
rect 21272 8848 21324 8900
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 4712 8576 4764 8628
rect 7380 8619 7432 8628
rect 7380 8585 7389 8619
rect 7389 8585 7423 8619
rect 7423 8585 7432 8619
rect 7380 8576 7432 8585
rect 8576 8576 8628 8628
rect 9404 8619 9456 8628
rect 9404 8585 9413 8619
rect 9413 8585 9447 8619
rect 9447 8585 9456 8619
rect 9404 8576 9456 8585
rect 9772 8576 9824 8628
rect 10968 8576 11020 8628
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 21088 8576 21140 8628
rect 21272 8619 21324 8628
rect 21272 8585 21281 8619
rect 21281 8585 21315 8619
rect 21315 8585 21324 8619
rect 21272 8576 21324 8585
rect 5632 8551 5684 8560
rect 5632 8517 5641 8551
rect 5641 8517 5675 8551
rect 5675 8517 5684 8551
rect 5632 8508 5684 8517
rect 8668 8508 8720 8560
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 8392 8440 8444 8492
rect 5540 8372 5592 8424
rect 7104 8372 7156 8424
rect 7932 8372 7984 8424
rect 8116 8372 8168 8424
rect 8208 8372 8260 8424
rect 10140 8440 10192 8492
rect 10048 8372 10100 8424
rect 10876 8372 10928 8424
rect 12256 8508 12308 8560
rect 11704 8440 11756 8492
rect 6368 8279 6420 8288
rect 6368 8245 6377 8279
rect 6377 8245 6411 8279
rect 6411 8245 6420 8279
rect 6368 8236 6420 8245
rect 8024 8236 8076 8288
rect 9956 8304 10008 8356
rect 10692 8304 10744 8356
rect 12072 8304 12124 8356
rect 13268 8372 13320 8424
rect 18512 8508 18564 8560
rect 10324 8236 10376 8288
rect 15016 8236 15068 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 6000 8075 6052 8084
rect 6000 8041 6009 8075
rect 6009 8041 6043 8075
rect 6043 8041 6052 8075
rect 6000 8032 6052 8041
rect 8668 8032 8720 8084
rect 10048 8032 10100 8084
rect 11060 8032 11112 8084
rect 13268 8075 13320 8084
rect 4620 7964 4672 8016
rect 8116 7964 8168 8016
rect 10324 7964 10376 8016
rect 11152 7964 11204 8016
rect 11704 7964 11756 8016
rect 11888 8007 11940 8016
rect 11888 7973 11897 8007
rect 11897 7973 11931 8007
rect 11931 7973 11940 8007
rect 11888 7964 11940 7973
rect 6368 7896 6420 7948
rect 6644 7939 6696 7948
rect 6644 7905 6653 7939
rect 6653 7905 6687 7939
rect 6687 7905 6696 7939
rect 6644 7896 6696 7905
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 8208 7896 8260 7948
rect 9588 7939 9640 7948
rect 9588 7905 9597 7939
rect 9597 7905 9631 7939
rect 9631 7905 9640 7939
rect 9588 7896 9640 7905
rect 6736 7828 6788 7880
rect 10140 7828 10192 7880
rect 13268 8041 13277 8075
rect 13277 8041 13311 8075
rect 13311 8041 13320 8075
rect 13268 8032 13320 8041
rect 12532 7828 12584 7880
rect 5540 7692 5592 7744
rect 7012 7692 7064 7744
rect 9404 7735 9456 7744
rect 9404 7701 9413 7735
rect 9413 7701 9447 7735
rect 9447 7701 9456 7735
rect 9404 7692 9456 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 6644 7488 6696 7540
rect 7012 7531 7064 7540
rect 7012 7497 7021 7531
rect 7021 7497 7055 7531
rect 7055 7497 7064 7531
rect 7012 7488 7064 7497
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 8392 7531 8444 7540
rect 8392 7497 8401 7531
rect 8401 7497 8435 7531
rect 8435 7497 8444 7531
rect 8392 7488 8444 7497
rect 9588 7488 9640 7540
rect 18696 7488 18748 7540
rect 7104 7420 7156 7472
rect 5724 7352 5776 7404
rect 10324 7420 10376 7472
rect 9128 7352 9180 7404
rect 6828 7284 6880 7336
rect 7564 7327 7616 7336
rect 7564 7293 7573 7327
rect 7573 7293 7607 7327
rect 7607 7293 7616 7327
rect 7564 7284 7616 7293
rect 9588 7284 9640 7336
rect 8484 7216 8536 7268
rect 5724 7148 5776 7200
rect 10968 7148 11020 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 3424 6944 3476 6996
rect 9404 6944 9456 6996
rect 10324 6987 10376 6996
rect 10324 6953 10333 6987
rect 10333 6953 10367 6987
rect 10367 6953 10376 6987
rect 10324 6944 10376 6953
rect 10876 6876 10928 6928
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 5908 6740 5960 6792
rect 7564 6851 7616 6860
rect 7564 6817 7573 6851
rect 7573 6817 7607 6851
rect 7607 6817 7616 6851
rect 7564 6808 7616 6817
rect 8208 6808 8260 6860
rect 9772 6808 9824 6860
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 11980 6808 12032 6860
rect 19892 6740 19944 6792
rect 21548 6672 21600 6724
rect 6920 6604 6972 6656
rect 7012 6647 7064 6656
rect 7012 6613 7021 6647
rect 7021 6613 7055 6647
rect 7055 6613 7064 6647
rect 7380 6647 7432 6656
rect 7012 6604 7064 6613
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 7472 6647 7524 6656
rect 7472 6613 7481 6647
rect 7481 6613 7515 6647
rect 7515 6613 7524 6647
rect 7472 6604 7524 6613
rect 8208 6604 8260 6656
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 10140 6604 10192 6656
rect 10876 6604 10928 6656
rect 10968 6604 11020 6656
rect 18972 6604 19024 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 4068 6400 4120 6452
rect 5632 6400 5684 6452
rect 7748 6400 7800 6452
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 10140 6443 10192 6452
rect 10140 6409 10149 6443
rect 10149 6409 10183 6443
rect 10183 6409 10192 6443
rect 10140 6400 10192 6409
rect 10968 6400 11020 6452
rect 6920 6332 6972 6384
rect 21456 6400 21508 6452
rect 7564 6264 7616 6316
rect 8484 6264 8536 6316
rect 4068 6196 4120 6248
rect 5908 6239 5960 6248
rect 5908 6205 5917 6239
rect 5917 6205 5951 6239
rect 5951 6205 5960 6239
rect 5908 6196 5960 6205
rect 5632 6128 5684 6180
rect 6828 6196 6880 6248
rect 9312 6196 9364 6248
rect 9772 6239 9824 6248
rect 9772 6205 9781 6239
rect 9781 6205 9815 6239
rect 9815 6205 9824 6239
rect 9772 6196 9824 6205
rect 4160 6060 4212 6112
rect 7380 6128 7432 6180
rect 7196 6103 7248 6112
rect 7196 6069 7205 6103
rect 7205 6069 7239 6103
rect 7239 6069 7248 6103
rect 7196 6060 7248 6069
rect 7472 6060 7524 6112
rect 9496 6060 9548 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 7380 5856 7432 5908
rect 8208 5856 8260 5908
rect 9312 5899 9364 5908
rect 9312 5865 9321 5899
rect 9321 5865 9355 5899
rect 9355 5865 9364 5899
rect 9312 5856 9364 5865
rect 8484 5831 8536 5840
rect 8484 5797 8493 5831
rect 8493 5797 8527 5831
rect 8527 5797 8536 5831
rect 8484 5788 8536 5797
rect 4068 5584 4120 5636
rect 10876 5584 10928 5636
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 4068 5312 4120 5364
rect 7656 5312 7708 5364
rect 3976 5244 4028 5296
rect 7196 5244 7248 5296
rect 10876 5219 10928 5228
rect 10876 5185 10885 5219
rect 10885 5185 10919 5219
rect 10919 5185 10928 5219
rect 10876 5176 10928 5185
rect 21180 5040 21232 5092
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 4068 4088 4120 4140
rect 5724 4088 5776 4140
rect 3424 4020 3476 4072
rect 8300 4020 8352 4072
rect 3976 3952 4028 4004
rect 9956 3952 10008 4004
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 3516 2592 3568 2644
rect 11888 2592 11940 2644
rect 4068 2524 4120 2576
rect 5632 2524 5684 2576
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 2872 1776 2924 1828
rect 5540 1776 5592 1828
<< metal2 >>
rect 202 22200 258 23000
rect 400 22222 612 22250
rect 216 18630 244 22200
rect 204 18624 256 18630
rect 204 18566 256 18572
rect 400 11830 428 22222
rect 584 22114 612 22222
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2962 22200 3018 23000
rect 3422 22200 3478 23000
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 5920 22222 6132 22250
rect 676 22114 704 22200
rect 584 22086 704 22114
rect 1136 19174 1164 22200
rect 1490 20088 1546 20097
rect 1490 20023 1492 20032
rect 1544 20023 1546 20032
rect 1492 19994 1544 20000
rect 1400 19984 1452 19990
rect 1400 19926 1452 19932
rect 1124 19168 1176 19174
rect 1124 19110 1176 19116
rect 1412 14074 1440 19926
rect 1596 19446 1624 22200
rect 1950 21312 2006 21321
rect 1950 21247 2006 21256
rect 1964 19938 1992 21247
rect 2056 20584 2084 22200
rect 2056 20556 2176 20584
rect 2042 20496 2098 20505
rect 2042 20431 2098 20440
rect 2056 20058 2084 20431
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 1964 19910 2084 19938
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1688 19446 1716 19790
rect 1950 19680 2006 19689
rect 1950 19615 2006 19624
rect 1964 19514 1992 19615
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1584 19440 1636 19446
rect 1584 19382 1636 19388
rect 1676 19440 1728 19446
rect 1676 19382 1728 19388
rect 1950 18048 2006 18057
rect 1950 17983 2006 17992
rect 1964 17882 1992 17983
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 1950 17640 2006 17649
rect 1950 17575 2006 17584
rect 1766 17504 1822 17513
rect 1766 17439 1822 17448
rect 1674 16688 1730 16697
rect 1674 16623 1730 16632
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1412 13394 1440 14010
rect 1400 13388 1452 13394
rect 1400 13330 1452 13336
rect 388 11824 440 11830
rect 388 11766 440 11772
rect 1504 11218 1532 16050
rect 1582 13152 1638 13161
rect 1582 13087 1638 13096
rect 1596 12442 1624 13087
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1504 10470 1532 10610
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1504 7857 1532 10406
rect 1688 9382 1716 16623
rect 1780 10810 1808 17439
rect 1964 17338 1992 17575
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 1950 17232 2006 17241
rect 1950 17167 2006 17176
rect 1858 16824 1914 16833
rect 1964 16794 1992 17167
rect 1858 16759 1914 16768
rect 1952 16788 2004 16794
rect 1872 15706 1900 16759
rect 1952 16730 2004 16736
rect 2056 16250 2084 19910
rect 2148 18970 2176 20556
rect 2516 19990 2544 22200
rect 2778 20904 2834 20913
rect 2778 20839 2834 20848
rect 2792 20058 2820 20839
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2136 18964 2188 18970
rect 2136 18906 2188 18912
rect 2320 18896 2372 18902
rect 2318 18864 2320 18873
rect 2372 18864 2374 18873
rect 2318 18799 2374 18808
rect 2410 18456 2466 18465
rect 2410 18391 2466 18400
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 1950 16008 2006 16017
rect 1950 15943 2006 15952
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1964 14618 1992 15943
rect 2424 15706 2452 18391
rect 2516 18358 2544 19790
rect 2870 19272 2926 19281
rect 2870 19207 2926 19216
rect 2504 18352 2556 18358
rect 2504 18294 2556 18300
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2700 17270 2728 17614
rect 2792 17338 2820 18226
rect 2884 17882 2912 19207
rect 2976 18902 3004 22200
rect 3436 19530 3464 22200
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3896 19530 3924 22200
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 3436 19502 3556 19530
rect 3896 19502 4016 19530
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2964 18896 3016 18902
rect 2964 18838 3016 18844
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2688 17264 2740 17270
rect 2688 17206 2740 17212
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2884 16590 2912 17138
rect 3068 16794 3096 19246
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3160 16810 3188 18770
rect 3436 18358 3464 19314
rect 3528 19174 3556 19502
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 3238 18184 3294 18193
rect 3238 18119 3240 18128
rect 3292 18119 3294 18128
rect 3424 18148 3476 18154
rect 3240 18090 3292 18096
rect 3424 18090 3476 18096
rect 3252 17066 3280 18090
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 3056 16788 3108 16794
rect 2976 16748 3056 16776
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2792 16182 2820 16526
rect 2870 16416 2926 16425
rect 2870 16351 2926 16360
rect 2780 16176 2832 16182
rect 2780 16118 2832 16124
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2502 15600 2558 15609
rect 2502 15535 2558 15544
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 2148 15094 2176 15438
rect 2136 15088 2188 15094
rect 2136 15030 2188 15036
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2332 14822 2360 14962
rect 2320 14816 2372 14822
rect 2042 14784 2098 14793
rect 2320 14758 2372 14764
rect 2042 14719 2098 14728
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1860 13796 1912 13802
rect 1860 13738 1912 13744
rect 1872 13190 1900 13738
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12646 1900 13126
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 2056 10266 2084 14719
rect 2516 14618 2544 15535
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2134 13560 2190 13569
rect 2134 13495 2190 13504
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 2148 9178 2176 13495
rect 2240 12306 2268 14350
rect 2504 14340 2556 14346
rect 2504 14282 2556 14288
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2332 13530 2360 13806
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2424 13394 2452 13670
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2424 13258 2452 13330
rect 2412 13252 2464 13258
rect 2412 13194 2464 13200
rect 2424 12850 2452 13194
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2332 11694 2360 12786
rect 2410 12336 2466 12345
rect 2410 12271 2466 12280
rect 2424 12238 2452 12271
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2516 10606 2544 14282
rect 2608 12918 2636 14962
rect 2596 12912 2648 12918
rect 2596 12854 2648 12860
rect 2700 10742 2728 15438
rect 2884 15162 2912 16351
rect 2976 15706 3004 16748
rect 3160 16782 3280 16810
rect 3056 16730 3108 16736
rect 3148 16040 3200 16046
rect 3068 15988 3148 15994
rect 3068 15982 3200 15988
rect 3068 15966 3188 15982
rect 3068 15910 3096 15966
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2962 15192 3018 15201
rect 2872 15156 2924 15162
rect 2962 15127 3018 15136
rect 2872 15098 2924 15104
rect 2870 14376 2926 14385
rect 2870 14311 2926 14320
rect 2778 13968 2834 13977
rect 2778 13903 2834 13912
rect 2792 11354 2820 13903
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2884 10826 2912 14311
rect 2976 11898 3004 15127
rect 3068 13297 3096 15846
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3160 14346 3188 15642
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3160 13326 3188 14282
rect 3148 13320 3200 13326
rect 3054 13288 3110 13297
rect 3148 13262 3200 13268
rect 3054 13223 3110 13232
rect 3160 12986 3188 13262
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 3068 12238 3096 12718
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3160 12306 3188 12582
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3146 12200 3202 12209
rect 3146 12135 3202 12144
rect 3160 12102 3188 12135
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3160 11898 3188 12038
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3056 11552 3108 11558
rect 3160 11529 3188 11630
rect 3056 11494 3108 11500
rect 3146 11520 3202 11529
rect 2884 10798 3004 10826
rect 2688 10736 2740 10742
rect 2688 10678 2740 10684
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2884 10266 2912 10610
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2332 8974 2360 9454
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 1490 7848 1546 7857
rect 1490 7783 1546 7792
rect 2792 7449 2820 9522
rect 2976 9450 3004 10798
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 3068 8265 3096 11494
rect 3146 11455 3202 11464
rect 3252 11121 3280 16782
rect 3344 16250 3372 17070
rect 3436 16250 3464 18090
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3896 17882 3924 19314
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3620 17338 3648 17478
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3700 16720 3752 16726
rect 3700 16662 3752 16668
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3344 15473 3372 16050
rect 3436 15638 3464 16186
rect 3712 16182 3740 16662
rect 3700 16176 3752 16182
rect 3700 16118 3752 16124
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3424 15632 3476 15638
rect 3424 15574 3476 15580
rect 3330 15464 3386 15473
rect 3330 15399 3386 15408
rect 3424 15428 3476 15434
rect 3424 15370 3476 15376
rect 3436 15094 3464 15370
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 3988 15042 4016 19502
rect 4172 18970 4200 19926
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4172 18426 4200 18906
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 4080 16182 4108 17546
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4172 16794 4200 17138
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4080 15178 4108 15982
rect 4080 15150 4200 15178
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3344 14414 3372 14894
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3344 13802 3372 14214
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 3344 13394 3372 13738
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3238 11112 3294 11121
rect 3238 11047 3294 11056
rect 3344 9897 3372 12786
rect 3436 10713 3464 15030
rect 3884 15020 3936 15026
rect 3988 15014 4108 15042
rect 3884 14962 3936 14968
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 3528 14074 3556 14486
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3712 13870 3740 14350
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3896 13530 3924 14962
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3988 14618 4016 14894
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 4080 13802 4108 15014
rect 4172 14618 4200 15150
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4264 14550 4292 19110
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 4252 14340 4304 14346
rect 4252 14282 4304 14288
rect 4264 14074 4292 14282
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4080 13410 4108 13466
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3896 13382 4108 13410
rect 3528 12646 3556 13330
rect 3896 12753 3924 13382
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3988 12918 4016 13126
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 3882 12744 3938 12753
rect 3882 12679 3938 12688
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3804 11778 3832 12242
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3896 11937 3924 12106
rect 3882 11928 3938 11937
rect 3988 11898 4016 12854
rect 4172 12442 4200 13874
rect 4264 13394 4292 14010
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 3882 11863 3938 11872
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3804 11750 3924 11778
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3896 11121 3924 11750
rect 4080 11558 4108 12310
rect 4264 11642 4292 13126
rect 4172 11614 4292 11642
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4172 11286 4200 11614
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 4068 11144 4120 11150
rect 3514 11112 3570 11121
rect 3514 11047 3516 11056
rect 3568 11047 3570 11056
rect 3882 11112 3938 11121
rect 4068 11086 4120 11092
rect 3882 11047 3938 11056
rect 3516 11018 3568 11024
rect 4080 10742 4108 11086
rect 4068 10736 4120 10742
rect 3422 10704 3478 10713
rect 3422 10639 3478 10648
rect 3606 10704 3662 10713
rect 4068 10678 4120 10684
rect 4172 10674 4200 11222
rect 4264 11150 4292 11494
rect 4356 11150 4384 22200
rect 4528 19440 4580 19446
rect 4528 19382 4580 19388
rect 4540 19174 4568 19382
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4540 18902 4568 19110
rect 4528 18896 4580 18902
rect 4528 18838 4580 18844
rect 4436 18216 4488 18222
rect 4436 18158 4488 18164
rect 4448 17678 4476 18158
rect 4540 17882 4568 18838
rect 4712 18216 4764 18222
rect 4632 18164 4712 18170
rect 4632 18158 4764 18164
rect 4632 18142 4752 18158
rect 4816 18154 4844 22200
rect 5276 20602 5304 22200
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 5184 19514 5212 19994
rect 5276 19786 5304 20538
rect 5368 19854 5396 20538
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5460 19417 5488 19654
rect 5446 19408 5502 19417
rect 5446 19343 5502 19352
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 4804 18148 4856 18154
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 4540 17338 4568 17478
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4632 17218 4660 18142
rect 4804 18090 4856 18096
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4540 17190 4660 17218
rect 4434 15056 4490 15065
rect 4434 14991 4490 15000
rect 4448 14958 4476 14991
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4448 13462 4476 14486
rect 4540 13530 4568 17190
rect 4724 16794 4752 17818
rect 4908 17678 4936 18022
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4908 17270 4936 17614
rect 5000 17338 5028 18906
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 5092 17814 5120 18566
rect 5080 17808 5132 17814
rect 5080 17750 5132 17756
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 5092 16658 5120 17750
rect 5276 17746 5304 19110
rect 5552 18698 5580 20334
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5644 19242 5672 20198
rect 5632 19236 5684 19242
rect 5632 19178 5684 19184
rect 5540 18692 5592 18698
rect 5540 18634 5592 18640
rect 5644 18612 5672 19178
rect 5736 18970 5764 22200
rect 5816 20324 5868 20330
rect 5816 20266 5868 20272
rect 5828 19854 5856 20266
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5724 18624 5776 18630
rect 5644 18584 5724 18612
rect 5724 18566 5776 18572
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 5184 17270 5212 17478
rect 5172 17264 5224 17270
rect 5172 17206 5224 17212
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5184 16969 5212 17070
rect 5170 16960 5226 16969
rect 5170 16895 5226 16904
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 5184 16114 5212 16730
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5000 15502 5028 15846
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4620 14884 4672 14890
rect 4620 14826 4672 14832
rect 4632 14278 4660 14826
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5000 14550 5028 14758
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4816 13870 4844 14010
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4436 13456 4488 13462
rect 4436 13398 4488 13404
rect 4448 13274 4476 13398
rect 4632 13326 4660 13670
rect 4620 13320 4672 13326
rect 4448 13246 4568 13274
rect 4620 13262 4672 13268
rect 4540 13190 4568 13246
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4448 12238 4476 12718
rect 4632 12434 4660 13262
rect 4540 12406 4660 12434
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4540 11694 4568 12406
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4356 10810 4384 11086
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 3606 10639 3608 10648
rect 3660 10639 3662 10648
rect 4160 10668 4212 10674
rect 3608 10610 3660 10616
rect 4160 10610 4212 10616
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3422 10296 3478 10305
rect 3549 10299 3857 10308
rect 3422 10231 3478 10240
rect 3436 10198 3464 10231
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 3330 9888 3386 9897
rect 3330 9823 3386 9832
rect 3974 9480 4030 9489
rect 3974 9415 4030 9424
rect 4068 9444 4120 9450
rect 3988 9382 4016 9415
rect 4068 9386 4120 9392
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3976 9104 4028 9110
rect 4080 9081 4108 9386
rect 3976 9046 4028 9052
rect 4066 9072 4122 9081
rect 3988 8673 4016 9046
rect 4066 9007 4122 9016
rect 3974 8664 4030 8673
rect 3974 8599 4030 8608
rect 3054 8256 3110 8265
rect 3054 8191 3110 8200
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 2778 7440 2834 7449
rect 2778 7375 2834 7384
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3422 7032 3478 7041
rect 3549 7035 3857 7044
rect 3422 6967 3424 6976
rect 3476 6967 3478 6976
rect 3424 6938 3476 6944
rect 4066 6624 4122 6633
rect 4066 6559 4122 6568
rect 4080 6458 4108 6559
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4068 6248 4120 6254
rect 4066 6216 4068 6225
rect 4120 6216 4122 6225
rect 4066 6151 4122 6160
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 4080 5642 4108 5743
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 4066 5400 4122 5409
rect 4066 5335 4068 5344
rect 4120 5335 4122 5344
rect 4068 5306 4120 5312
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3988 4185 4016 5238
rect 4172 5137 4200 6054
rect 4158 5128 4214 5137
rect 4158 5063 4214 5072
rect 4448 4593 4476 11290
rect 4632 10810 4660 12242
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4540 9178 4568 9522
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4632 8022 4660 9862
rect 4724 8634 4752 13738
rect 4816 12306 4844 13806
rect 5092 13734 5120 15506
rect 5184 13977 5212 16050
rect 5276 16017 5304 17682
rect 5368 16250 5396 18362
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5460 17882 5488 18226
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5262 16008 5318 16017
rect 5262 15943 5318 15952
rect 5368 15434 5396 16186
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5446 15056 5502 15065
rect 5446 14991 5502 15000
rect 5460 14618 5488 14991
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5170 13968 5226 13977
rect 5170 13903 5226 13912
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 5184 13394 5212 13806
rect 5368 13394 5396 14350
rect 5552 14074 5580 17138
rect 5644 17134 5672 18022
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5736 15502 5764 18566
rect 5828 17241 5856 19790
rect 5920 18426 5948 22222
rect 6104 22114 6132 22222
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20088 22222 20392 22250
rect 6196 22114 6224 22200
rect 6104 22086 6224 22114
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6012 19514 6040 20402
rect 6184 20392 6236 20398
rect 6184 20334 6236 20340
rect 6196 19718 6224 20334
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6552 19712 6604 19718
rect 6552 19654 6604 19660
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 6564 19514 6592 19654
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6288 18630 6316 18770
rect 6276 18624 6328 18630
rect 6276 18566 6328 18572
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 6104 17785 6132 18022
rect 6090 17776 6146 17785
rect 6090 17711 6092 17720
rect 6144 17711 6146 17720
rect 6092 17682 6144 17688
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5920 17338 5948 17478
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5814 17232 5870 17241
rect 5814 17167 5870 17176
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 13433 5488 13738
rect 5446 13424 5502 13433
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5356 13388 5408 13394
rect 5446 13359 5502 13368
rect 5356 13330 5408 13336
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5276 12986 5304 13194
rect 5368 12986 5396 13330
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5170 12880 5226 12889
rect 5170 12815 5226 12824
rect 5184 12782 5212 12815
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5644 12442 5672 14962
rect 5736 14906 5764 15302
rect 5828 15162 5856 16526
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 5736 14878 5856 14906
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 4986 12336 5042 12345
rect 4804 12300 4856 12306
rect 4986 12271 4988 12280
rect 4804 12242 4856 12248
rect 5040 12271 5042 12280
rect 4988 12242 5040 12248
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 5092 11898 5120 12038
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5460 11354 5488 11630
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5184 11150 5212 11290
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 5000 10062 5028 11018
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5184 9518 5212 11086
rect 5538 10568 5594 10577
rect 5538 10503 5594 10512
rect 5552 10130 5580 10503
rect 5644 10266 5672 11154
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5736 10198 5764 14758
rect 5828 14618 5856 14878
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5920 12434 5948 17070
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6012 16250 6040 16662
rect 6564 16590 6592 19314
rect 6656 16794 6684 22200
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 6736 20324 6788 20330
rect 6736 20266 6788 20272
rect 6748 19854 6776 20266
rect 6828 20256 6880 20262
rect 6826 20224 6828 20233
rect 6880 20224 6882 20233
rect 6826 20159 6882 20168
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6656 16046 6684 16730
rect 6748 16425 6776 19790
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6840 18698 6868 19722
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6840 17338 6868 18362
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6932 17134 6960 18022
rect 7024 17270 7052 20402
rect 7116 17882 7144 22200
rect 7576 19802 7604 22200
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7576 19774 7788 19802
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7484 19514 7512 19654
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7576 19446 7604 19654
rect 7564 19440 7616 19446
rect 7286 19408 7342 19417
rect 7564 19382 7616 19388
rect 7286 19343 7342 19352
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 7116 16726 7144 17818
rect 7300 17728 7328 19343
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7392 18358 7420 18566
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 7300 17700 7420 17728
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7104 16720 7156 16726
rect 7104 16662 7156 16668
rect 7194 16688 7250 16697
rect 7194 16623 7196 16632
rect 7248 16623 7250 16632
rect 7196 16594 7248 16600
rect 6920 16448 6972 16454
rect 6734 16416 6790 16425
rect 6920 16390 6972 16396
rect 6734 16351 6790 16360
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6000 15972 6052 15978
rect 6000 15914 6052 15920
rect 6012 13530 6040 15914
rect 6288 15570 6316 15982
rect 6748 15706 6776 16351
rect 6932 16250 6960 16390
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6276 15564 6328 15570
rect 6748 15552 6776 15642
rect 6276 15506 6328 15512
rect 6656 15524 6776 15552
rect 6288 15366 6316 15506
rect 6656 15434 6684 15524
rect 6644 15428 6696 15434
rect 6644 15370 6696 15376
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6550 15328 6606 15337
rect 6148 15260 6456 15269
rect 6550 15263 6606 15272
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6104 14793 6132 14894
rect 6090 14784 6146 14793
rect 6090 14719 6146 14728
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6564 13462 6592 15263
rect 6644 14884 6696 14890
rect 6644 14826 6696 14832
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 5920 12406 6040 12434
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5828 9926 5856 10950
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5828 9450 5856 9862
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5920 9382 5948 11494
rect 6012 10169 6040 12406
rect 6288 12306 6316 12786
rect 6460 12776 6512 12782
rect 6564 12764 6592 13262
rect 6656 12918 6684 14826
rect 6748 14822 6776 15370
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6840 14278 6868 16118
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6840 13274 6868 14214
rect 6932 13734 6960 15302
rect 7116 15094 7144 15574
rect 7104 15088 7156 15094
rect 7104 15030 7156 15036
rect 7012 14952 7064 14958
rect 7010 14920 7012 14929
rect 7064 14920 7066 14929
rect 7010 14855 7066 14864
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7024 14074 7052 14214
rect 7116 14074 7144 14758
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7010 13968 7066 13977
rect 7010 13903 7066 13912
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6840 13246 6960 13274
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6512 12736 6592 12764
rect 6644 12776 6696 12782
rect 6460 12718 6512 12724
rect 6644 12718 6696 12724
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6656 12170 6684 12718
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6656 11898 6684 12106
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6642 11656 6698 11665
rect 6642 11591 6698 11600
rect 6182 11248 6238 11257
rect 6182 11183 6184 11192
rect 6236 11183 6238 11192
rect 6184 11154 6236 11160
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6564 10198 6592 10542
rect 6552 10192 6604 10198
rect 5998 10160 6054 10169
rect 6552 10134 6604 10140
rect 6656 10146 6684 11591
rect 6748 11558 6776 12038
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6748 10810 6776 11154
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6734 10704 6790 10713
rect 6734 10639 6790 10648
rect 6748 10538 6776 10639
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6840 10266 6868 13126
rect 6932 11665 6960 13246
rect 7024 12170 7052 13903
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 7116 13297 7144 13738
rect 7208 13462 7236 15914
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 7102 13288 7158 13297
rect 7102 13223 7158 13232
rect 7300 12986 7328 17546
rect 7392 15994 7420 17700
rect 7576 17134 7604 19246
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7668 17338 7696 18226
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7654 16416 7710 16425
rect 7392 15966 7512 15994
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7392 15706 7420 15846
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7392 12866 7420 15370
rect 7484 14657 7512 15966
rect 7576 15366 7604 16390
rect 7654 16351 7710 16360
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7470 14648 7526 14657
rect 7470 14583 7526 14592
rect 7576 14414 7604 14962
rect 7668 14618 7696 16351
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7668 14226 7696 14418
rect 7208 12838 7420 12866
rect 7576 14198 7696 14226
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 7208 11898 7236 12838
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 6918 11656 6974 11665
rect 6918 11591 6974 11600
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6656 10118 6868 10146
rect 5998 10095 6054 10104
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 6012 9722 6040 9930
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5170 9072 5226 9081
rect 5170 9007 5172 9016
rect 5224 9007 5226 9016
rect 5632 9036 5684 9042
rect 5172 8978 5224 8984
rect 5632 8978 5684 8984
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 5644 8566 5672 8978
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 5552 7750 5580 8366
rect 6012 8090 6040 8910
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6380 7954 6408 8230
rect 6656 7954 6684 8978
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 4434 4584 4490 4593
rect 4434 4519 4490 4528
rect 3974 4176 4030 4185
rect 3974 4111 4030 4120
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3436 3777 3464 4014
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3422 3768 3478 3777
rect 3549 3771 3857 3780
rect 3422 3703 3478 3712
rect 3988 2961 4016 3946
rect 4080 3369 4108 4082
rect 4066 3360 4122 3369
rect 4066 3295 4122 3304
rect 3974 2952 4030 2961
rect 3974 2887 4030 2896
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3528 2145 3556 2586
rect 4068 2576 4120 2582
rect 4066 2544 4068 2553
rect 4120 2544 4122 2553
rect 4066 2479 4122 2488
rect 3514 2136 3570 2145
rect 3514 2071 3570 2080
rect 5552 1834 5580 7686
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6656 7546 6684 7890
rect 6748 7886 6776 8434
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5736 7206 5764 7346
rect 6840 7342 6868 10118
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9518 6960 9862
rect 6920 9512 6972 9518
rect 7024 9500 7052 10678
rect 7300 10470 7328 11766
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7484 10266 7512 11086
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7116 9654 7144 9930
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7104 9512 7156 9518
rect 7024 9472 7104 9500
rect 6920 9454 6972 9460
rect 7104 9454 7156 9460
rect 6932 9178 6960 9454
rect 7116 9194 7144 9454
rect 7208 9382 7236 10134
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 6920 9172 6972 9178
rect 7116 9166 7236 9194
rect 6920 9114 6972 9120
rect 7208 8838 7236 9166
rect 7300 8906 7328 9454
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5644 6458 5672 6734
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5644 2582 5672 6122
rect 5736 4146 5764 7142
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 6254 5948 6734
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6840 6254 6868 7278
rect 6932 7018 6960 8774
rect 7208 8514 7236 8774
rect 7392 8634 7420 9522
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7208 8486 7420 8514
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7024 7546 7052 7686
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7116 7478 7144 8366
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 6932 6990 7052 7018
rect 7024 6662 7052 6990
rect 7392 6662 7420 8486
rect 7576 7426 7604 14198
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7668 12102 7696 13126
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7484 7398 7604 7426
rect 7484 6662 7512 7398
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7576 6866 7604 7278
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 6932 6390 6960 6598
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 7392 6186 7420 6598
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 7208 5302 7236 6054
rect 7392 5914 7420 6122
rect 7484 6118 7512 6598
rect 7576 6322 7604 6802
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7668 5370 7696 12038
rect 7760 7954 7788 19774
rect 7944 19310 7972 20198
rect 7932 19304 7984 19310
rect 7932 19246 7984 19252
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7852 18426 7880 19110
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7944 18306 7972 19110
rect 7852 18278 7972 18306
rect 7852 18222 7880 18278
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 7852 14521 7880 18158
rect 8036 17921 8064 22200
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8116 18692 8168 18698
rect 8116 18634 8168 18640
rect 8022 17912 8078 17921
rect 8022 17847 8078 17856
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 7944 17338 7972 17478
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 8036 16810 8064 17478
rect 7944 16782 8064 16810
rect 7944 16250 7972 16782
rect 8022 16688 8078 16697
rect 8022 16623 8024 16632
rect 8076 16623 8078 16632
rect 8024 16594 8076 16600
rect 8128 16590 8156 18634
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8220 18426 8248 18566
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8220 16454 8248 17002
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 8022 15600 8078 15609
rect 8022 15535 8024 15544
rect 8076 15535 8078 15544
rect 8024 15506 8076 15512
rect 8220 15502 8248 16390
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 7932 15360 7984 15366
rect 8116 15360 8168 15366
rect 7984 15320 8064 15348
rect 7932 15302 7984 15308
rect 7930 15192 7986 15201
rect 8036 15162 8064 15320
rect 8116 15302 8168 15308
rect 7930 15127 7986 15136
rect 8024 15156 8076 15162
rect 7838 14512 7894 14521
rect 7838 14447 7894 14456
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7852 13530 7880 13806
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 7852 12646 7880 12854
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7838 11792 7894 11801
rect 7838 11727 7840 11736
rect 7892 11727 7894 11736
rect 7840 11698 7892 11704
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9761 7880 9862
rect 7838 9752 7894 9761
rect 7838 9687 7840 9696
rect 7892 9687 7894 9696
rect 7840 9658 7892 9664
rect 7944 8430 7972 15127
rect 8024 15098 8076 15104
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 8036 14482 8064 14962
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 8128 14074 8156 15302
rect 8208 14884 8260 14890
rect 8208 14826 8260 14832
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8220 13682 8248 14826
rect 8312 14482 8340 20402
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8404 15337 8432 16594
rect 8496 15502 8524 22200
rect 8956 20346 8984 22200
rect 9416 20346 9444 22200
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 8956 20318 9168 20346
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8588 18154 8616 19314
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8680 17762 8708 18022
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 8680 17734 8800 17762
rect 8772 17678 8800 17734
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8588 17202 8616 17478
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8390 15328 8446 15337
rect 8390 15263 8446 15272
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 8404 14793 8432 15098
rect 8496 15094 8524 15438
rect 8484 15088 8536 15094
rect 8484 15030 8536 15036
rect 8390 14784 8446 14793
rect 8390 14719 8446 14728
rect 8482 14648 8538 14657
rect 8392 14612 8444 14618
rect 8482 14583 8538 14592
rect 8392 14554 8444 14560
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8404 13938 8432 14554
rect 8496 14414 8524 14583
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8588 14074 8616 16186
rect 8680 16153 8708 17614
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8864 17270 8892 17546
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8956 17338 8984 17478
rect 9048 17338 9076 17682
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 8852 17264 8904 17270
rect 8852 17206 8904 17212
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 9034 16416 9090 16425
rect 9034 16351 9090 16360
rect 8666 16144 8722 16153
rect 9048 16114 9076 16351
rect 8666 16079 8722 16088
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 8668 15632 8720 15638
rect 8666 15600 8668 15609
rect 8720 15600 8722 15609
rect 8666 15535 8722 15544
rect 8850 15464 8906 15473
rect 8850 15399 8906 15408
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8128 13654 8248 13682
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 8036 12306 8064 12786
rect 8128 12434 8156 13654
rect 8404 13394 8432 13670
rect 8588 13530 8616 14010
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8208 12776 8260 12782
rect 8206 12744 8208 12753
rect 8260 12744 8262 12753
rect 8206 12679 8262 12688
rect 8128 12406 8248 12434
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8022 12200 8078 12209
rect 8022 12135 8078 12144
rect 8036 10606 8064 12135
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8128 11354 8156 12038
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 8220 10418 8248 12406
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8036 10390 8248 10418
rect 8036 9654 8064 10390
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 8220 9602 8248 10202
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8312 9722 8340 9862
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8220 9574 8340 9602
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8036 8974 8064 9114
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 8036 8294 8064 8910
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8220 8430 8248 8842
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8128 8022 8156 8366
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7760 6458 7788 7890
rect 8128 7546 8156 7958
rect 8220 7954 8248 8366
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8220 6866 8248 7890
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 8220 5914 8248 6598
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 8312 4078 8340 9574
rect 8404 9450 8432 10610
rect 8496 10130 8524 10678
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8588 10010 8616 12786
rect 8680 11354 8708 15302
rect 8864 14890 8892 15399
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9140 14482 9168 20318
rect 9232 20318 9444 20346
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 9140 11150 9168 14010
rect 9232 12986 9260 20318
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9324 19281 9352 20198
rect 9404 19984 9456 19990
rect 9402 19952 9404 19961
rect 9456 19952 9458 19961
rect 9402 19887 9458 19896
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9310 19272 9366 19281
rect 9310 19207 9366 19216
rect 9416 19156 9444 19790
rect 9324 19128 9444 19156
rect 9324 17746 9352 19128
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9312 17740 9364 17746
rect 9312 17682 9364 17688
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9324 16250 9352 17138
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9310 16144 9366 16153
rect 9310 16079 9366 16088
rect 9324 15042 9352 16079
rect 9416 15706 9444 18226
rect 9508 17270 9536 20402
rect 9876 19990 9904 22200
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 9864 19984 9916 19990
rect 9864 19926 9916 19932
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9508 15201 9536 15642
rect 9600 15502 9628 19314
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9692 16590 9720 18634
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9494 15192 9550 15201
rect 9494 15127 9550 15136
rect 9324 15014 9444 15042
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9324 14618 9352 14894
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9324 14074 9352 14350
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9416 13716 9444 15014
rect 9692 13938 9720 16118
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9324 13688 9444 13716
rect 9324 13530 9352 13688
rect 9402 13560 9458 13569
rect 9312 13524 9364 13530
rect 9402 13495 9458 13504
rect 9312 13466 9364 13472
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9220 12844 9272 12850
rect 9324 12832 9352 13466
rect 9272 12804 9352 12832
rect 9220 12786 9272 12792
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9140 10470 9168 10950
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 8496 9982 8616 10010
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8404 7546 8432 8434
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8496 7274 8524 9982
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8588 8634 8616 9862
rect 9034 9616 9090 9625
rect 9034 9551 9090 9560
rect 9048 9518 9076 9551
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 9140 9110 9168 10406
rect 9232 9994 9260 12378
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9324 11898 9352 12038
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9324 10062 9352 10542
rect 9416 10130 9444 13495
rect 9508 11218 9536 13738
rect 9678 13696 9734 13705
rect 9678 13631 9734 13640
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9508 10266 9536 11018
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9508 9926 9536 10202
rect 9600 10130 9628 12718
rect 9692 10266 9720 13631
rect 9784 12442 9812 18702
rect 9876 16182 9904 19790
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9862 15464 9918 15473
rect 9862 15399 9918 15408
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9600 9178 9628 9522
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9692 9178 9720 9386
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9416 8634 9444 8774
rect 9784 8634 9812 10746
rect 9876 9042 9904 15399
rect 9968 15094 9996 19314
rect 10060 18766 10088 20334
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10152 18358 10180 20402
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 10244 18766 10272 19246
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 10336 17354 10364 22200
rect 10416 19984 10468 19990
rect 10416 19926 10468 19932
rect 10152 17326 10364 17354
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 10060 14074 10088 16526
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9968 12782 9996 13330
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9968 11830 9996 12038
rect 10060 11830 10088 13874
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 10048 11688 10100 11694
rect 10046 11656 10048 11665
rect 10100 11656 10102 11665
rect 10046 11591 10102 11600
rect 10060 11150 10088 11591
rect 10152 11218 10180 17326
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10244 16114 10272 16390
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10244 13394 10272 13874
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10336 12238 10364 13806
rect 10428 13530 10456 19926
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10598 18728 10654 18737
rect 10598 18663 10654 18672
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10520 16114 10548 18022
rect 10612 17270 10640 18663
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 15502 10548 15846
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10612 13258 10640 17070
rect 10704 16182 10732 19790
rect 10796 18408 10824 22200
rect 11256 19938 11284 22200
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11072 19910 11284 19938
rect 10796 18380 10916 18408
rect 10784 18284 10836 18290
rect 10784 18226 10836 18232
rect 10796 17678 10824 18226
rect 10888 18086 10916 18380
rect 10966 18320 11022 18329
rect 10966 18255 11022 18264
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10796 16028 10824 17002
rect 10888 16590 10916 17070
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10704 16000 10824 16028
rect 10704 14906 10732 16000
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10796 15026 10824 15302
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10704 14878 10824 14906
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10704 14482 10732 14758
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10796 14362 10824 14878
rect 10888 14618 10916 15302
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10704 14334 10824 14362
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10612 12986 10640 13194
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10704 12374 10732 14334
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10796 12714 10824 14214
rect 10888 14074 10916 14214
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10980 14006 11008 18255
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10888 11898 10916 13126
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10244 10810 10272 10950
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 10198 9996 10406
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 10060 9518 10088 9930
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8680 8090 8708 8502
rect 10060 8430 10088 9454
rect 10336 9081 10364 10950
rect 10980 10010 11008 13194
rect 10704 9982 11008 10010
rect 10704 9518 10732 9982
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10796 9722 10824 9862
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10796 9586 10824 9658
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10322 9072 10378 9081
rect 10322 9007 10378 9016
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 8496 6322 8524 7210
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9140 6458 9168 7346
rect 9416 7002 9444 7686
rect 9600 7546 9628 7890
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9600 7342 9628 7482
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8496 5846 8524 6258
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 9324 5914 9352 6190
rect 9508 6118 9536 6598
rect 9784 6254 9812 6802
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 9968 4010 9996 8298
rect 10060 8090 10088 8366
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10152 7886 10180 8434
rect 10704 8362 10732 9454
rect 10796 8974 10824 9522
rect 10888 9382 10916 9862
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10888 8430 10916 9318
rect 10980 9178 11008 9454
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 11072 9024 11100 19910
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11256 17746 11284 19790
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11244 17604 11296 17610
rect 11244 17546 11296 17552
rect 11164 13705 11192 17546
rect 11256 15042 11284 17546
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11716 17270 11744 22200
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11808 18358 11836 18566
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11704 17264 11756 17270
rect 11704 17206 11756 17212
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11348 15366 11376 15982
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11256 15014 11376 15042
rect 11716 15026 11744 16934
rect 11348 14498 11376 15014
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11532 14618 11560 14962
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11256 14470 11376 14498
rect 11150 13696 11206 13705
rect 11150 13631 11206 13640
rect 11150 13152 11206 13161
rect 11150 13087 11206 13096
rect 11164 12986 11192 13087
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11256 12345 11284 14470
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11242 12336 11298 12345
rect 11242 12271 11298 12280
rect 11532 12152 11560 12582
rect 11808 12442 11836 18022
rect 11888 17536 11940 17542
rect 11886 17504 11888 17513
rect 11940 17504 11942 17513
rect 11886 17439 11942 17448
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 16250 11928 16390
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11992 15094 12020 19858
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12084 17610 12112 18566
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 12176 16538 12204 22200
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12544 18970 12572 20538
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12452 18873 12480 18906
rect 12438 18864 12494 18873
rect 12438 18799 12494 18808
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12544 18698 12572 18770
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12438 18592 12494 18601
rect 12438 18527 12494 18536
rect 12452 18426 12480 18527
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12544 17882 12572 18362
rect 12636 18057 12664 22200
rect 13096 20534 13124 22200
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 13556 20262 13584 22200
rect 14016 20618 14044 22200
rect 13832 20590 14044 20618
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12728 19378 12756 19858
rect 12808 19848 12860 19854
rect 13832 19802 13860 20590
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 12808 19790 12860 19796
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12820 19174 12848 19790
rect 13648 19774 13860 19802
rect 13648 19514 13676 19774
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13740 19514 13768 19654
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 13004 19258 13032 19314
rect 12912 19230 13032 19258
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12728 18358 12756 18566
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12622 18048 12678 18057
rect 12622 17983 12678 17992
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12084 16510 12204 16538
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 11978 13288 12034 13297
rect 11978 13223 12034 13232
rect 11992 12986 12020 13223
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11992 12442 12020 12718
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11808 12306 11836 12378
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11164 12124 11560 12152
rect 11164 12073 11192 12124
rect 11704 12096 11756 12102
rect 11150 12064 11206 12073
rect 11704 12038 11756 12044
rect 11150 11999 11206 12008
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 10980 8996 11192 9024
rect 10980 8634 11008 8996
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10336 8022 10364 8230
rect 11072 8090 11100 8774
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11164 8022 11192 8996
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11716 8634 11744 12038
rect 12084 11642 12112 16510
rect 12268 13870 12296 17818
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12176 12646 12204 13262
rect 12268 13258 12296 13670
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12268 12782 12296 13194
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12360 12434 12388 17206
rect 12452 16454 12480 17750
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12530 17232 12586 17241
rect 12530 17167 12586 17176
rect 12544 16697 12572 17167
rect 12530 16688 12586 16697
rect 12530 16623 12586 16632
rect 12636 16522 12664 17478
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12268 12406 12388 12434
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12176 11801 12204 12038
rect 12162 11792 12218 11801
rect 12162 11727 12218 11736
rect 11992 11614 12112 11642
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11716 8498 11744 8570
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11716 8022 11744 8434
rect 10324 8016 10376 8022
rect 10324 7958 10376 7964
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11888 8016 11940 8022
rect 11888 7958 11940 7964
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10152 6662 10180 7822
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 10336 7002 10364 7414
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10888 6662 10916 6870
rect 10980 6866 11008 7142
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 6662 11008 6802
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10152 6458 10180 6598
rect 10980 6458 11008 6598
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10888 5234 10916 5578
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 11900 2650 11928 7958
rect 11992 6866 12020 11614
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12084 10606 12112 11494
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12084 8362 12112 8774
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12176 2774 12204 11727
rect 12268 8566 12296 12406
rect 12452 12238 12480 12922
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12360 11286 12388 11630
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12360 10062 12388 11222
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12452 8634 12480 9590
rect 12544 9042 12572 13942
rect 12636 13705 12664 16458
rect 12622 13696 12678 13705
rect 12622 13631 12678 13640
rect 12728 12170 12756 18294
rect 12820 14822 12848 19110
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12912 12889 12940 19230
rect 13740 18766 13768 19450
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 13452 18692 13504 18698
rect 13452 18634 13504 18640
rect 13280 17542 13308 18634
rect 13464 18290 13492 18634
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13372 17105 13400 17138
rect 13358 17096 13414 17105
rect 13358 17031 13414 17040
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13280 15910 13308 16458
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12898 12880 12954 12889
rect 12898 12815 12954 12824
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12912 12209 12940 12582
rect 12898 12200 12954 12209
rect 12716 12164 12768 12170
rect 12898 12135 12954 12144
rect 12716 12106 12768 12112
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12728 11218 12756 11698
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 13004 10810 13032 14894
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 12238 13124 13126
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 13188 11150 13216 13466
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13004 9654 13032 10746
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 13280 9178 13308 15846
rect 13464 15638 13492 18226
rect 13740 18086 13768 18702
rect 14188 18624 14240 18630
rect 14186 18592 14188 18601
rect 14240 18592 14242 18601
rect 14186 18527 14242 18536
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13740 17678 13768 18022
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13740 17134 13768 17614
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13740 16998 13768 17070
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 16794 13768 16934
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13832 16674 13860 18022
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 14186 17504 14242 17513
rect 14186 17439 14242 17448
rect 14200 16980 14228 17439
rect 14292 17202 14320 19450
rect 14476 18698 14504 22200
rect 14936 20330 14964 22200
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14464 18692 14516 18698
rect 14464 18634 14516 18640
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14476 17270 14504 17682
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14464 17264 14516 17270
rect 14464 17206 14516 17212
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14200 16952 14320 16980
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13556 16646 13860 16674
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 13556 15502 13584 16646
rect 13820 16584 13872 16590
rect 13634 16552 13690 16561
rect 13820 16526 13872 16532
rect 13634 16487 13690 16496
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13556 14074 13584 14350
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13372 11762 13400 13126
rect 13464 12986 13492 13874
rect 13648 13258 13676 16487
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13740 16250 13768 16390
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13740 15706 13768 16186
rect 13832 16182 13860 16526
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13832 15502 13860 16118
rect 14016 16114 14044 16730
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13832 15178 13860 15438
rect 14108 15366 14136 15642
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 13740 15150 13860 15178
rect 13740 15094 13768 15150
rect 14292 15094 14320 16952
rect 14384 16522 14412 17002
rect 14372 16516 14424 16522
rect 14372 16458 14424 16464
rect 14464 16516 14516 16522
rect 14464 16458 14516 16464
rect 14476 15434 14504 16458
rect 14464 15428 14516 15434
rect 14464 15370 14516 15376
rect 14476 15162 14504 15370
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 13740 14414 13768 15030
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13820 14544 13872 14550
rect 14292 14521 14320 14758
rect 13820 14486 13872 14492
rect 14278 14512 14334 14521
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 14278 13768 14350
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13740 13870 13768 14214
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13740 13326 13768 13806
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13740 12646 13768 13262
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13740 12238 13768 12582
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13464 11354 13492 12106
rect 13740 11830 13768 12174
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13740 11218 13768 11766
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13832 10674 13860 14486
rect 14278 14447 14334 14456
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13924 12850 13952 13466
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 14292 11257 14320 14447
rect 14476 13938 14504 14826
rect 14568 14346 14596 17478
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14476 12918 14504 13194
rect 14568 13161 14596 14282
rect 14554 13152 14610 13161
rect 14554 13087 14610 13096
rect 14464 12912 14516 12918
rect 14464 12854 14516 12860
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14476 12102 14504 12242
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14278 11248 14334 11257
rect 14278 11183 14334 11192
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 14292 10674 14320 11018
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 13832 10198 13860 10610
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 14384 10266 14412 11086
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13924 9722 13952 9998
rect 14096 9920 14148 9926
rect 14568 9908 14596 12786
rect 14660 12306 14688 19654
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 15212 18426 15240 19314
rect 15304 18698 15332 19790
rect 15396 19786 15424 22200
rect 15856 19990 15884 22200
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 16316 19922 16344 22200
rect 16776 20890 16804 22200
rect 16776 20862 16988 20890
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16764 19440 16816 19446
rect 16816 19400 16896 19428
rect 16764 19382 16816 19388
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15568 18896 15620 18902
rect 15382 18864 15438 18873
rect 15568 18838 15620 18844
rect 15382 18799 15438 18808
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 15396 18426 15424 18799
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 14740 17604 14792 17610
rect 14740 17546 14792 17552
rect 14752 14822 14780 17546
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 14936 15026 14964 15846
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14752 13530 14780 14758
rect 14936 14634 14964 14962
rect 14844 14606 14964 14634
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14752 12209 14780 12854
rect 14738 12200 14794 12209
rect 14738 12135 14794 12144
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14752 10742 14780 11494
rect 14844 11354 14872 14606
rect 15120 14521 15148 15846
rect 15106 14512 15162 14521
rect 15106 14447 15162 14456
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14148 9880 14596 9908
rect 14096 9862 14148 9868
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12544 7886 12572 8978
rect 13280 8430 13308 9114
rect 14936 9110 14964 14010
rect 15028 14006 15056 14350
rect 15016 14000 15068 14006
rect 15016 13942 15068 13948
rect 15120 13852 15148 14447
rect 15028 13824 15148 13852
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 15028 8294 15056 13824
rect 15304 13530 15332 17478
rect 15488 16726 15516 18226
rect 15580 18086 15608 18838
rect 15764 18766 15792 19246
rect 16592 18986 16620 19314
rect 16500 18958 16620 18986
rect 16500 18902 16528 18958
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15764 18086 15792 18702
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16132 18086 16160 18634
rect 16868 18612 16896 19400
rect 16960 19174 16988 20862
rect 17236 19961 17264 22200
rect 17222 19952 17278 19961
rect 17222 19887 17278 19896
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16868 18584 16988 18612
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16960 18154 16988 18584
rect 17512 18290 17540 19450
rect 17696 18358 17724 22200
rect 18156 19281 18184 22200
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18236 19304 18288 19310
rect 18142 19272 18198 19281
rect 17960 19236 18012 19242
rect 18236 19246 18288 19252
rect 18142 19207 18198 19216
rect 17960 19178 18012 19184
rect 17684 18352 17736 18358
rect 17684 18294 17736 18300
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 16948 18148 17000 18154
rect 16948 18090 17000 18096
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 15764 17542 15792 18022
rect 15844 17604 15896 17610
rect 15844 17546 15896 17552
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15764 17066 15792 17478
rect 15752 17060 15804 17066
rect 15752 17002 15804 17008
rect 15476 16720 15528 16726
rect 15476 16662 15528 16668
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15106 13288 15162 13297
rect 15106 13223 15162 13232
rect 15120 11762 15148 13223
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15212 9994 15240 11290
rect 15304 10470 15332 12106
rect 15396 10810 15424 15914
rect 15488 13734 15516 16662
rect 15856 15706 15884 17546
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 16132 15366 16160 18022
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 17144 16454 17172 17682
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 17338 17448 17478
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16488 16176 16540 16182
rect 16488 16118 16540 16124
rect 16500 15978 16528 16118
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16408 15094 16436 15302
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 15842 14920 15898 14929
rect 15842 14855 15898 14864
rect 15856 14618 15884 14855
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15474 12744 15530 12753
rect 15474 12679 15530 12688
rect 15488 11354 15516 12679
rect 16408 12442 16436 15030
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16592 14550 16620 14894
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16592 14278 16620 14486
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16960 12850 16988 15846
rect 17040 15428 17092 15434
rect 17040 15370 17092 15376
rect 17052 14074 17080 15370
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15764 11286 15792 11766
rect 16132 11694 16160 12174
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16132 11558 16160 11630
rect 16316 11558 16344 11698
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 16132 11150 16160 11494
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 16132 10606 16160 11086
rect 17052 11082 17080 13466
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 17144 10724 17172 16390
rect 17236 11830 17264 17206
rect 17788 16794 17816 18226
rect 17972 17649 18000 19178
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 17958 17640 18014 17649
rect 17958 17575 18014 17584
rect 18064 17542 18092 18158
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 18248 17241 18276 19246
rect 18340 19174 18368 19654
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18340 18766 18368 19110
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18432 18329 18460 18566
rect 18418 18320 18474 18329
rect 18418 18255 18474 18264
rect 18524 18193 18552 19790
rect 18616 18970 18644 22200
rect 19076 20346 19104 22200
rect 18984 20318 19104 20346
rect 18984 20058 19012 20318
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 19076 19854 19104 20198
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19338 19272 19394 19281
rect 19338 19207 19340 19216
rect 19392 19207 19394 19216
rect 19444 19224 19472 19654
rect 19536 19281 19564 22200
rect 19996 19802 20024 22200
rect 19904 19774 20024 19802
rect 19904 19310 19932 19774
rect 19892 19304 19944 19310
rect 19522 19272 19578 19281
rect 19444 19196 19492 19224
rect 19892 19246 19944 19252
rect 19522 19207 19578 19216
rect 19340 19178 19392 19184
rect 19464 19156 19492 19196
rect 19616 19168 19668 19174
rect 19464 19128 19555 19156
rect 19527 19122 19555 19128
rect 19527 19094 19564 19122
rect 19616 19110 19668 19116
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18708 18737 18736 18906
rect 18694 18728 18750 18737
rect 18694 18663 18750 18672
rect 19340 18692 19392 18698
rect 19536 18680 19564 19094
rect 19392 18652 19564 18680
rect 19340 18634 19392 18640
rect 19628 18290 19656 19110
rect 19720 18698 19748 19110
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19616 18284 19668 18290
rect 19668 18244 19748 18272
rect 19616 18226 19668 18232
rect 18510 18184 18566 18193
rect 18510 18119 18566 18128
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 18602 17776 18658 17785
rect 18602 17711 18658 17720
rect 19616 17740 19668 17746
rect 18234 17232 18290 17241
rect 18144 17196 18196 17202
rect 18234 17167 18290 17176
rect 18144 17138 18196 17144
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 18156 15366 18184 17138
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18248 16522 18276 16934
rect 18236 16516 18288 16522
rect 18236 16458 18288 16464
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17972 14822 18000 14962
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17960 14544 18012 14550
rect 17958 14512 17960 14521
rect 18012 14512 18014 14521
rect 17958 14447 18014 14456
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 16776 10696 17172 10724
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 10266 15792 10406
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 16132 10062 16160 10542
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 16132 9722 16160 9998
rect 16776 9926 16804 10696
rect 17236 10674 17264 11766
rect 17328 11082 17356 14214
rect 17420 14074 17448 14282
rect 17696 14074 17724 14282
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17696 13433 17724 14010
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 17682 13424 17738 13433
rect 17682 13359 17738 13368
rect 18064 13326 18092 13670
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18064 12850 18092 13262
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 15842 9480 15898 9489
rect 15842 9415 15844 9424
rect 15896 9415 15898 9424
rect 15844 9386 15896 9392
rect 16132 9382 16160 9658
rect 16960 9450 16988 9862
rect 17236 9722 17264 10610
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17880 10169 17908 10406
rect 17866 10160 17922 10169
rect 17866 10095 17922 10104
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17420 9722 17448 9998
rect 17880 9994 17908 10095
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 18156 9625 18184 15302
rect 18248 14278 18276 16458
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18340 15910 18368 16050
rect 18328 15904 18380 15910
rect 18328 15846 18380 15852
rect 18340 15502 18368 15846
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 18340 15026 18368 15438
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18340 11014 18368 14758
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18432 10742 18460 11494
rect 18420 10736 18472 10742
rect 18420 10678 18472 10684
rect 18432 9654 18460 10678
rect 18420 9648 18472 9654
rect 18142 9616 18198 9625
rect 18420 9590 18472 9596
rect 18142 9551 18198 9560
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16132 8838 16160 9318
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 18524 8566 18552 12038
rect 18616 10266 18644 17711
rect 19616 17682 19668 17688
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18696 17060 18748 17066
rect 18696 17002 18748 17008
rect 18708 16182 18736 17002
rect 19076 16998 19104 17478
rect 19628 17270 19656 17682
rect 19720 17542 19748 18244
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 18880 16584 18932 16590
rect 18880 16526 18932 16532
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 18892 16114 18920 16526
rect 18984 16182 19012 16934
rect 19076 16658 19104 16934
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19430 16688 19486 16697
rect 19064 16652 19116 16658
rect 19430 16623 19486 16632
rect 19064 16594 19116 16600
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18984 15366 19012 16118
rect 19444 15994 19472 16623
rect 19536 16590 19564 16934
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19536 16250 19564 16526
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19444 15966 19564 15994
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13266 8120 13322 8129
rect 13945 8123 14253 8132
rect 13266 8055 13268 8064
rect 13320 8055 13322 8064
rect 13268 8026 13320 8032
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 18708 7546 18736 14214
rect 18786 13832 18842 13841
rect 18786 13767 18842 13776
rect 18800 11830 18828 13767
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18892 12918 18920 13398
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18892 12102 18920 12854
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18788 11824 18840 11830
rect 18788 11766 18840 11772
rect 18800 11354 18828 11766
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18892 11121 18920 12038
rect 18878 11112 18934 11121
rect 18878 11047 18934 11056
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 18984 6662 19012 15302
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19062 13832 19118 13841
rect 19062 13767 19118 13776
rect 19076 13734 19104 13767
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19536 13530 19564 15966
rect 19616 15496 19668 15502
rect 19614 15464 19616 15473
rect 19668 15464 19670 15473
rect 19614 15399 19670 15408
rect 19720 15314 19748 17478
rect 20088 17354 20116 22222
rect 20364 22114 20392 22222
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 20456 22114 20484 22200
rect 20364 22086 20484 22114
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 19904 17326 20116 17354
rect 19628 15286 19748 15314
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19628 15065 19656 15286
rect 19614 15056 19670 15065
rect 19614 14991 19670 15000
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19720 14618 19748 14962
rect 19812 14822 19840 15302
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19708 14612 19760 14618
rect 19708 14554 19760 14560
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19352 12986 19380 13194
rect 19616 13184 19668 13190
rect 19616 13126 19668 13132
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 19076 11762 19104 12174
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 19076 11218 19104 11698
rect 19260 11665 19288 12378
rect 19628 11898 19656 13126
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19246 11656 19302 11665
rect 19246 11591 19302 11600
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19522 11248 19578 11257
rect 19064 11212 19116 11218
rect 19522 11183 19578 11192
rect 19064 11154 19116 11160
rect 19536 11150 19564 11183
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 19076 9178 19104 9998
rect 19536 9654 19564 11086
rect 19628 10266 19656 11290
rect 19720 10810 19748 14418
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19812 12986 19840 14010
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19800 9988 19852 9994
rect 19800 9930 19852 9936
rect 19812 9722 19840 9930
rect 19800 9716 19852 9722
rect 19800 9658 19852 9664
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19904 6798 19932 17326
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19996 13258 20024 14758
rect 20180 14482 20208 19722
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18290 20300 18566
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20272 17882 20300 18226
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20732 17678 20760 19654
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20824 17610 20852 19314
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20916 17338 20944 22200
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 20996 19780 21048 19786
rect 20996 19722 21048 19728
rect 21008 18426 21036 19722
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21100 18766 21128 19246
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20456 14346 20484 15846
rect 20640 15434 20668 16390
rect 20824 15910 20852 16526
rect 21086 16008 21142 16017
rect 21086 15943 21088 15952
rect 21140 15943 21142 15952
rect 21088 15914 21140 15920
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20824 15502 20852 15846
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20628 15428 20680 15434
rect 20628 15370 20680 15376
rect 20824 15094 20852 15438
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20824 14346 20852 15030
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20180 13530 20208 13874
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 20076 13252 20128 13258
rect 20076 13194 20128 13200
rect 20088 10810 20116 13194
rect 20732 12434 20760 14010
rect 20824 13938 20852 14282
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20824 13326 20852 13874
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 21100 13258 21128 15914
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 20732 12406 20852 12434
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11762 20484 12038
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 20456 10554 20484 11698
rect 20824 11354 20852 12406
rect 21088 12164 21140 12170
rect 21088 12106 21140 12112
rect 21100 11898 21128 12106
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20534 10568 20590 10577
rect 20456 10526 20534 10554
rect 20534 10503 20590 10512
rect 20548 9654 20576 10503
rect 20720 10056 20772 10062
rect 21100 10033 21128 10610
rect 20720 9998 20772 10004
rect 21086 10024 21142 10033
rect 20732 9722 20760 9998
rect 21086 9959 21142 9968
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 21100 8634 21128 9959
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 21192 5098 21220 20742
rect 21376 20482 21404 22200
rect 21836 20806 21864 22200
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21376 20454 21496 20482
rect 22296 20466 22324 22200
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21376 19854 21404 20334
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21376 19310 21404 19790
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21376 17134 21404 17614
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21376 16590 21404 17070
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21284 12238 21312 12718
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21284 11762 21312 12174
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21284 11354 21312 11698
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21284 10674 21312 11290
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21284 10062 21312 10610
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21362 10024 21418 10033
rect 21362 9959 21418 9968
rect 21376 9926 21404 9959
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21272 8900 21324 8906
rect 21272 8842 21324 8848
rect 21284 8634 21312 8842
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21468 6458 21496 20454
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 22756 18970 22784 22200
rect 22744 18964 22796 18970
rect 22744 18906 22796 18912
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 21560 6730 21588 17274
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21180 5092 21232 5098
rect 21180 5034 21232 5040
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 12084 2746 12204 2774
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 2872 1828 2924 1834
rect 2872 1770 2924 1776
rect 5540 1828 5592 1834
rect 5540 1770 5592 1776
rect 2884 1737 2912 1770
rect 2870 1728 2926 1737
rect 2870 1663 2926 1672
rect 12084 898 12112 2746
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 11440 870 11560 898
rect 11440 800 11468 870
rect 11426 0 11482 800
rect 11532 762 11560 870
rect 11808 870 12112 898
rect 11808 762 11836 870
rect 11532 734 11836 762
<< via2 >>
rect 1490 20052 1546 20088
rect 1490 20032 1492 20052
rect 1492 20032 1544 20052
rect 1544 20032 1546 20052
rect 1950 21256 2006 21312
rect 2042 20440 2098 20496
rect 1950 19624 2006 19680
rect 1950 17992 2006 18048
rect 1950 17584 2006 17640
rect 1766 17448 1822 17504
rect 1674 16632 1730 16688
rect 1582 13096 1638 13152
rect 1950 17176 2006 17232
rect 1858 16768 1914 16824
rect 2778 20848 2834 20904
rect 2318 18844 2320 18864
rect 2320 18844 2372 18864
rect 2372 18844 2374 18864
rect 2318 18808 2374 18844
rect 2410 18400 2466 18456
rect 1950 15952 2006 16008
rect 2870 19216 2926 19272
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3238 18148 3294 18184
rect 3238 18128 3240 18148
rect 3240 18128 3292 18148
rect 3292 18128 3294 18148
rect 2870 16360 2926 16416
rect 2502 15544 2558 15600
rect 2042 14728 2098 14784
rect 2134 13504 2190 13560
rect 2410 12280 2466 12336
rect 2962 15136 3018 15192
rect 2870 14320 2926 14376
rect 2778 13912 2834 13968
rect 3054 13232 3110 13288
rect 3146 12144 3202 12200
rect 1490 7792 1546 7848
rect 3146 11464 3202 11520
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3330 15408 3386 15464
rect 3238 11056 3294 11112
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3882 12688 3938 12744
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3882 11872 3938 11928
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3514 11076 3570 11112
rect 3514 11056 3516 11076
rect 3516 11056 3568 11076
rect 3568 11056 3570 11076
rect 3882 11056 3938 11112
rect 3422 10648 3478 10704
rect 3606 10668 3662 10704
rect 5446 19352 5502 19408
rect 4434 15000 4490 15056
rect 5170 16904 5226 16960
rect 3606 10648 3608 10668
rect 3608 10648 3660 10668
rect 3660 10648 3662 10668
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3422 10240 3478 10296
rect 3330 9832 3386 9888
rect 3974 9424 4030 9480
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 4066 9016 4122 9072
rect 3974 8608 4030 8664
rect 3054 8200 3110 8256
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 2778 7384 2834 7440
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3422 6996 3478 7032
rect 3422 6976 3424 6996
rect 3424 6976 3476 6996
rect 3476 6976 3478 6996
rect 4066 6568 4122 6624
rect 4066 6196 4068 6216
rect 4068 6196 4120 6216
rect 4120 6196 4122 6216
rect 4066 6160 4122 6196
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 4066 5752 4122 5808
rect 4066 5364 4122 5400
rect 4066 5344 4068 5364
rect 4068 5344 4120 5364
rect 4120 5344 4122 5364
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 4158 5072 4214 5128
rect 5262 15952 5318 16008
rect 5446 15000 5502 15056
rect 5170 13912 5226 13968
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6090 17740 6146 17776
rect 6090 17720 6092 17740
rect 6092 17720 6144 17740
rect 6144 17720 6146 17740
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 5814 17176 5870 17232
rect 5446 13368 5502 13424
rect 5170 12824 5226 12880
rect 4986 12300 5042 12336
rect 4986 12280 4988 12300
rect 4988 12280 5040 12300
rect 5040 12280 5042 12300
rect 5538 10512 5594 10568
rect 6826 20204 6828 20224
rect 6828 20204 6880 20224
rect 6880 20204 6882 20224
rect 6826 20168 6882 20204
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 7286 19352 7342 19408
rect 7194 16652 7250 16688
rect 7194 16632 7196 16652
rect 7196 16632 7248 16652
rect 7248 16632 7250 16652
rect 6734 16360 6790 16416
rect 6550 15272 6606 15328
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6090 14728 6146 14784
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 7010 14900 7012 14920
rect 7012 14900 7064 14920
rect 7064 14900 7066 14920
rect 7010 14864 7066 14900
rect 7010 13912 7066 13968
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6642 11600 6698 11656
rect 6182 11212 6238 11248
rect 6182 11192 6184 11212
rect 6184 11192 6236 11212
rect 6236 11192 6238 11212
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 5998 10104 6054 10160
rect 6734 10648 6790 10704
rect 7102 13232 7158 13288
rect 7654 16360 7710 16416
rect 7470 14592 7526 14648
rect 6918 11600 6974 11656
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 5170 9036 5226 9072
rect 5170 9016 5172 9036
rect 5172 9016 5224 9036
rect 5224 9016 5226 9036
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 4434 4528 4490 4584
rect 3974 4120 4030 4176
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3422 3712 3478 3768
rect 4066 3304 4122 3360
rect 3974 2896 4030 2952
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 4066 2524 4068 2544
rect 4068 2524 4120 2544
rect 4120 2524 4122 2544
rect 4066 2488 4122 2524
rect 3514 2080 3570 2136
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 8022 17856 8078 17912
rect 8022 16652 8078 16688
rect 8022 16632 8024 16652
rect 8024 16632 8076 16652
rect 8076 16632 8078 16652
rect 8022 15564 8078 15600
rect 8022 15544 8024 15564
rect 8024 15544 8076 15564
rect 8076 15544 8078 15564
rect 7930 15136 7986 15192
rect 7838 14456 7894 14512
rect 7838 11756 7894 11792
rect 7838 11736 7840 11756
rect 7840 11736 7892 11756
rect 7892 11736 7894 11756
rect 7838 9716 7894 9752
rect 7838 9696 7840 9716
rect 7840 9696 7892 9716
rect 7892 9696 7894 9716
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8390 15272 8446 15328
rect 8390 14728 8446 14784
rect 8482 14592 8538 14648
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 9034 16360 9090 16416
rect 8666 16088 8722 16144
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8666 15580 8668 15600
rect 8668 15580 8720 15600
rect 8720 15580 8722 15600
rect 8666 15544 8722 15580
rect 8850 15408 8906 15464
rect 8206 12724 8208 12744
rect 8208 12724 8260 12744
rect 8260 12724 8262 12744
rect 8206 12688 8262 12724
rect 8022 12144 8078 12200
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 9402 19932 9404 19952
rect 9404 19932 9456 19952
rect 9456 19932 9458 19952
rect 9402 19896 9458 19932
rect 9310 19216 9366 19272
rect 9310 16088 9366 16144
rect 9494 15136 9550 15192
rect 9402 13504 9458 13560
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 9034 9560 9090 9616
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 9678 13640 9734 13696
rect 9862 15408 9918 15464
rect 10046 11636 10048 11656
rect 10048 11636 10100 11656
rect 10100 11636 10102 11656
rect 10046 11600 10102 11636
rect 10598 18672 10654 18728
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 10966 18264 11022 18320
rect 10322 9016 10378 9072
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11150 13640 11206 13696
rect 11150 13096 11206 13152
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11242 12280 11298 12336
rect 11886 17484 11888 17504
rect 11888 17484 11940 17504
rect 11940 17484 11942 17504
rect 11886 17448 11942 17484
rect 12438 18808 12494 18864
rect 12438 18536 12494 18592
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 12622 17992 12678 18048
rect 11978 13232 12034 13288
rect 11150 12008 11206 12064
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 12530 17176 12586 17232
rect 12530 16632 12586 16688
rect 12162 11736 12218 11792
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 12622 13640 12678 13696
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13358 17040 13414 17096
rect 12898 12824 12954 12880
rect 12898 12144 12954 12200
rect 14186 18572 14188 18592
rect 14188 18572 14240 18592
rect 14240 18572 14242 18592
rect 14186 18536 14242 18572
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 14186 17448 14242 17504
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13634 16496 13690 16552
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 14278 14456 14334 14512
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 14554 13096 14610 13152
rect 14278 11192 14334 11248
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 15382 18808 15438 18864
rect 14738 12144 14794 12200
rect 15106 14456 15162 14512
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 17222 19896 17278 19952
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 18142 19216 18198 19272
rect 15106 13232 15162 13288
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 15842 14864 15898 14920
rect 15474 12688 15530 12744
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 17958 17584 18014 17640
rect 18418 18264 18474 18320
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19338 19236 19394 19272
rect 19338 19216 19340 19236
rect 19340 19216 19392 19236
rect 19392 19216 19394 19236
rect 19522 19216 19578 19272
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 18694 18672 18750 18728
rect 18510 18128 18566 18184
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 18602 17720 18658 17776
rect 18234 17176 18290 17232
rect 17958 14492 17960 14512
rect 17960 14492 18012 14512
rect 18012 14492 18014 14512
rect 17958 14456 18014 14492
rect 17682 13368 17738 13424
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 15842 9444 15898 9480
rect 15842 9424 15844 9444
rect 15844 9424 15896 9444
rect 15896 9424 15898 9444
rect 17866 10104 17922 10160
rect 18142 9560 18198 9616
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19430 16632 19486 16688
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13266 8084 13322 8120
rect 13266 8064 13268 8084
rect 13268 8064 13320 8084
rect 13320 8064 13322 8084
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 18786 13776 18842 13832
rect 18878 11056 18934 11112
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19062 13776 19118 13832
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19614 15444 19616 15464
rect 19616 15444 19668 15464
rect 19668 15444 19670 15464
rect 19614 15408 19670 15444
rect 19614 15000 19670 15056
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19246 11600 19302 11656
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19522 11192 19578 11248
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 21086 15972 21142 16008
rect 21086 15952 21088 15972
rect 21088 15952 21140 15972
rect 21140 15952 21142 15972
rect 20534 10512 20590 10568
rect 21086 9968 21142 10024
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21362 9968 21418 10024
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 2870 1672 2926 1728
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 0 21314 800 21344
rect 1945 21314 2011 21317
rect 0 21312 2011 21314
rect 0 21256 1950 21312
rect 2006 21256 2011 21312
rect 0 21254 2011 21256
rect 0 21224 800 21254
rect 1945 21251 2011 21254
rect 0 20906 800 20936
rect 2773 20906 2839 20909
rect 0 20904 2839 20906
rect 0 20848 2778 20904
rect 2834 20848 2839 20904
rect 0 20846 2839 20848
rect 0 20816 800 20846
rect 2773 20843 2839 20846
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 0 20498 800 20528
rect 2037 20498 2103 20501
rect 0 20496 2103 20498
rect 0 20440 2042 20496
rect 2098 20440 2103 20496
rect 0 20438 2103 20440
rect 0 20408 800 20438
rect 2037 20435 2103 20438
rect 6821 20228 6887 20229
rect 6821 20226 6868 20228
rect 6776 20224 6868 20226
rect 6776 20168 6826 20224
rect 6776 20166 6868 20168
rect 6821 20164 6868 20166
rect 6932 20164 6938 20228
rect 6821 20163 6887 20164
rect 3545 20160 3861 20161
rect 0 20090 800 20120
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 1485 20090 1551 20093
rect 0 20088 1551 20090
rect 0 20032 1490 20088
rect 1546 20032 1551 20088
rect 0 20030 1551 20032
rect 0 20000 800 20030
rect 1485 20027 1551 20030
rect 9397 19954 9463 19957
rect 17217 19954 17283 19957
rect 9397 19952 17283 19954
rect 9397 19896 9402 19952
rect 9458 19896 17222 19952
rect 17278 19896 17283 19952
rect 9397 19894 17283 19896
rect 9397 19891 9463 19894
rect 17217 19891 17283 19894
rect 0 19682 800 19712
rect 1945 19682 2011 19685
rect 0 19680 2011 19682
rect 0 19624 1950 19680
rect 2006 19624 2011 19680
rect 0 19622 2011 19624
rect 0 19592 800 19622
rect 1945 19619 2011 19622
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 5441 19410 5507 19413
rect 7281 19410 7347 19413
rect 5441 19408 7347 19410
rect 5441 19352 5446 19408
rect 5502 19352 7286 19408
rect 7342 19352 7347 19408
rect 5441 19350 7347 19352
rect 5441 19347 5507 19350
rect 7281 19347 7347 19350
rect 0 19274 800 19304
rect 2865 19274 2931 19277
rect 0 19272 2931 19274
rect 0 19216 2870 19272
rect 2926 19216 2931 19272
rect 0 19214 2931 19216
rect 0 19184 800 19214
rect 2865 19211 2931 19214
rect 9305 19274 9371 19277
rect 18137 19274 18203 19277
rect 9305 19272 18203 19274
rect 9305 19216 9310 19272
rect 9366 19216 18142 19272
rect 18198 19216 18203 19272
rect 9305 19214 18203 19216
rect 9305 19211 9371 19214
rect 18137 19211 18203 19214
rect 19333 19274 19399 19277
rect 19517 19274 19583 19277
rect 19333 19272 19583 19274
rect 19333 19216 19338 19272
rect 19394 19216 19522 19272
rect 19578 19216 19583 19272
rect 19333 19214 19583 19216
rect 19333 19211 19399 19214
rect 19517 19211 19583 19214
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 0 18866 800 18896
rect 2313 18866 2379 18869
rect 0 18864 2379 18866
rect 0 18808 2318 18864
rect 2374 18808 2379 18864
rect 0 18806 2379 18808
rect 0 18776 800 18806
rect 2313 18803 2379 18806
rect 12433 18866 12499 18869
rect 15377 18866 15443 18869
rect 12433 18864 15443 18866
rect 12433 18808 12438 18864
rect 12494 18808 15382 18864
rect 15438 18808 15443 18864
rect 12433 18806 15443 18808
rect 12433 18803 12499 18806
rect 15377 18803 15443 18806
rect 10593 18730 10659 18733
rect 18689 18730 18755 18733
rect 10593 18728 18755 18730
rect 10593 18672 10598 18728
rect 10654 18672 18694 18728
rect 18750 18672 18755 18728
rect 10593 18670 18755 18672
rect 10593 18667 10659 18670
rect 18689 18667 18755 18670
rect 12433 18594 12499 18597
rect 14181 18594 14247 18597
rect 12433 18592 14247 18594
rect 12433 18536 12438 18592
rect 12494 18536 14186 18592
rect 14242 18536 14247 18592
rect 12433 18534 14247 18536
rect 12433 18531 12499 18534
rect 14181 18531 14247 18534
rect 6144 18528 6460 18529
rect 0 18458 800 18488
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 2405 18458 2471 18461
rect 0 18456 2471 18458
rect 0 18400 2410 18456
rect 2466 18400 2471 18456
rect 0 18398 2471 18400
rect 0 18368 800 18398
rect 2405 18395 2471 18398
rect 10961 18322 11027 18325
rect 18413 18322 18479 18325
rect 10961 18320 18479 18322
rect 10961 18264 10966 18320
rect 11022 18264 18418 18320
rect 18474 18264 18479 18320
rect 10961 18262 18479 18264
rect 10961 18259 11027 18262
rect 18413 18259 18479 18262
rect 3233 18186 3299 18189
rect 18505 18186 18571 18189
rect 3233 18184 18571 18186
rect 3233 18128 3238 18184
rect 3294 18128 18510 18184
rect 18566 18128 18571 18184
rect 3233 18126 18571 18128
rect 3233 18123 3299 18126
rect 18505 18123 18571 18126
rect 0 18050 800 18080
rect 1945 18050 2011 18053
rect 0 18048 2011 18050
rect 0 17992 1950 18048
rect 2006 17992 2011 18048
rect 0 17990 2011 17992
rect 0 17960 800 17990
rect 1945 17987 2011 17990
rect 12617 18050 12683 18053
rect 13302 18050 13308 18052
rect 12617 18048 13308 18050
rect 12617 17992 12622 18048
rect 12678 17992 13308 18048
rect 12617 17990 13308 17992
rect 12617 17987 12683 17990
rect 13302 17988 13308 17990
rect 13372 17988 13378 18052
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 8017 17916 8083 17917
rect 7966 17914 7972 17916
rect 7926 17854 7972 17914
rect 8036 17912 8083 17916
rect 8078 17856 8083 17912
rect 7966 17852 7972 17854
rect 8036 17852 8083 17856
rect 8017 17851 8083 17852
rect 6085 17778 6151 17781
rect 18597 17778 18663 17781
rect 6085 17776 18663 17778
rect 6085 17720 6090 17776
rect 6146 17720 18602 17776
rect 18658 17720 18663 17776
rect 6085 17718 18663 17720
rect 6085 17715 6151 17718
rect 18597 17715 18663 17718
rect 0 17642 800 17672
rect 1945 17642 2011 17645
rect 17953 17642 18019 17645
rect 0 17640 2011 17642
rect 0 17584 1950 17640
rect 2006 17584 2011 17640
rect 0 17582 2011 17584
rect 0 17552 800 17582
rect 1945 17579 2011 17582
rect 2086 17640 18019 17642
rect 2086 17584 17958 17640
rect 18014 17584 18019 17640
rect 2086 17582 18019 17584
rect 1761 17506 1827 17509
rect 2086 17506 2146 17582
rect 17953 17579 18019 17582
rect 1761 17504 2146 17506
rect 1761 17448 1766 17504
rect 1822 17448 2146 17504
rect 1761 17446 2146 17448
rect 11881 17506 11947 17509
rect 14181 17506 14247 17509
rect 11881 17504 14247 17506
rect 11881 17448 11886 17504
rect 11942 17448 14186 17504
rect 14242 17448 14247 17504
rect 11881 17446 14247 17448
rect 1761 17443 1827 17446
rect 11881 17443 11947 17446
rect 14181 17443 14247 17446
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 0 17234 800 17264
rect 1945 17234 2011 17237
rect 0 17232 2011 17234
rect 0 17176 1950 17232
rect 2006 17176 2011 17232
rect 0 17174 2011 17176
rect 0 17144 800 17174
rect 1945 17171 2011 17174
rect 5809 17234 5875 17237
rect 12525 17234 12591 17237
rect 18229 17234 18295 17237
rect 5809 17232 12591 17234
rect 5809 17176 5814 17232
rect 5870 17176 12530 17232
rect 12586 17176 12591 17232
rect 5809 17174 12591 17176
rect 5809 17171 5875 17174
rect 12525 17171 12591 17174
rect 12942 17232 18295 17234
rect 12942 17176 18234 17232
rect 18290 17176 18295 17232
rect 12942 17174 18295 17176
rect 12942 17098 13002 17174
rect 18229 17171 18295 17174
rect 2730 17038 13002 17098
rect 0 16826 800 16856
rect 1853 16826 1919 16829
rect 0 16824 1919 16826
rect 0 16768 1858 16824
rect 1914 16768 1919 16824
rect 0 16766 1919 16768
rect 0 16736 800 16766
rect 1853 16763 1919 16766
rect 1669 16690 1735 16693
rect 2730 16690 2790 17038
rect 13118 17036 13124 17100
rect 13188 17098 13194 17100
rect 13353 17098 13419 17101
rect 13188 17096 13419 17098
rect 13188 17040 13358 17096
rect 13414 17040 13419 17096
rect 13188 17038 13419 17040
rect 13188 17036 13194 17038
rect 13353 17035 13419 17038
rect 5165 16964 5231 16965
rect 5165 16962 5212 16964
rect 5120 16960 5212 16962
rect 5120 16904 5170 16960
rect 5120 16902 5212 16904
rect 5165 16900 5212 16902
rect 5276 16900 5282 16964
rect 5165 16899 5231 16900
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 7189 16692 7255 16693
rect 7189 16690 7236 16692
rect 1669 16688 2790 16690
rect 1669 16632 1674 16688
rect 1730 16632 2790 16688
rect 1669 16630 2790 16632
rect 7144 16688 7236 16690
rect 7144 16632 7194 16688
rect 7144 16630 7236 16632
rect 1669 16627 1735 16630
rect 7189 16628 7236 16630
rect 7300 16628 7306 16692
rect 8017 16690 8083 16693
rect 12525 16690 12591 16693
rect 19425 16690 19491 16693
rect 8017 16688 12450 16690
rect 8017 16632 8022 16688
rect 8078 16632 12450 16688
rect 8017 16630 12450 16632
rect 7189 16627 7255 16628
rect 8017 16627 8083 16630
rect 12390 16554 12450 16630
rect 12525 16688 19491 16690
rect 12525 16632 12530 16688
rect 12586 16632 19430 16688
rect 19486 16632 19491 16688
rect 12525 16630 19491 16632
rect 12525 16627 12591 16630
rect 19425 16627 19491 16630
rect 13629 16554 13695 16557
rect 12390 16552 13695 16554
rect 12390 16496 13634 16552
rect 13690 16496 13695 16552
rect 12390 16494 13695 16496
rect 13629 16491 13695 16494
rect 0 16418 800 16448
rect 2865 16418 2931 16421
rect 0 16416 2931 16418
rect 0 16360 2870 16416
rect 2926 16360 2931 16416
rect 0 16358 2931 16360
rect 0 16328 800 16358
rect 2865 16355 2931 16358
rect 6729 16418 6795 16421
rect 7649 16418 7715 16421
rect 9029 16418 9095 16421
rect 6729 16416 9095 16418
rect 6729 16360 6734 16416
rect 6790 16360 7654 16416
rect 7710 16360 9034 16416
rect 9090 16360 9095 16416
rect 6729 16358 9095 16360
rect 6729 16355 6795 16358
rect 7649 16355 7715 16358
rect 9029 16355 9095 16358
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 8661 16146 8727 16149
rect 9305 16146 9371 16149
rect 8661 16144 9371 16146
rect 8661 16088 8666 16144
rect 8722 16088 9310 16144
rect 9366 16088 9371 16144
rect 8661 16086 9371 16088
rect 8661 16083 8727 16086
rect 9305 16083 9371 16086
rect 0 16010 800 16040
rect 1945 16010 2011 16013
rect 0 16008 2011 16010
rect 0 15952 1950 16008
rect 2006 15952 2011 16008
rect 0 15950 2011 15952
rect 0 15920 800 15950
rect 1945 15947 2011 15950
rect 5257 16010 5323 16013
rect 21081 16010 21147 16013
rect 5257 16008 21147 16010
rect 5257 15952 5262 16008
rect 5318 15952 21086 16008
rect 21142 15952 21147 16008
rect 5257 15950 21147 15952
rect 5257 15947 5323 15950
rect 21081 15947 21147 15950
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 0 15602 800 15632
rect 2497 15602 2563 15605
rect 0 15600 2563 15602
rect 0 15544 2502 15600
rect 2558 15544 2563 15600
rect 0 15542 2563 15544
rect 0 15512 800 15542
rect 2497 15539 2563 15542
rect 8017 15602 8083 15605
rect 8661 15602 8727 15605
rect 8017 15600 8727 15602
rect 8017 15544 8022 15600
rect 8078 15544 8666 15600
rect 8722 15544 8727 15600
rect 8017 15542 8727 15544
rect 8017 15539 8083 15542
rect 8661 15539 8727 15542
rect 3325 15466 3391 15469
rect 8845 15466 8911 15469
rect 3325 15464 8911 15466
rect 3325 15408 3330 15464
rect 3386 15408 8850 15464
rect 8906 15408 8911 15464
rect 3325 15406 8911 15408
rect 3325 15403 3391 15406
rect 8845 15403 8911 15406
rect 9857 15466 9923 15469
rect 19609 15466 19675 15469
rect 9857 15464 19675 15466
rect 9857 15408 9862 15464
rect 9918 15408 19614 15464
rect 19670 15408 19675 15464
rect 9857 15406 19675 15408
rect 9857 15403 9923 15406
rect 19609 15403 19675 15406
rect 6545 15330 6611 15333
rect 8385 15330 8451 15333
rect 6545 15328 8451 15330
rect 6545 15272 6550 15328
rect 6606 15272 8390 15328
rect 8446 15272 8451 15328
rect 6545 15270 8451 15272
rect 6545 15267 6611 15270
rect 8385 15267 8451 15270
rect 6144 15264 6460 15265
rect 0 15194 800 15224
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 2957 15194 3023 15197
rect 0 15192 3023 15194
rect 0 15136 2962 15192
rect 3018 15136 3023 15192
rect 0 15134 3023 15136
rect 0 15104 800 15134
rect 2957 15131 3023 15134
rect 7925 15194 7991 15197
rect 9489 15194 9555 15197
rect 7925 15192 9555 15194
rect 7925 15136 7930 15192
rect 7986 15136 9494 15192
rect 9550 15136 9555 15192
rect 7925 15134 9555 15136
rect 7925 15131 7991 15134
rect 9489 15131 9555 15134
rect 4429 15058 4495 15061
rect 5441 15058 5507 15061
rect 19609 15058 19675 15061
rect 4429 15056 19675 15058
rect 4429 15000 4434 15056
rect 4490 15000 5446 15056
rect 5502 15000 19614 15056
rect 19670 15000 19675 15056
rect 4429 14998 19675 15000
rect 4429 14995 4495 14998
rect 5441 14995 5507 14998
rect 19609 14995 19675 14998
rect 7005 14922 7071 14925
rect 15837 14922 15903 14925
rect 7005 14920 15903 14922
rect 7005 14864 7010 14920
rect 7066 14864 15842 14920
rect 15898 14864 15903 14920
rect 7005 14862 15903 14864
rect 7005 14859 7071 14862
rect 15837 14859 15903 14862
rect 0 14786 800 14816
rect 2037 14786 2103 14789
rect 0 14784 2103 14786
rect 0 14728 2042 14784
rect 2098 14728 2103 14784
rect 0 14726 2103 14728
rect 0 14696 800 14726
rect 2037 14723 2103 14726
rect 6085 14786 6151 14789
rect 8385 14786 8451 14789
rect 6085 14784 8451 14786
rect 6085 14728 6090 14784
rect 6146 14728 8390 14784
rect 8446 14728 8451 14784
rect 6085 14726 8451 14728
rect 6085 14723 6151 14726
rect 8385 14723 8451 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 7465 14650 7531 14653
rect 8477 14650 8543 14653
rect 7465 14648 8543 14650
rect 7465 14592 7470 14648
rect 7526 14592 8482 14648
rect 8538 14592 8543 14648
rect 7465 14590 8543 14592
rect 7465 14587 7531 14590
rect 8477 14587 8543 14590
rect 7833 14514 7899 14517
rect 14273 14514 14339 14517
rect 7833 14512 14339 14514
rect 7833 14456 7838 14512
rect 7894 14456 14278 14512
rect 14334 14456 14339 14512
rect 7833 14454 14339 14456
rect 7833 14451 7899 14454
rect 14273 14451 14339 14454
rect 15101 14514 15167 14517
rect 17953 14514 18019 14517
rect 15101 14512 18019 14514
rect 15101 14456 15106 14512
rect 15162 14456 17958 14512
rect 18014 14456 18019 14512
rect 15101 14454 18019 14456
rect 15101 14451 15167 14454
rect 17953 14451 18019 14454
rect 0 14378 800 14408
rect 2865 14378 2931 14381
rect 0 14376 2931 14378
rect 0 14320 2870 14376
rect 2926 14320 2931 14376
rect 0 14318 2931 14320
rect 0 14288 800 14318
rect 2865 14315 2931 14318
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 0 13970 800 14000
rect 2773 13970 2839 13973
rect 0 13968 2839 13970
rect 0 13912 2778 13968
rect 2834 13912 2839 13968
rect 0 13910 2839 13912
rect 0 13880 800 13910
rect 2773 13907 2839 13910
rect 5165 13970 5231 13973
rect 7005 13970 7071 13973
rect 5165 13968 7071 13970
rect 5165 13912 5170 13968
rect 5226 13912 7010 13968
rect 7066 13912 7071 13968
rect 5165 13910 7071 13912
rect 5165 13907 5231 13910
rect 7005 13907 7071 13910
rect 6862 13772 6868 13836
rect 6932 13834 6938 13836
rect 18781 13834 18847 13837
rect 19057 13834 19123 13837
rect 6932 13832 19123 13834
rect 6932 13776 18786 13832
rect 18842 13776 19062 13832
rect 19118 13776 19123 13832
rect 6932 13774 19123 13776
rect 6932 13772 6938 13774
rect 18781 13771 18847 13774
rect 19057 13771 19123 13774
rect 9673 13698 9739 13701
rect 11145 13698 11211 13701
rect 12617 13698 12683 13701
rect 9673 13696 11211 13698
rect 9673 13640 9678 13696
rect 9734 13640 11150 13696
rect 11206 13640 11211 13696
rect 9673 13638 11211 13640
rect 9673 13635 9739 13638
rect 11145 13635 11211 13638
rect 12390 13696 12683 13698
rect 12390 13640 12622 13696
rect 12678 13640 12683 13696
rect 12390 13638 12683 13640
rect 3545 13632 3861 13633
rect 0 13562 800 13592
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 2129 13562 2195 13565
rect 0 13560 2195 13562
rect 0 13504 2134 13560
rect 2190 13504 2195 13560
rect 0 13502 2195 13504
rect 0 13472 800 13502
rect 2129 13499 2195 13502
rect 9397 13562 9463 13565
rect 12390 13562 12450 13638
rect 12617 13635 12683 13638
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 9397 13560 12450 13562
rect 9397 13504 9402 13560
rect 9458 13504 12450 13560
rect 9397 13502 12450 13504
rect 9397 13499 9463 13502
rect 5441 13426 5507 13429
rect 17677 13426 17743 13429
rect 5441 13424 17743 13426
rect 5441 13368 5446 13424
rect 5502 13368 17682 13424
rect 17738 13368 17743 13424
rect 5441 13366 17743 13368
rect 5441 13363 5507 13366
rect 17677 13363 17743 13366
rect 3049 13290 3115 13293
rect 7097 13290 7163 13293
rect 11973 13290 12039 13293
rect 15101 13290 15167 13293
rect 3049 13288 6746 13290
rect 3049 13232 3054 13288
rect 3110 13232 6746 13288
rect 3049 13230 6746 13232
rect 3049 13227 3115 13230
rect 0 13154 800 13184
rect 1577 13154 1643 13157
rect 0 13152 1643 13154
rect 0 13096 1582 13152
rect 1638 13096 1643 13152
rect 0 13094 1643 13096
rect 6686 13154 6746 13230
rect 7097 13288 11898 13290
rect 7097 13232 7102 13288
rect 7158 13232 11898 13288
rect 7097 13230 11898 13232
rect 7097 13227 7163 13230
rect 11145 13154 11211 13157
rect 6686 13152 11211 13154
rect 6686 13096 11150 13152
rect 11206 13096 11211 13152
rect 6686 13094 11211 13096
rect 11838 13154 11898 13230
rect 11973 13288 15167 13290
rect 11973 13232 11978 13288
rect 12034 13232 15106 13288
rect 15162 13232 15167 13288
rect 11973 13230 15167 13232
rect 11973 13227 12039 13230
rect 15101 13227 15167 13230
rect 14549 13154 14615 13157
rect 11838 13152 14615 13154
rect 11838 13096 14554 13152
rect 14610 13096 14615 13152
rect 11838 13094 14615 13096
rect 0 13064 800 13094
rect 1577 13091 1643 13094
rect 11145 13091 11211 13094
rect 14549 13091 14615 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 5165 12882 5231 12885
rect 12893 12882 12959 12885
rect 5165 12880 12959 12882
rect 5165 12824 5170 12880
rect 5226 12824 12898 12880
rect 12954 12824 12959 12880
rect 5165 12822 12959 12824
rect 5165 12819 5231 12822
rect 12893 12819 12959 12822
rect 0 12746 800 12776
rect 3877 12746 3943 12749
rect 0 12744 3943 12746
rect 0 12688 3882 12744
rect 3938 12688 3943 12744
rect 0 12686 3943 12688
rect 0 12656 800 12686
rect 3877 12683 3943 12686
rect 8201 12746 8267 12749
rect 15469 12746 15535 12749
rect 8201 12744 15535 12746
rect 8201 12688 8206 12744
rect 8262 12688 15474 12744
rect 15530 12688 15535 12744
rect 8201 12686 15535 12688
rect 8201 12683 8267 12686
rect 15469 12683 15535 12686
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 0 12338 800 12368
rect 2405 12338 2471 12341
rect 4981 12338 5047 12341
rect 11237 12338 11303 12341
rect 0 12278 2330 12338
rect 0 12248 800 12278
rect 2270 12202 2330 12278
rect 2405 12336 4906 12338
rect 2405 12280 2410 12336
rect 2466 12280 4906 12336
rect 2405 12278 4906 12280
rect 2405 12275 2471 12278
rect 3141 12202 3207 12205
rect 2270 12200 3207 12202
rect 2270 12144 3146 12200
rect 3202 12144 3207 12200
rect 2270 12142 3207 12144
rect 4846 12202 4906 12278
rect 4981 12336 11303 12338
rect 4981 12280 4986 12336
rect 5042 12280 11242 12336
rect 11298 12280 11303 12336
rect 4981 12278 11303 12280
rect 4981 12275 5047 12278
rect 11237 12275 11303 12278
rect 8017 12202 8083 12205
rect 12893 12202 12959 12205
rect 14733 12202 14799 12205
rect 4846 12142 6746 12202
rect 3141 12139 3207 12142
rect 6686 12066 6746 12142
rect 8017 12200 14799 12202
rect 8017 12144 8022 12200
rect 8078 12144 12898 12200
rect 12954 12144 14738 12200
rect 14794 12144 14799 12200
rect 8017 12142 14799 12144
rect 8017 12139 8083 12142
rect 12893 12139 12959 12142
rect 14733 12139 14799 12142
rect 11145 12066 11211 12069
rect 6686 12064 11211 12066
rect 6686 12008 11150 12064
rect 11206 12008 11211 12064
rect 6686 12006 11211 12008
rect 11145 12003 11211 12006
rect 6144 12000 6460 12001
rect 0 11930 800 11960
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 3877 11930 3943 11933
rect 0 11928 3943 11930
rect 0 11872 3882 11928
rect 3938 11872 3943 11928
rect 0 11870 3943 11872
rect 0 11840 800 11870
rect 3877 11867 3943 11870
rect 7833 11794 7899 11797
rect 12157 11794 12223 11797
rect 7833 11792 12223 11794
rect 7833 11736 7838 11792
rect 7894 11736 12162 11792
rect 12218 11736 12223 11792
rect 7833 11734 12223 11736
rect 7833 11731 7899 11734
rect 12157 11731 12223 11734
rect 6637 11658 6703 11661
rect 6913 11658 6979 11661
rect 10041 11658 10107 11661
rect 6637 11656 10107 11658
rect 6637 11600 6642 11656
rect 6698 11600 6918 11656
rect 6974 11600 10046 11656
rect 10102 11600 10107 11656
rect 6637 11598 10107 11600
rect 6637 11595 6703 11598
rect 6913 11595 6979 11598
rect 10041 11595 10107 11598
rect 19241 11658 19307 11661
rect 19241 11656 19626 11658
rect 19241 11600 19246 11656
rect 19302 11600 19626 11656
rect 19241 11598 19626 11600
rect 19241 11595 19307 11598
rect 0 11522 800 11552
rect 3141 11522 3207 11525
rect 0 11520 3207 11522
rect 0 11464 3146 11520
rect 3202 11464 3207 11520
rect 0 11462 3207 11464
rect 19566 11522 19626 11598
rect 22200 11522 23000 11552
rect 19566 11462 23000 11522
rect 0 11432 800 11462
rect 3141 11459 3207 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 22200 11432 23000 11462
rect 19139 11391 19455 11392
rect 6177 11250 6243 11253
rect 13118 11250 13124 11252
rect 6177 11248 13124 11250
rect 6177 11192 6182 11248
rect 6238 11192 13124 11248
rect 6177 11190 13124 11192
rect 6177 11187 6243 11190
rect 13118 11188 13124 11190
rect 13188 11188 13194 11252
rect 14273 11250 14339 11253
rect 19517 11250 19583 11253
rect 14273 11248 19583 11250
rect 14273 11192 14278 11248
rect 14334 11192 19522 11248
rect 19578 11192 19583 11248
rect 14273 11190 19583 11192
rect 14273 11187 14339 11190
rect 19517 11187 19583 11190
rect 0 11114 800 11144
rect 3233 11114 3299 11117
rect 0 11112 3299 11114
rect 0 11056 3238 11112
rect 3294 11056 3299 11112
rect 0 11054 3299 11056
rect 0 11024 800 11054
rect 3233 11051 3299 11054
rect 3509 11114 3575 11117
rect 3877 11114 3943 11117
rect 18873 11114 18939 11117
rect 3509 11112 18939 11114
rect 3509 11056 3514 11112
rect 3570 11056 3882 11112
rect 3938 11056 18878 11112
rect 18934 11056 18939 11112
rect 3509 11054 18939 11056
rect 3509 11051 3575 11054
rect 3877 11051 3943 11054
rect 18873 11051 18939 11054
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 0 10706 800 10736
rect 3417 10706 3483 10709
rect 0 10704 3483 10706
rect 0 10648 3422 10704
rect 3478 10648 3483 10704
rect 0 10646 3483 10648
rect 0 10616 800 10646
rect 3417 10643 3483 10646
rect 3601 10706 3667 10709
rect 6729 10706 6795 10709
rect 3601 10704 6795 10706
rect 3601 10648 3606 10704
rect 3662 10648 6734 10704
rect 6790 10648 6795 10704
rect 3601 10646 6795 10648
rect 3601 10643 3667 10646
rect 6729 10643 6795 10646
rect 5533 10570 5599 10573
rect 20529 10570 20595 10573
rect 5533 10568 20595 10570
rect 5533 10512 5538 10568
rect 5594 10512 20534 10568
rect 20590 10512 20595 10568
rect 5533 10510 20595 10512
rect 5533 10507 5599 10510
rect 20529 10507 20595 10510
rect 3545 10368 3861 10369
rect 0 10298 800 10328
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 3417 10298 3483 10301
rect 0 10296 3483 10298
rect 0 10240 3422 10296
rect 3478 10240 3483 10296
rect 0 10238 3483 10240
rect 0 10208 800 10238
rect 3417 10235 3483 10238
rect 5993 10162 6059 10165
rect 17861 10162 17927 10165
rect 5993 10160 17927 10162
rect 5993 10104 5998 10160
rect 6054 10104 17866 10160
rect 17922 10104 17927 10160
rect 5993 10102 17927 10104
rect 5993 10099 6059 10102
rect 17861 10099 17927 10102
rect 5206 9964 5212 10028
rect 5276 10026 5282 10028
rect 21081 10026 21147 10029
rect 21357 10026 21423 10029
rect 5276 10024 21423 10026
rect 5276 9968 21086 10024
rect 21142 9968 21362 10024
rect 21418 9968 21423 10024
rect 5276 9966 21423 9968
rect 5276 9964 5282 9966
rect 21081 9963 21147 9966
rect 21357 9963 21423 9966
rect 0 9890 800 9920
rect 3325 9890 3391 9893
rect 0 9888 3391 9890
rect 0 9832 3330 9888
rect 3386 9832 3391 9888
rect 0 9830 3391 9832
rect 0 9800 800 9830
rect 3325 9827 3391 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 7833 9754 7899 9757
rect 7966 9754 7972 9756
rect 7833 9752 7972 9754
rect 7833 9696 7838 9752
rect 7894 9696 7972 9752
rect 7833 9694 7972 9696
rect 7833 9691 7899 9694
rect 7966 9692 7972 9694
rect 8036 9692 8042 9756
rect 9029 9618 9095 9621
rect 18137 9618 18203 9621
rect 9029 9616 18203 9618
rect 9029 9560 9034 9616
rect 9090 9560 18142 9616
rect 18198 9560 18203 9616
rect 9029 9558 18203 9560
rect 9029 9555 9095 9558
rect 18137 9555 18203 9558
rect 0 9482 800 9512
rect 3969 9482 4035 9485
rect 0 9480 4035 9482
rect 0 9424 3974 9480
rect 4030 9424 4035 9480
rect 0 9422 4035 9424
rect 0 9392 800 9422
rect 3969 9419 4035 9422
rect 7230 9420 7236 9484
rect 7300 9482 7306 9484
rect 15837 9482 15903 9485
rect 7300 9480 15903 9482
rect 7300 9424 15842 9480
rect 15898 9424 15903 9480
rect 7300 9422 15903 9424
rect 7300 9420 7306 9422
rect 15837 9419 15903 9422
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 0 9074 800 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 800 9014
rect 4061 9011 4127 9014
rect 5165 9074 5231 9077
rect 10317 9074 10383 9077
rect 5165 9072 10383 9074
rect 5165 9016 5170 9072
rect 5226 9016 10322 9072
rect 10378 9016 10383 9072
rect 5165 9014 10383 9016
rect 5165 9011 5231 9014
rect 10317 9011 10383 9014
rect 6144 8736 6460 8737
rect 0 8666 800 8696
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 3969 8666 4035 8669
rect 0 8664 4035 8666
rect 0 8608 3974 8664
rect 4030 8608 4035 8664
rect 0 8606 4035 8608
rect 0 8576 800 8606
rect 3969 8603 4035 8606
rect 0 8258 800 8288
rect 3049 8258 3115 8261
rect 0 8256 3115 8258
rect 0 8200 3054 8256
rect 3110 8200 3115 8256
rect 0 8198 3115 8200
rect 0 8168 800 8198
rect 3049 8195 3115 8198
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 13261 8124 13327 8125
rect 13261 8122 13308 8124
rect 13216 8120 13308 8122
rect 13216 8064 13266 8120
rect 13216 8062 13308 8064
rect 13261 8060 13308 8062
rect 13372 8060 13378 8124
rect 13261 8059 13327 8060
rect 0 7850 800 7880
rect 1485 7850 1551 7853
rect 0 7848 1551 7850
rect 0 7792 1490 7848
rect 1546 7792 1551 7848
rect 0 7790 1551 7792
rect 0 7760 800 7790
rect 1485 7787 1551 7790
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 0 7442 800 7472
rect 2773 7442 2839 7445
rect 0 7440 2839 7442
rect 0 7384 2778 7440
rect 2834 7384 2839 7440
rect 0 7382 2839 7384
rect 0 7352 800 7382
rect 2773 7379 2839 7382
rect 3545 7104 3861 7105
rect 0 7034 800 7064
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 3417 7034 3483 7037
rect 0 7032 3483 7034
rect 0 6976 3422 7032
rect 3478 6976 3483 7032
rect 0 6974 3483 6976
rect 0 6944 800 6974
rect 3417 6971 3483 6974
rect 0 6626 800 6656
rect 4061 6626 4127 6629
rect 0 6624 4127 6626
rect 0 6568 4066 6624
rect 4122 6568 4127 6624
rect 0 6566 4127 6568
rect 0 6536 800 6566
rect 4061 6563 4127 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 0 6218 800 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 800 6158
rect 4061 6155 4127 6158
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 0 5810 800 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 800 5750
rect 4061 5747 4127 5750
rect 6144 5472 6460 5473
rect 0 5402 800 5432
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 4061 5402 4127 5405
rect 0 5400 4127 5402
rect 0 5344 4066 5400
rect 4122 5344 4127 5400
rect 0 5342 4127 5344
rect 0 5312 800 5342
rect 4061 5339 4127 5342
rect 4153 5130 4219 5133
rect 2730 5128 4219 5130
rect 2730 5072 4158 5128
rect 4214 5072 4219 5128
rect 2730 5070 4219 5072
rect 0 4994 800 5024
rect 2730 4994 2790 5070
rect 4153 5067 4219 5070
rect 0 4934 2790 4994
rect 0 4904 800 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 0 4586 800 4616
rect 4429 4586 4495 4589
rect 0 4584 4495 4586
rect 0 4528 4434 4584
rect 4490 4528 4495 4584
rect 0 4526 4495 4528
rect 0 4496 800 4526
rect 4429 4523 4495 4526
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 0 4178 800 4208
rect 3969 4178 4035 4181
rect 0 4176 4035 4178
rect 0 4120 3974 4176
rect 4030 4120 4035 4176
rect 0 4118 4035 4120
rect 0 4088 800 4118
rect 3969 4115 4035 4118
rect 3545 3840 3861 3841
rect 0 3770 800 3800
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 3417 3770 3483 3773
rect 0 3768 3483 3770
rect 0 3712 3422 3768
rect 3478 3712 3483 3768
rect 0 3710 3483 3712
rect 0 3680 800 3710
rect 3417 3707 3483 3710
rect 0 3362 800 3392
rect 4061 3362 4127 3365
rect 0 3360 4127 3362
rect 0 3304 4066 3360
rect 4122 3304 4127 3360
rect 0 3302 4127 3304
rect 0 3272 800 3302
rect 4061 3299 4127 3302
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 0 2954 800 2984
rect 3969 2954 4035 2957
rect 0 2952 4035 2954
rect 0 2896 3974 2952
rect 4030 2896 4035 2952
rect 0 2894 4035 2896
rect 0 2864 800 2894
rect 3969 2891 4035 2894
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 0 2546 800 2576
rect 4061 2546 4127 2549
rect 0 2544 4127 2546
rect 0 2488 4066 2544
rect 4122 2488 4127 2544
rect 0 2486 4127 2488
rect 0 2456 800 2486
rect 4061 2483 4127 2486
rect 6144 2208 6460 2209
rect 0 2138 800 2168
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 3509 2138 3575 2141
rect 0 2136 3575 2138
rect 0 2080 3514 2136
rect 3570 2080 3575 2136
rect 0 2078 3575 2080
rect 0 2048 800 2078
rect 3509 2075 3575 2078
rect 0 1730 800 1760
rect 2865 1730 2931 1733
rect 0 1728 2931 1730
rect 0 1672 2870 1728
rect 2926 1672 2931 1728
rect 0 1670 2931 1672
rect 0 1640 800 1670
rect 2865 1667 2931 1670
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 6868 20224 6932 20228
rect 6868 20168 6882 20224
rect 6882 20168 6932 20224
rect 6868 20164 6932 20168
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 13308 17988 13372 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 7972 17912 8036 17916
rect 7972 17856 8022 17912
rect 8022 17856 8036 17912
rect 7972 17852 8036 17856
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 13124 17036 13188 17100
rect 5212 16960 5276 16964
rect 5212 16904 5226 16960
rect 5226 16904 5276 16960
rect 5212 16900 5276 16904
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 7236 16688 7300 16692
rect 7236 16632 7250 16688
rect 7250 16632 7300 16688
rect 7236 16628 7300 16632
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 6868 13772 6932 13836
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 13124 11188 13188 11252
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 5212 9964 5276 10028
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 7972 9692 8036 9756
rect 7236 9420 7300 9484
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 13308 8120 13372 8124
rect 13308 8064 13322 8120
rect 13322 8064 13372 8120
rect 13308 8060 13372 8064
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6867 20228 6933 20229
rect 6867 20164 6868 20228
rect 6932 20164 6933 20228
rect 6867 20163 6933 20164
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 5211 16964 5277 16965
rect 5211 16900 5212 16964
rect 5276 16900 5277 16964
rect 5211 16899 5277 16900
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 5214 10029 5274 16899
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6870 13837 6930 20163
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 7971 17916 8037 17917
rect 7971 17852 7972 17916
rect 8036 17852 8037 17916
rect 7971 17851 8037 17852
rect 7235 16692 7301 16693
rect 7235 16628 7236 16692
rect 7300 16628 7301 16692
rect 7235 16627 7301 16628
rect 6867 13836 6933 13837
rect 6867 13772 6868 13836
rect 6932 13772 6933 13836
rect 6867 13771 6933 13772
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 5211 10028 5277 10029
rect 5211 9964 5212 10028
rect 5276 9964 5277 10028
rect 5211 9963 5277 9964
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 7238 9485 7298 16627
rect 7974 9757 8034 17851
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 7971 9756 8037 9757
rect 7971 9692 7972 9756
rect 8036 9692 8037 9756
rect 7971 9691 8037 9692
rect 7235 9484 7301 9485
rect 7235 9420 7236 9484
rect 7300 9420 7301 9484
rect 7235 9419 7301 9420
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13307 18052 13373 18053
rect 13307 17988 13308 18052
rect 13372 17988 13373 18052
rect 13307 17987 13373 17988
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 13123 17100 13189 17101
rect 13123 17036 13124 17100
rect 13188 17036 13189 17100
rect 13123 17035 13189 17036
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 13126 11253 13186 17035
rect 13123 11252 13189 11253
rect 13123 11188 13124 11252
rect 13188 11188 13189 11252
rect 13123 11187 13189 11188
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 13310 8125 13370 17987
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13307 8124 13373 8125
rect 13307 8060 13308 8124
rect 13372 8060 13373 8124
rect 13307 8059 13373 8060
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1472 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform -1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1649977179
transform 1 0 4692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1649977179
transform -1 0 5612 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1649977179
transform -1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20884 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 19780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 19596 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 19596 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 19780 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 18676 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16652 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20884 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 20700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17204 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 19964 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 19964 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 21160 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 21344 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 19504 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20148 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 18676 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 19780 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16100 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20792 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 19504 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18216 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 19596 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 20700 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 19228 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 17020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17756 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18952 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18768 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 19504 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17756 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12328 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15548 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4784 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 5520 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6808 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 6624 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6440 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 7912 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1649977179
transform -1 0 4324 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 12788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 11316 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 10488 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 10120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1649977179
transform -1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10212 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 10580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 8004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 10764 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 11408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5152 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10028 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 11408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9844 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9384 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10120 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 7912 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 7544 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 7176 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6624 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 5152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 5244 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 7084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 5704 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 5060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 4048 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 4600 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 4968 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 5336 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 1656 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 1656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 1656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 3312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 4048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 5612 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 7544 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 2760 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7636 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 1564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 2668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 2668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 2944 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 1840 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 1564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5888 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 4508 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4232 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 5612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 8924 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 9752 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 9936 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 8096 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1649977179
transform -1 0 8280 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 2300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 4324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 1656 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 3312 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 4784 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 6992 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4048 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 5888 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 6440 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5888 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 3128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 5520 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6440 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6440 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3220 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 3036 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 7360 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 8188 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7728 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 9568 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_115
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_127
timestamp 1649977179
transform 1 0 12788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_139
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_151
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1649977179
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_87
timestamp 1649977179
transform 1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_91
timestamp 1649977179
transform 1 0 9476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_103
timestamp 1649977179
transform 1 0 10580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_115
timestamp 1649977179
transform 1 0 11684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_127
timestamp 1649977179
transform 1 0 12788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_49
timestamp 1649977179
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_60
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_64
timestamp 1649977179
transform 1 0 6992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_68
timestamp 1649977179
transform 1 0 7360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1649977179
transform 1 0 8280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_82
timestamp 1649977179
transform 1 0 8648 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_85
timestamp 1649977179
transform 1 0 8924 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_100
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_37
timestamp 1649977179
transform 1 0 4508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_47
timestamp 1649977179
transform 1 0 5428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_59
timestamp 1649977179
transform 1 0 6532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_63
timestamp 1649977179
transform 1 0 6900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_73
timestamp 1649977179
transform 1 0 7820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_95
timestamp 1649977179
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1649977179
transform 1 0 10212 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_113
timestamp 1649977179
transform 1 0 11500 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_117
timestamp 1649977179
transform 1 0 11868 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_129
timestamp 1649977179
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1649977179
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_47
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_50
timestamp 1649977179
transform 1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1649977179
transform 1 0 6808 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_73
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_77
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_88
timestamp 1649977179
transform 1 0 9200 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_92
timestamp 1649977179
transform 1 0 9568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_96
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_100
timestamp 1649977179
transform 1 0 10304 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_51
timestamp 1649977179
transform 1 0 5796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_62
timestamp 1649977179
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_66
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_76
timestamp 1649977179
transform 1 0 8096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_94
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_98
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_101
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_105
timestamp 1649977179
transform 1 0 10764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_112
timestamp 1649977179
transform 1 0 11408 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_116
timestamp 1649977179
transform 1 0 11776 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_130
timestamp 1649977179
transform 1 0 13064 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1649977179
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_42
timestamp 1649977179
transform 1 0 4968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_46
timestamp 1649977179
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_50
timestamp 1649977179
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1649977179
transform 1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_95
timestamp 1649977179
transform 1 0 9844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_99
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_117
timestamp 1649977179
transform 1 0 11868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_121
timestamp 1649977179
transform 1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_132
timestamp 1649977179
transform 1 0 13248 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_144
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_156
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_213
timestamp 1649977179
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1649977179
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_14
timestamp 1649977179
transform 1 0 2392 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1649977179
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_35
timestamp 1649977179
transform 1 0 4324 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 1649977179
transform 1 0 5336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_57
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_62
timestamp 1649977179
transform 1 0 6808 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_66
timestamp 1649977179
transform 1 0 7176 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_72
timestamp 1649977179
transform 1 0 7728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_112
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_123
timestamp 1649977179
transform 1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_127
timestamp 1649977179
transform 1 0 12788 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_135
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_163
timestamp 1649977179
transform 1 0 16100 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_175
timestamp 1649977179
transform 1 0 17204 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1649977179
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_199
timestamp 1649977179
transform 1 0 19412 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_205
timestamp 1649977179
transform 1 0 19964 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_211
timestamp 1649977179
transform 1 0 20516 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1649977179
transform 1 0 20884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1649977179
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_13
timestamp 1649977179
transform 1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_19
timestamp 1649977179
transform 1 0 2852 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_23
timestamp 1649977179
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp 1649977179
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_43
timestamp 1649977179
transform 1 0 5060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_47
timestamp 1649977179
transform 1 0 5428 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1649977179
transform 1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1649977179
transform 1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_74
timestamp 1649977179
transform 1 0 7912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_78
timestamp 1649977179
transform 1 0 8280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_88
timestamp 1649977179
transform 1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1649977179
transform 1 0 10212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1649977179
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1649977179
transform 1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_140
timestamp 1649977179
transform 1 0 13984 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_144
timestamp 1649977179
transform 1 0 14352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1649977179
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1649977179
transform 1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_179
timestamp 1649977179
transform 1 0 17572 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_187
timestamp 1649977179
transform 1 0 18308 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_191
timestamp 1649977179
transform 1 0 18676 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_195
timestamp 1649977179
transform 1 0 19044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_201
timestamp 1649977179
transform 1 0 19596 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_209
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_213
timestamp 1649977179
transform 1 0 20700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_13
timestamp 1649977179
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1649977179
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_31
timestamp 1649977179
transform 1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_42
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1649977179
transform 1 0 5336 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_49
timestamp 1649977179
transform 1 0 5612 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_60
timestamp 1649977179
transform 1 0 6624 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1649977179
transform 1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_94
timestamp 1649977179
transform 1 0 9752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_98
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_101
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_105
timestamp 1649977179
transform 1 0 10764 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_157
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_175
timestamp 1649977179
transform 1 0 17204 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1649977179
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_200
timestamp 1649977179
transform 1 0 19504 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_204
timestamp 1649977179
transform 1 0 19872 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_6
timestamp 1649977179
transform 1 0 1656 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_12
timestamp 1649977179
transform 1 0 2208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_20
timestamp 1649977179
transform 1 0 2944 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_28
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_32
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_40
timestamp 1649977179
transform 1 0 4784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_46
timestamp 1649977179
transform 1 0 5336 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_83
timestamp 1649977179
transform 1 0 8740 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_88
timestamp 1649977179
transform 1 0 9200 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_92
timestamp 1649977179
transform 1 0 9568 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_104
timestamp 1649977179
transform 1 0 10672 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_127
timestamp 1649977179
transform 1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1649977179
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_203
timestamp 1649977179
transform 1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_13
timestamp 1649977179
transform 1 0 2300 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_19
timestamp 1649977179
transform 1 0 2852 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_22
timestamp 1649977179
transform 1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_35
timestamp 1649977179
transform 1 0 4324 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_39
timestamp 1649977179
transform 1 0 4692 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_49
timestamp 1649977179
transform 1 0 5612 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_62
timestamp 1649977179
transform 1 0 6808 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_70
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_75
timestamp 1649977179
transform 1 0 8004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_94
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_98
timestamp 1649977179
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_108
timestamp 1649977179
transform 1 0 11040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_112
timestamp 1649977179
transform 1 0 11408 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1649977179
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_157
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_175
timestamp 1649977179
transform 1 0 17204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp 1649977179
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1649977179
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_217
timestamp 1649977179
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_13
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_17
timestamp 1649977179
transform 1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_21
timestamp 1649977179
transform 1 0 3036 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_24
timestamp 1649977179
transform 1 0 3312 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_28
timestamp 1649977179
transform 1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_32
timestamp 1649977179
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_60
timestamp 1649977179
transform 1 0 6624 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_64
timestamp 1649977179
transform 1 0 6992 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_68
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_72
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_89
timestamp 1649977179
transform 1 0 9292 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1649977179
transform 1 0 10212 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_116
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_135
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_143
timestamp 1649977179
transform 1 0 14260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1649977179
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_171
timestamp 1649977179
transform 1 0 16836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_177
timestamp 1649977179
transform 1 0 17388 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_196
timestamp 1649977179
transform 1 0 19136 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_200
timestamp 1649977179
transform 1 0 19504 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_7
timestamp 1649977179
transform 1 0 1748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_38
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_49
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_57
timestamp 1649977179
transform 1 0 6348 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_68
timestamp 1649977179
transform 1 0 7360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_73
timestamp 1649977179
transform 1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_94
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_102
timestamp 1649977179
transform 1 0 10488 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_105
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_120
timestamp 1649977179
transform 1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_147
timestamp 1649977179
transform 1 0 14628 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1649977179
transform 1 0 16468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_171
timestamp 1649977179
transform 1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1649977179
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_199
timestamp 1649977179
transform 1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_5
timestamp 1649977179
transform 1 0 1564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_13
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1649977179
transform 1 0 2668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_21
timestamp 1649977179
transform 1 0 3036 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_25
timestamp 1649977179
transform 1 0 3404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_30
timestamp 1649977179
transform 1 0 3864 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_34
timestamp 1649977179
transform 1 0 4232 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_66
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_70
timestamp 1649977179
transform 1 0 7544 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_80
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1649977179
transform 1 0 9476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_95
timestamp 1649977179
transform 1 0 9844 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_101
timestamp 1649977179
transform 1 0 10396 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_104
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1649977179
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_146
timestamp 1649977179
transform 1 0 14536 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_150
timestamp 1649977179
transform 1 0 14904 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_185
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_196
timestamp 1649977179
transform 1 0 19136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_200
timestamp 1649977179
transform 1 0 19504 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1649977179
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1649977179
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_40
timestamp 1649977179
transform 1 0 4784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_52
timestamp 1649977179
transform 1 0 5888 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_56
timestamp 1649977179
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1649977179
transform 1 0 7176 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp 1649977179
transform 1 0 7636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1649977179
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_87
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_91
timestamp 1649977179
transform 1 0 9476 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_100
timestamp 1649977179
transform 1 0 10304 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_104
timestamp 1649977179
transform 1 0 10672 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1649977179
transform 1 0 11684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_119
timestamp 1649977179
transform 1 0 12052 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_157
timestamp 1649977179
transform 1 0 15548 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_161
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_173
timestamp 1649977179
transform 1 0 17020 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_216
timestamp 1649977179
transform 1 0 20976 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_220
timestamp 1649977179
transform 1 0 21344 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_8
timestamp 1649977179
transform 1 0 1840 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_19
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_30
timestamp 1649977179
transform 1 0 3864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_35
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_50
timestamp 1649977179
transform 1 0 5704 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_67
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_72
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_84
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_88
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_92
timestamp 1649977179
transform 1 0 9568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 1649977179
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1649977179
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1649977179
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_154
timestamp 1649977179
transform 1 0 15272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1649977179
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_171
timestamp 1649977179
transform 1 0 16836 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1649977179
transform 1 0 20516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1649977179
transform 1 0 20884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1649977179
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_12
timestamp 1649977179
transform 1 0 2208 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_18
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_22
timestamp 1649977179
transform 1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_40
timestamp 1649977179
transform 1 0 4784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_44
timestamp 1649977179
transform 1 0 5152 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_48
timestamp 1649977179
transform 1 0 5520 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_52
timestamp 1649977179
transform 1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_58
timestamp 1649977179
transform 1 0 6440 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_62
timestamp 1649977179
transform 1 0 6808 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_70
timestamp 1649977179
transform 1 0 7544 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_74
timestamp 1649977179
transform 1 0 7912 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_94
timestamp 1649977179
transform 1 0 9752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_98
timestamp 1649977179
transform 1 0 10120 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_111
timestamp 1649977179
transform 1 0 11316 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_123
timestamp 1649977179
transform 1 0 12420 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_135
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1649977179
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_161
timestamp 1649977179
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_184
timestamp 1649977179
transform 1 0 18032 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_188
timestamp 1649977179
transform 1 0 18400 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1649977179
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_199
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_203
timestamp 1649977179
transform 1 0 19780 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_220
timestamp 1649977179
transform 1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_6
timestamp 1649977179
transform 1 0 1656 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_14
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_20
timestamp 1649977179
transform 1 0 2944 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1649977179
transform 1 0 4048 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_60
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1649977179
transform 1 0 7636 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_82
timestamp 1649977179
transform 1 0 8648 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_98
timestamp 1649977179
transform 1 0 10120 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_106
timestamp 1649977179
transform 1 0 10856 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_119
timestamp 1649977179
transform 1 0 12052 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_147
timestamp 1649977179
transform 1 0 14628 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1649977179
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_187
timestamp 1649977179
transform 1 0 18308 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_191
timestamp 1649977179
transform 1 0 18676 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_195
timestamp 1649977179
transform 1 0 19044 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_203
timestamp 1649977179
transform 1 0 19780 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1649977179
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_6
timestamp 1649977179
transform 1 0 1656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_12
timestamp 1649977179
transform 1 0 2208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_18
timestamp 1649977179
transform 1 0 2760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_22
timestamp 1649977179
transform 1 0 3128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1649977179
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1649977179
transform 1 0 4048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_36
timestamp 1649977179
transform 1 0 4416 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_47
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_58
timestamp 1649977179
transform 1 0 6440 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_69
timestamp 1649977179
transform 1 0 7452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_87
timestamp 1649977179
transform 1 0 9108 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_95
timestamp 1649977179
transform 1 0 9844 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_103
timestamp 1649977179
transform 1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_114
timestamp 1649977179
transform 1 0 11592 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_119
timestamp 1649977179
transform 1 0 12052 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_131
timestamp 1649977179
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_161
timestamp 1649977179
transform 1 0 15916 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_168
timestamp 1649977179
transform 1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1649977179
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_190
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_199
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_6
timestamp 1649977179
transform 1 0 1656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_12
timestamp 1649977179
transform 1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_22
timestamp 1649977179
transform 1 0 3128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_33
timestamp 1649977179
transform 1 0 4140 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_41
timestamp 1649977179
transform 1 0 4876 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1649977179
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_66
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_71
timestamp 1649977179
transform 1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_83
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_87
timestamp 1649977179
transform 1 0 9108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_91
timestamp 1649977179
transform 1 0 9476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1649977179
transform 1 0 10304 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_122
timestamp 1649977179
transform 1 0 12328 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_130
timestamp 1649977179
transform 1 0 13064 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_147
timestamp 1649977179
transform 1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_151
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1649977179
transform 1 0 15364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_159
timestamp 1649977179
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_185
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_189
timestamp 1649977179
transform 1 0 18492 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_211
timestamp 1649977179
transform 1 0 20516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_216
timestamp 1649977179
transform 1 0 20976 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_220
timestamp 1649977179
transform 1 0 21344 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_6
timestamp 1649977179
transform 1 0 1656 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_12
timestamp 1649977179
transform 1 0 2208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_18
timestamp 1649977179
transform 1 0 2760 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1649977179
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_31
timestamp 1649977179
transform 1 0 3956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_42
timestamp 1649977179
transform 1 0 4968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1649977179
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1649977179
transform 1 0 6348 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1649977179
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_72
timestamp 1649977179
transform 1 0 7728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1649977179
transform 1 0 9476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_98
timestamp 1649977179
transform 1 0 10120 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_111
timestamp 1649977179
transform 1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_116
timestamp 1649977179
transform 1 0 11776 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_175
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1649977179
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_12
timestamp 1649977179
transform 1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_21
timestamp 1649977179
transform 1 0 3036 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_32
timestamp 1649977179
transform 1 0 4048 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_36
timestamp 1649977179
transform 1 0 4416 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_46
timestamp 1649977179
transform 1 0 5336 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_66
timestamp 1649977179
transform 1 0 7176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_79
timestamp 1649977179
transform 1 0 8372 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_83
timestamp 1649977179
transform 1 0 8740 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_91
timestamp 1649977179
transform 1 0 9476 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_96
timestamp 1649977179
transform 1 0 9936 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_100
timestamp 1649977179
transform 1 0 10304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1649977179
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_145
timestamp 1649977179
transform 1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_159
timestamp 1649977179
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_173
timestamp 1649977179
transform 1 0 17020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1649977179
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_195
timestamp 1649977179
transform 1 0 19044 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_199
timestamp 1649977179
transform 1 0 19412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp 1649977179
transform 1 0 19780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_12
timestamp 1649977179
transform 1 0 2208 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_18
timestamp 1649977179
transform 1 0 2760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_22
timestamp 1649977179
transform 1 0 3128 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_45
timestamp 1649977179
transform 1 0 5244 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_56
timestamp 1649977179
transform 1 0 6256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_61
timestamp 1649977179
transform 1 0 6716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_66
timestamp 1649977179
transform 1 0 7176 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_71
timestamp 1649977179
transform 1 0 7636 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_94
timestamp 1649977179
transform 1 0 9752 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1649977179
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_102
timestamp 1649977179
transform 1 0 10488 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_114
timestamp 1649977179
transform 1 0 11592 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_157
timestamp 1649977179
transform 1 0 15548 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_161
timestamp 1649977179
transform 1 0 15916 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_179
timestamp 1649977179
transform 1 0 17572 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1649977179
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_187
timestamp 1649977179
transform 1 0 18308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_191
timestamp 1649977179
transform 1 0 18676 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_199
timestamp 1649977179
transform 1 0 19412 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_203
timestamp 1649977179
transform 1 0 19780 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_19
timestamp 1649977179
transform 1 0 2852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_24
timestamp 1649977179
transform 1 0 3312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_28
timestamp 1649977179
transform 1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1649977179
transform 1 0 4416 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_41
timestamp 1649977179
transform 1 0 4876 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_45
timestamp 1649977179
transform 1 0 5244 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_50
timestamp 1649977179
transform 1 0 5704 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_59
timestamp 1649977179
transform 1 0 6532 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_65
timestamp 1649977179
transform 1 0 7084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_76
timestamp 1649977179
transform 1 0 8096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_85
timestamp 1649977179
transform 1 0 8924 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_89
timestamp 1649977179
transform 1 0 9292 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1649977179
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_100
timestamp 1649977179
transform 1 0 10304 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1649977179
transform 1 0 12236 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_124
timestamp 1649977179
transform 1 0 12512 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_142
timestamp 1649977179
transform 1 0 14168 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_160
timestamp 1649977179
transform 1 0 15824 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_185
timestamp 1649977179
transform 1 0 18124 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1649977179
transform 1 0 19780 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_11
timestamp 1649977179
transform 1 0 2116 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_16
timestamp 1649977179
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_33
timestamp 1649977179
transform 1 0 4140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_40
timestamp 1649977179
transform 1 0 4784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_44
timestamp 1649977179
transform 1 0 5152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_48
timestamp 1649977179
transform 1 0 5520 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_54
timestamp 1649977179
transform 1 0 6072 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_58
timestamp 1649977179
transform 1 0 6440 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_69
timestamp 1649977179
transform 1 0 7452 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_90
timestamp 1649977179
transform 1 0 9384 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_100
timestamp 1649977179
transform 1 0 10304 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_112
timestamp 1649977179
transform 1 0 11408 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1649977179
transform 1 0 12144 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_157
timestamp 1649977179
transform 1 0 15548 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_161
timestamp 1649977179
transform 1 0 15916 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_179
timestamp 1649977179
transform 1 0 17572 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_183
timestamp 1649977179
transform 1 0 17940 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_187
timestamp 1649977179
transform 1 0 18308 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1649977179
transform 1 0 18584 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_213
timestamp 1649977179
transform 1 0 20700 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_217
timestamp 1649977179
transform 1 0 21068 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_12
timestamp 1649977179
transform 1 0 2208 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_24
timestamp 1649977179
transform 1 0 3312 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_31
timestamp 1649977179
transform 1 0 3956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_43
timestamp 1649977179
transform 1 0 5060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_49
timestamp 1649977179
transform 1 0 5612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1649977179
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_63
timestamp 1649977179
transform 1 0 6900 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_74
timestamp 1649977179
transform 1 0 7912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_78
timestamp 1649977179
transform 1 0 8280 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_87
timestamp 1649977179
transform 1 0 9108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_99
timestamp 1649977179
transform 1 0 10212 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_121
timestamp 1649977179
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_157
timestamp 1649977179
transform 1 0 15548 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_185
timestamp 1649977179
transform 1 0 18124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_189
timestamp 1649977179
transform 1 0 18492 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_196
timestamp 1649977179
transform 1 0 19136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_200
timestamp 1649977179
transform 1 0 19504 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_218
timestamp 1649977179
transform 1 0 21160 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1649977179
transform 1 0 21528 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_13
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1649977179
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1649977179
transform 1 0 4048 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_36
timestamp 1649977179
transform 1 0 4416 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_44
timestamp 1649977179
transform 1 0 5152 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_55
timestamp 1649977179
transform 1 0 6164 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_66
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1649977179
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_87
timestamp 1649977179
transform 1 0 9108 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1649977179
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_99
timestamp 1649977179
transform 1 0 10212 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_105
timestamp 1649977179
transform 1 0 10764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_114
timestamp 1649977179
transform 1 0 11592 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_126
timestamp 1649977179
transform 1 0 12696 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1649977179
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_143
timestamp 1649977179
transform 1 0 14260 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_147
timestamp 1649977179
transform 1 0 14628 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_159
timestamp 1649977179
transform 1 0 15732 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_171
timestamp 1649977179
transform 1 0 16836 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1649977179
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_199
timestamp 1649977179
transform 1 0 19412 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1649977179
transform 1 0 19780 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_35
timestamp 1649977179
transform 1 0 4324 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_38
timestamp 1649977179
transform 1 0 4600 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_42
timestamp 1649977179
transform 1 0 4968 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_46
timestamp 1649977179
transform 1 0 5336 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_50
timestamp 1649977179
transform 1 0 5704 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_66
timestamp 1649977179
transform 1 0 7176 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_72
timestamp 1649977179
transform 1 0 7728 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_76
timestamp 1649977179
transform 1 0 8096 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_82
timestamp 1649977179
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_89
timestamp 1649977179
transform 1 0 9292 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_95
timestamp 1649977179
transform 1 0 9844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1649977179
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1649977179
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1649977179
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_189
timestamp 1649977179
transform 1 0 18492 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_194
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_199
timestamp 1649977179
transform 1 0 19412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_203
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_207
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1649977179
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1649977179
transform 1 0 4600 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1649977179
transform -1 0 6072 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1649977179
transform -1 0 3496 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1649977179
transform -1 0 8648 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1649977179
transform -1 0 8648 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1649977179
transform 1 0 7728 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1649977179
transform -1 0 10948 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1649977179
transform 1 0 11316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1649977179
transform 1 0 11776 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1649977179
transform -1 0 11776 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1649977179
transform -1 0 10304 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1649977179
transform -1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1649977179
transform -1 0 8648 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1649977179
transform -1 0 9200 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1649977179
transform -1 0 7636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1649977179
transform 1 0 4416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1649977179
transform -1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1649977179
transform 1 0 6532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1649977179
transform -1 0 11224 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1649977179
transform 1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1649977179
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1649977179
transform 1 0 9844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1649977179
transform 1 0 7360 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1649977179
transform 1 0 7360 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1649977179
transform -1 0 6624 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1649977179
transform 1 0 8280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1649977179
transform 1 0 5152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _068_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2392 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1649977179
transform -1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1649977179
transform -1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1649977179
transform -1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1649977179
transform 1 0 2392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1649977179
transform -1 0 2208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1649977179
transform 1 0 2576 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1649977179
transform -1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1649977179
transform -1 0 2208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1649977179
transform -1 0 2208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1649977179
transform -1 0 2760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1649977179
transform -1 0 2576 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1649977179
transform -1 0 2760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1649977179
transform -1 0 2208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1649977179
transform -1 0 2300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1649977179
transform -1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1649977179
transform 1 0 8280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1649977179
transform 1 0 7360 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1649977179
transform 1 0 10396 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1649977179
transform 1 0 6532 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1649977179
transform 1 0 9476 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1649977179
transform 1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1649977179
transform -1 0 10764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1649977179
transform -1 0 10212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1649977179
transform -1 0 9660 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1649977179
transform -1 0 9660 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1649977179
transform -1 0 9384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1649977179
transform -1 0 9292 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1649977179
transform 1 0 10120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1649977179
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1649977179
transform 1 0 1840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1649977179
transform 1 0 5060 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1649977179
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1649977179
transform 1 0 6164 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1649977179
transform 1 0 10856 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19412 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21436 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18308 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13800 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16744 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17572 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19044 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21344 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14628 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21436 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14536 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13616 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12144 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13524 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16100 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13800 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14444 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13616 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17204 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14996 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21068 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17204 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14536 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19964 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20976 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20516 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19136 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18308 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18676 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16376 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14444 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21252 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18032 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13156 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19596 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18952 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16100 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21160 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19780 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17572 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13892 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12696 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13708 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15824 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13800 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6992 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5520 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4508 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4508 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8372 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6072 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9108 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9016 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8372 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6072 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12420 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7544 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4784 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12144 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10212 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3680 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10856 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7636 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2392 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8832 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3128 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3496 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6808 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4876 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7268 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6716 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2944 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4784 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3036 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5428 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4416 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4048 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6164 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5152 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3220 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2852 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5612 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5060 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5428 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7268 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7636 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8096 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2668 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3036 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2852 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3496 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5704 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5520 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7544 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7176 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7912 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8096 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3956 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3956 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4048 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4600 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6072 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7912 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8924 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5888 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10488 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10304 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7452 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10488 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5060 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10764 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10856 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7452 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10580 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5796 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11316 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7360 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10120 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6808 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9752 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8004 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9384 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5612 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10580 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
<< labels >>
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 22200 11432 23000 11552 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 4 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 5 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 6 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 7 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 8 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 9 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 10 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 11 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 12 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 13 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 14 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 15 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 16 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 17 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 18 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 19 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 20 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 21 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 22 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 23 nsew signal input
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 24 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 25 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 26 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 27 nsew signal tristate
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 28 nsew signal tristate
flabel metal3 s 0 19184 800 19304 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 29 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 30 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 31 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 32 nsew signal tristate
flabel metal3 s 0 20816 800 20936 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 33 nsew signal tristate
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 34 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 35 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 36 nsew signal tristate
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 37 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 38 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 39 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 40 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 41 nsew signal tristate
flabel metal3 s 0 16736 800 16856 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 42 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 43 nsew signal tristate
flabel metal2 s 3882 22200 3938 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 44 nsew signal input
flabel metal2 s 8482 22200 8538 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 45 nsew signal input
flabel metal2 s 8942 22200 8998 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 46 nsew signal input
flabel metal2 s 9402 22200 9458 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 47 nsew signal input
flabel metal2 s 9862 22200 9918 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 48 nsew signal input
flabel metal2 s 10322 22200 10378 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 49 nsew signal input
flabel metal2 s 10782 22200 10838 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 50 nsew signal input
flabel metal2 s 11242 22200 11298 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 51 nsew signal input
flabel metal2 s 11702 22200 11758 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 52 nsew signal input
flabel metal2 s 12162 22200 12218 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 53 nsew signal input
flabel metal2 s 12622 22200 12678 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 54 nsew signal input
flabel metal2 s 4342 22200 4398 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 55 nsew signal input
flabel metal2 s 4802 22200 4858 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 56 nsew signal input
flabel metal2 s 5262 22200 5318 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 57 nsew signal input
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 58 nsew signal input
flabel metal2 s 6182 22200 6238 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 59 nsew signal input
flabel metal2 s 6642 22200 6698 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 60 nsew signal input
flabel metal2 s 7102 22200 7158 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 61 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 62 nsew signal input
flabel metal2 s 8022 22200 8078 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 63 nsew signal input
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 64 nsew signal tristate
flabel metal2 s 17682 22200 17738 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 65 nsew signal tristate
flabel metal2 s 18142 22200 18198 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 66 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 67 nsew signal tristate
flabel metal2 s 19062 22200 19118 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 68 nsew signal tristate
flabel metal2 s 19522 22200 19578 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 69 nsew signal tristate
flabel metal2 s 19982 22200 20038 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 70 nsew signal tristate
flabel metal2 s 20442 22200 20498 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 71 nsew signal tristate
flabel metal2 s 20902 22200 20958 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 72 nsew signal tristate
flabel metal2 s 21362 22200 21418 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 73 nsew signal tristate
flabel metal2 s 21822 22200 21878 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 74 nsew signal tristate
flabel metal2 s 13542 22200 13598 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 75 nsew signal tristate
flabel metal2 s 14002 22200 14058 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 76 nsew signal tristate
flabel metal2 s 14462 22200 14518 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 77 nsew signal tristate
flabel metal2 s 14922 22200 14978 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 78 nsew signal tristate
flabel metal2 s 15382 22200 15438 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 79 nsew signal tristate
flabel metal2 s 15842 22200 15898 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 80 nsew signal tristate
flabel metal2 s 16302 22200 16358 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 81 nsew signal tristate
flabel metal2 s 16762 22200 16818 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 82 nsew signal tristate
flabel metal2 s 17222 22200 17278 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 83 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 left_bottom_grid_pin_11_
port 84 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 left_bottom_grid_pin_13_
port 85 nsew signal input
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 left_bottom_grid_pin_15_
port 86 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 left_bottom_grid_pin_17_
port 87 nsew signal input
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 left_bottom_grid_pin_1_
port 88 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 left_bottom_grid_pin_3_
port 89 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 left_bottom_grid_pin_5_
port 90 nsew signal input
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 left_bottom_grid_pin_7_
port 91 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 left_bottom_grid_pin_9_
port 92 nsew signal input
flabel metal2 s 22282 22200 22338 23000 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 93 nsew signal input
flabel metal2 s 202 22200 258 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_42_
port 94 nsew signal input
flabel metal2 s 662 22200 718 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_43_
port 95 nsew signal input
flabel metal2 s 1122 22200 1178 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_44_
port 96 nsew signal input
flabel metal2 s 1582 22200 1638 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_45_
port 97 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_46_
port 98 nsew signal input
flabel metal2 s 2502 22200 2558 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_47_
port 99 nsew signal input
flabel metal2 s 2962 22200 3018 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_48_
port 100 nsew signal input
flabel metal2 s 3422 22200 3478 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_49_
port 101 nsew signal input
flabel metal2 s 22742 22200 22798 23000 0 FreeSans 224 90 0 0 top_right_grid_pin_1_
port 102 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
